magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect 1158 -1981 1192 -1905
rect 1158 -2071 1192 -2065
rect 1544 -1981 1578 -1905
rect 1544 -2071 1578 -2065
rect 1650 -2105 1684 -1905
rect 1650 -2195 1684 -2189
rect 2036 -2105 2070 -1905
rect 2036 -2195 2070 -2189
<< viali >>
rect 1158 -2065 1192 -1981
rect 1544 -2065 1578 -1981
rect 1650 -2189 1684 -2105
rect 2036 -2189 2070 -2105
<< metal1 >>
rect 1322 -882 1342 -830
rect 1394 -882 1414 -830
rect 1252 -972 1258 -920
rect 1310 -972 1316 -920
rect 1252 -1044 1316 -972
rect 1252 -1096 1258 -1044
rect 1310 -1096 1316 -1044
rect 1252 -1168 1316 -1096
rect 1252 -1220 1258 -1168
rect 1310 -1220 1316 -1168
rect 1420 -972 1426 -920
rect 1478 -972 1484 -920
rect 1420 -1044 1484 -972
rect 1420 -1096 1426 -1044
rect 1478 -1096 1484 -1044
rect 1420 -1168 1484 -1096
rect 1420 -1220 1426 -1168
rect 1478 -1220 1484 -1168
rect 1322 -1310 1342 -1258
rect 1394 -1310 1414 -1258
rect 1814 -1318 1834 -1266
rect 1886 -1318 1906 -1266
rect 1322 -1418 1342 -1366
rect 1394 -1418 1414 -1366
rect 1744 -1395 1808 -1347
rect 1744 -1447 1750 -1395
rect 1802 -1447 1808 -1395
rect 1912 -1395 1976 -1347
rect 1912 -1447 1918 -1395
rect 1970 -1447 1976 -1395
rect 1252 -1508 1258 -1456
rect 1310 -1508 1316 -1456
rect 1252 -1580 1316 -1508
rect 1252 -1632 1258 -1580
rect 1310 -1632 1316 -1580
rect 1252 -1704 1316 -1632
rect 1252 -1756 1258 -1704
rect 1310 -1756 1316 -1704
rect 1420 -1508 1426 -1456
rect 1478 -1508 1484 -1456
rect 1420 -1580 1484 -1508
rect 1814 -1528 1834 -1476
rect 1886 -1528 1906 -1476
rect 1420 -1632 1426 -1580
rect 1478 -1632 1484 -1580
rect 1420 -1665 1484 -1632
rect 1814 -1636 1834 -1584
rect 1886 -1636 1906 -1584
rect 1420 -1704 1808 -1665
rect 1420 -1756 1426 -1704
rect 1478 -1713 1808 -1704
rect 1478 -1756 1750 -1713
rect 1420 -1765 1750 -1756
rect 1802 -1765 1808 -1713
rect 1912 -1713 1976 -1665
rect 1912 -1765 1918 -1713
rect 1970 -1765 1976 -1713
rect 1322 -1846 1342 -1794
rect 1394 -1846 1414 -1794
rect 1814 -1846 1834 -1794
rect 1886 -1846 1906 -1794
rect 1252 -1932 1258 -1880
rect 1310 -1932 1918 -1880
rect 1970 -1932 1976 -1880
rect 1122 -1981 2106 -1975
rect 1122 -2065 1158 -1981
rect 1192 -2065 1544 -1981
rect 1578 -2065 2106 -1981
rect 1122 -2071 2106 -2065
rect 1122 -2105 2106 -2099
rect 1122 -2189 1650 -2105
rect 1684 -2189 2036 -2105
rect 2070 -2189 2106 -2105
rect 1122 -2195 2106 -2189
rect 1122 -2275 1258 -2223
rect 1310 -2275 2106 -2223
rect 1122 -2281 2106 -2275
<< via1 >>
rect 1342 -882 1394 -830
rect 1258 -972 1310 -920
rect 1258 -1096 1310 -1044
rect 1258 -1220 1310 -1168
rect 1426 -972 1478 -920
rect 1426 -1096 1478 -1044
rect 1426 -1220 1478 -1168
rect 1342 -1310 1394 -1258
rect 1834 -1318 1886 -1266
rect 1342 -1418 1394 -1366
rect 1750 -1447 1802 -1395
rect 1918 -1447 1970 -1395
rect 1258 -1508 1310 -1456
rect 1258 -1632 1310 -1580
rect 1258 -1756 1310 -1704
rect 1426 -1508 1478 -1456
rect 1834 -1528 1886 -1476
rect 1426 -1632 1478 -1580
rect 1834 -1636 1886 -1584
rect 1426 -1756 1478 -1704
rect 1750 -1765 1802 -1713
rect 1918 -1765 1970 -1713
rect 1342 -1846 1394 -1794
rect 1834 -1846 1886 -1794
rect 1258 -1932 1310 -1880
rect 1918 -1932 1970 -1880
rect 1258 -2275 1310 -2223
<< metal2 >>
rect 1340 -830 1396 -824
rect 1340 -882 1342 -830
rect 1394 -882 1396 -830
rect 1256 -920 1312 -914
rect 1256 -972 1258 -920
rect 1310 -972 1312 -920
rect 1256 -1044 1312 -972
rect 1256 -1096 1258 -1044
rect 1310 -1096 1312 -1044
rect 1256 -1168 1312 -1096
rect 1256 -1220 1258 -1168
rect 1310 -1220 1312 -1168
rect 1256 -1456 1312 -1220
rect 1256 -1508 1258 -1456
rect 1310 -1508 1312 -1456
rect 1256 -1580 1312 -1508
rect 1256 -1632 1258 -1580
rect 1310 -1632 1312 -1580
rect 1256 -1704 1312 -1632
rect 1256 -1756 1258 -1704
rect 1310 -1756 1312 -1704
rect 1256 -1880 1312 -1756
rect 1340 -1258 1396 -882
rect 1340 -1310 1342 -1258
rect 1394 -1310 1396 -1258
rect 1340 -1366 1396 -1310
rect 1340 -1418 1342 -1366
rect 1394 -1418 1396 -1366
rect 1340 -1794 1396 -1418
rect 1424 -920 1480 -914
rect 1424 -972 1426 -920
rect 1478 -972 1480 -920
rect 1424 -1044 1480 -972
rect 1424 -1096 1426 -1044
rect 1478 -1096 1480 -1044
rect 1424 -1168 1480 -1096
rect 1424 -1220 1426 -1168
rect 1478 -1220 1480 -1168
rect 1424 -1456 1480 -1220
rect 1832 -1266 1888 -1260
rect 1832 -1318 1834 -1266
rect 1886 -1318 1888 -1266
rect 1424 -1508 1426 -1456
rect 1478 -1508 1480 -1456
rect 1424 -1580 1480 -1508
rect 1424 -1632 1426 -1580
rect 1478 -1632 1480 -1580
rect 1424 -1704 1480 -1632
rect 1424 -1756 1426 -1704
rect 1478 -1756 1480 -1704
rect 1424 -1762 1480 -1756
rect 1748 -1395 1804 -1389
rect 1748 -1447 1750 -1395
rect 1802 -1447 1804 -1395
rect 1748 -1713 1804 -1447
rect 1748 -1765 1750 -1713
rect 1802 -1765 1804 -1713
rect 1748 -1771 1804 -1765
rect 1832 -1476 1888 -1318
rect 1832 -1528 1834 -1476
rect 1886 -1528 1888 -1476
rect 1832 -1584 1888 -1528
rect 1832 -1636 1834 -1584
rect 1886 -1636 1888 -1584
rect 1340 -1846 1342 -1794
rect 1394 -1846 1396 -1794
rect 1340 -1852 1396 -1846
rect 1832 -1794 1888 -1636
rect 1832 -1846 1834 -1794
rect 1886 -1846 1888 -1794
rect 1832 -1852 1888 -1846
rect 1916 -1395 1972 -1389
rect 1916 -1447 1918 -1395
rect 1970 -1447 1972 -1395
rect 1916 -1713 1972 -1447
rect 1916 -1765 1918 -1713
rect 1970 -1765 1972 -1713
rect 1256 -1932 1258 -1880
rect 1310 -1932 1312 -1880
rect 1256 -2223 1312 -1932
rect 1916 -1880 1972 -1765
rect 1916 -1932 1918 -1880
rect 1970 -1932 1972 -1880
rect 1916 -1938 1972 -1932
rect 1256 -2275 1258 -2223
rect 1310 -2275 1312 -2223
rect 1256 -2281 1312 -2275
use sky130_fd_pr__nfet_01v8_DJGLWN  sky130_fd_pr__nfet_01v8_DJGLWN_0
timestamp 1730624594
transform 1 0 1860 0 1 -1556
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_TMYQY6  sky130_fd_pr__pfet_01v8_TMYQY6_0
timestamp 1730624594
transform 1 0 1368 0 1 -1338
box -246 -637 246 637
<< labels >>
flabel metal1 1122 -2071 1218 -1975 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel metal1 1122 -2195 1218 -2099 0 FreeSans 320 0 0 0 vssa
port 4 nsew
flabel metal1 1122 -2281 1180 -2223 0 FreeSans 320 0 0 0 in
port 5 nsew
flabel via1 1342 -1846 1394 -1794 0 FreeSans 320 0 0 0 swp
port 2 nsew
flabel via1 1834 -1846 1886 -1794 0 FreeSans 320 0 0 0 swn
port 3 nsew
flabel via1 1426 -972 1478 -920 0 FreeSans 320 0 0 0 out
port 6 nsew
<< end >>
