magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect 360 -2065 394 -1989
rect 360 -2155 394 -2149
rect 746 -2065 780 -1989
rect 746 -2155 780 -2149
rect 852 -2189 886 -1989
rect 852 -2279 886 -2273
rect 1238 -2189 1272 -1989
rect 1238 -2279 1272 -2273
<< viali >>
rect 360 -2149 394 -2065
rect 746 -2149 780 -2065
rect 852 -2273 886 -2189
rect 1238 -2273 1272 -2189
<< metal1 >>
rect 524 106 544 158
rect 596 106 616 158
rect 454 16 460 68
rect 512 16 518 68
rect 454 -56 518 16
rect 454 -108 460 -56
rect 512 -108 518 -56
rect 454 -180 518 -108
rect 454 -232 460 -180
rect 512 -232 518 -180
rect 622 16 628 68
rect 680 16 686 68
rect 622 -56 686 16
rect 622 -108 628 -56
rect 680 -108 686 -56
rect 622 -180 686 -108
rect 622 -232 628 -180
rect 680 -232 686 -180
rect 524 -322 544 -270
rect 596 -322 616 -270
rect 524 -430 544 -378
rect 596 -430 616 -378
rect 454 -520 460 -468
rect 512 -520 518 -468
rect 454 -592 518 -520
rect 454 -644 460 -592
rect 512 -644 518 -592
rect 454 -716 518 -644
rect 454 -768 460 -716
rect 512 -768 518 -716
rect 622 -520 628 -468
rect 680 -520 686 -468
rect 622 -592 686 -520
rect 622 -644 628 -592
rect 680 -644 686 -592
rect 622 -716 686 -644
rect 622 -768 628 -716
rect 680 -768 686 -716
rect 1016 -766 1036 -714
rect 1088 -766 1108 -714
rect 524 -858 544 -806
rect 596 -858 616 -806
rect 946 -843 1010 -795
rect 946 -895 952 -843
rect 1004 -895 1010 -843
rect 1114 -843 1178 -795
rect 1114 -895 1120 -843
rect 1172 -895 1178 -843
rect 524 -966 544 -914
rect 596 -966 616 -914
rect 1016 -976 1036 -924
rect 1088 -976 1108 -924
rect 454 -1056 460 -1004
rect 512 -1056 518 -1004
rect 454 -1128 518 -1056
rect 454 -1180 460 -1128
rect 512 -1180 518 -1128
rect 454 -1252 518 -1180
rect 454 -1304 460 -1252
rect 512 -1304 518 -1252
rect 622 -1056 628 -1004
rect 680 -1056 686 -1004
rect 622 -1113 686 -1056
rect 1016 -1084 1036 -1032
rect 1088 -1084 1108 -1032
rect 622 -1128 1010 -1113
rect 622 -1180 628 -1128
rect 680 -1161 1010 -1128
rect 680 -1180 952 -1161
rect 622 -1213 952 -1180
rect 1004 -1213 1010 -1161
rect 1114 -1161 1178 -1113
rect 1114 -1213 1120 -1161
rect 1172 -1213 1178 -1161
rect 622 -1252 686 -1213
rect 622 -1304 628 -1252
rect 680 -1304 686 -1252
rect 1016 -1294 1036 -1242
rect 1088 -1294 1108 -1242
rect 524 -1394 544 -1342
rect 596 -1394 616 -1342
rect 1016 -1402 1036 -1350
rect 1088 -1402 1108 -1350
rect 524 -1502 544 -1450
rect 596 -1502 616 -1450
rect 946 -1479 1010 -1431
rect 946 -1531 952 -1479
rect 1004 -1531 1010 -1479
rect 1114 -1479 1178 -1431
rect 1114 -1531 1120 -1479
rect 1172 -1531 1178 -1479
rect 454 -1592 460 -1540
rect 512 -1592 518 -1540
rect 454 -1664 518 -1592
rect 454 -1716 460 -1664
rect 512 -1716 518 -1664
rect 454 -1788 518 -1716
rect 454 -1840 460 -1788
rect 512 -1840 518 -1788
rect 622 -1592 628 -1540
rect 680 -1592 686 -1540
rect 622 -1664 686 -1592
rect 1016 -1612 1036 -1560
rect 1088 -1612 1108 -1560
rect 622 -1716 628 -1664
rect 680 -1716 686 -1664
rect 622 -1749 686 -1716
rect 1016 -1720 1036 -1668
rect 1088 -1720 1108 -1668
rect 622 -1788 1010 -1749
rect 622 -1840 628 -1788
rect 680 -1797 1010 -1788
rect 680 -1840 952 -1797
rect 622 -1849 952 -1840
rect 1004 -1849 1010 -1797
rect 1114 -1797 1178 -1749
rect 1114 -1849 1120 -1797
rect 1172 -1849 1178 -1797
rect 524 -1930 544 -1878
rect 596 -1930 616 -1878
rect 1016 -1930 1036 -1878
rect 1088 -1930 1108 -1878
rect 454 -2016 460 -1964
rect 512 -2016 1120 -1964
rect 1172 -2016 1178 -1964
rect 324 -2065 1308 -2059
rect 324 -2149 360 -2065
rect 394 -2149 746 -2065
rect 780 -2149 1308 -2065
rect 324 -2155 1308 -2149
rect 324 -2189 1308 -2183
rect 324 -2273 852 -2189
rect 886 -2273 1238 -2189
rect 1272 -2273 1308 -2189
rect 324 -2279 1308 -2273
rect 324 -2359 460 -2307
rect 512 -2359 1308 -2307
rect 324 -2365 1308 -2359
<< via1 >>
rect 544 106 596 158
rect 460 16 512 68
rect 460 -108 512 -56
rect 460 -232 512 -180
rect 628 16 680 68
rect 628 -108 680 -56
rect 628 -232 680 -180
rect 544 -322 596 -270
rect 544 -430 596 -378
rect 460 -520 512 -468
rect 460 -644 512 -592
rect 460 -768 512 -716
rect 628 -520 680 -468
rect 628 -644 680 -592
rect 628 -768 680 -716
rect 1036 -766 1088 -714
rect 544 -858 596 -806
rect 952 -895 1004 -843
rect 1120 -895 1172 -843
rect 544 -966 596 -914
rect 1036 -976 1088 -924
rect 460 -1056 512 -1004
rect 460 -1180 512 -1128
rect 460 -1304 512 -1252
rect 628 -1056 680 -1004
rect 1036 -1084 1088 -1032
rect 628 -1180 680 -1128
rect 952 -1213 1004 -1161
rect 1120 -1213 1172 -1161
rect 628 -1304 680 -1252
rect 1036 -1294 1088 -1242
rect 544 -1394 596 -1342
rect 1036 -1402 1088 -1350
rect 544 -1502 596 -1450
rect 952 -1531 1004 -1479
rect 1120 -1531 1172 -1479
rect 460 -1592 512 -1540
rect 460 -1716 512 -1664
rect 460 -1840 512 -1788
rect 628 -1592 680 -1540
rect 1036 -1612 1088 -1560
rect 628 -1716 680 -1664
rect 1036 -1720 1088 -1668
rect 628 -1840 680 -1788
rect 952 -1849 1004 -1797
rect 1120 -1849 1172 -1797
rect 544 -1930 596 -1878
rect 1036 -1930 1088 -1878
rect 460 -2016 512 -1964
rect 1120 -2016 1172 -1964
rect 460 -2359 512 -2307
<< metal2 >>
rect 542 158 598 164
rect 542 106 544 158
rect 596 106 598 158
rect 458 68 514 74
rect 458 16 460 68
rect 512 16 514 68
rect 458 -56 514 16
rect 458 -108 460 -56
rect 512 -108 514 -56
rect 458 -180 514 -108
rect 458 -232 460 -180
rect 512 -232 514 -180
rect 458 -468 514 -232
rect 458 -520 460 -468
rect 512 -520 514 -468
rect 458 -592 514 -520
rect 458 -644 460 -592
rect 512 -644 514 -592
rect 458 -716 514 -644
rect 458 -768 460 -716
rect 512 -768 514 -716
rect 458 -1004 514 -768
rect 458 -1056 460 -1004
rect 512 -1056 514 -1004
rect 458 -1128 514 -1056
rect 458 -1180 460 -1128
rect 512 -1180 514 -1128
rect 458 -1252 514 -1180
rect 458 -1304 460 -1252
rect 512 -1304 514 -1252
rect 458 -1540 514 -1304
rect 458 -1592 460 -1540
rect 512 -1592 514 -1540
rect 458 -1664 514 -1592
rect 458 -1716 460 -1664
rect 512 -1716 514 -1664
rect 458 -1788 514 -1716
rect 458 -1840 460 -1788
rect 512 -1840 514 -1788
rect 458 -1964 514 -1840
rect 542 -270 598 106
rect 542 -322 544 -270
rect 596 -322 598 -270
rect 542 -378 598 -322
rect 542 -430 544 -378
rect 596 -430 598 -378
rect 542 -806 598 -430
rect 542 -858 544 -806
rect 596 -858 598 -806
rect 542 -914 598 -858
rect 542 -966 544 -914
rect 596 -966 598 -914
rect 542 -1342 598 -966
rect 542 -1394 544 -1342
rect 596 -1394 598 -1342
rect 542 -1450 598 -1394
rect 542 -1502 544 -1450
rect 596 -1502 598 -1450
rect 542 -1878 598 -1502
rect 626 68 682 74
rect 626 16 628 68
rect 680 16 682 68
rect 626 -56 682 16
rect 626 -108 628 -56
rect 680 -108 682 -56
rect 626 -180 682 -108
rect 626 -232 628 -180
rect 680 -232 682 -180
rect 626 -468 682 -232
rect 626 -520 628 -468
rect 680 -520 682 -468
rect 626 -592 682 -520
rect 626 -644 628 -592
rect 680 -644 682 -592
rect 626 -716 682 -644
rect 626 -768 628 -716
rect 680 -768 682 -716
rect 626 -1004 682 -768
rect 1034 -714 1090 -708
rect 1034 -766 1036 -714
rect 1088 -766 1090 -714
rect 626 -1056 628 -1004
rect 680 -1056 682 -1004
rect 626 -1128 682 -1056
rect 626 -1180 628 -1128
rect 680 -1180 682 -1128
rect 626 -1252 682 -1180
rect 626 -1304 628 -1252
rect 680 -1304 682 -1252
rect 626 -1540 682 -1304
rect 626 -1592 628 -1540
rect 680 -1592 682 -1540
rect 626 -1664 682 -1592
rect 626 -1716 628 -1664
rect 680 -1716 682 -1664
rect 626 -1788 682 -1716
rect 626 -1840 628 -1788
rect 680 -1840 682 -1788
rect 626 -1846 682 -1840
rect 950 -843 1006 -789
rect 950 -895 952 -843
rect 1004 -895 1006 -843
rect 950 -1161 1006 -895
rect 950 -1213 952 -1161
rect 1004 -1213 1006 -1161
rect 950 -1479 1006 -1213
rect 950 -1531 952 -1479
rect 1004 -1531 1006 -1479
rect 950 -1797 1006 -1531
rect 950 -1849 952 -1797
rect 1004 -1849 1006 -1797
rect 950 -1855 1006 -1849
rect 1034 -924 1090 -766
rect 1034 -976 1036 -924
rect 1088 -976 1090 -924
rect 1034 -1032 1090 -976
rect 1034 -1084 1036 -1032
rect 1088 -1084 1090 -1032
rect 1034 -1242 1090 -1084
rect 1034 -1294 1036 -1242
rect 1088 -1294 1090 -1242
rect 1034 -1350 1090 -1294
rect 1034 -1402 1036 -1350
rect 1088 -1402 1090 -1350
rect 1034 -1560 1090 -1402
rect 1034 -1612 1036 -1560
rect 1088 -1612 1090 -1560
rect 1034 -1668 1090 -1612
rect 1034 -1720 1036 -1668
rect 1088 -1720 1090 -1668
rect 542 -1930 544 -1878
rect 596 -1930 598 -1878
rect 542 -1936 598 -1930
rect 1034 -1878 1090 -1720
rect 1034 -1930 1036 -1878
rect 1088 -1930 1090 -1878
rect 1034 -1936 1090 -1930
rect 1118 -843 1174 -789
rect 1118 -895 1120 -843
rect 1172 -895 1174 -843
rect 1118 -1161 1174 -895
rect 1118 -1213 1120 -1161
rect 1172 -1213 1174 -1161
rect 1118 -1479 1174 -1213
rect 1118 -1531 1120 -1479
rect 1172 -1531 1174 -1479
rect 1118 -1797 1174 -1531
rect 1118 -1849 1120 -1797
rect 1172 -1849 1174 -1797
rect 458 -2016 460 -1964
rect 512 -2016 514 -1964
rect 458 -2307 514 -2016
rect 1118 -1964 1174 -1849
rect 1118 -2016 1120 -1964
rect 1172 -2016 1174 -1964
rect 1118 -2022 1174 -2016
rect 458 -2359 460 -2307
rect 512 -2359 514 -2307
rect 458 -2365 514 -2359
use sky130_fd_pr__pfet_01v8_TMY429  XM1
timestamp 1730624594
transform 1 0 570 0 1 -886
box -246 -1173 246 1173
use sky130_fd_pr__nfet_01v8_XHGLWN  XM2
timestamp 1730624594
transform 1 0 1062 0 1 -1322
box -246 -737 246 737
<< labels >>
flabel metal1 324 -2155 420 -2059 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel metal1 324 -2279 420 -2183 0 FreeSans 320 0 0 0 vssa
port 4 nsew
flabel metal1 324 -2365 382 -2307 0 FreeSans 320 0 0 0 in
port 5 nsew
flabel via1 1036 -1930 1088 -1878 0 FreeSans 320 0 0 0 swn
port 3 nsew
flabel via1 544 -1930 596 -1878 0 FreeSans 320 0 0 0 swp
port 2 nsew
flabel via1 628 16 680 68 0 FreeSans 320 0 0 0 out
port 6 nsew
<< end >>
