magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect 315 -2043 349 -1967
rect 315 -2133 349 -2127
rect 701 -2043 735 -1967
rect 701 -2133 735 -2127
rect 1087 -2043 1121 -1967
rect 1087 -2133 1121 -2127
rect 1193 -2167 1227 -1967
rect 1193 -2257 1227 -2251
rect 1579 -2167 1613 -1967
rect 1579 -2257 1613 -2251
rect 1965 -2167 1999 -1967
rect 1965 -2257 1999 -2251
<< viali >>
rect 315 -2127 349 -2043
rect 701 -2127 735 -2043
rect 1087 -2127 1121 -2043
rect 1193 -2251 1227 -2167
rect 1579 -2251 1613 -2167
rect 1965 -2251 1999 -2167
<< metal1 >>
rect 479 128 499 180
rect 551 128 571 180
rect 865 128 885 180
rect 937 128 957 180
rect 409 38 415 90
rect 467 38 473 90
rect 409 -34 473 38
rect 409 -86 415 -34
rect 467 -86 473 -34
rect 409 -158 473 -86
rect 409 -210 415 -158
rect 467 -210 473 -158
rect 577 38 583 90
rect 635 38 801 90
rect 853 38 859 90
rect 577 -34 859 38
rect 577 -86 583 -34
rect 635 -86 801 -34
rect 853 -86 859 -34
rect 577 -158 859 -86
rect 577 -210 583 -158
rect 635 -210 801 -158
rect 853 -210 859 -158
rect 963 38 969 90
rect 1021 38 1027 90
rect 963 -34 1027 38
rect 963 -86 969 -34
rect 1021 -86 1027 -34
rect 963 -158 1027 -86
rect 963 -210 969 -158
rect 1021 -210 1027 -158
rect 479 -300 499 -248
rect 551 -300 571 -248
rect 865 -300 885 -248
rect 937 -300 957 -248
rect 479 -408 499 -356
rect 551 -408 571 -356
rect 865 -408 885 -356
rect 937 -408 957 -356
rect 409 -498 415 -446
rect 467 -498 473 -446
rect 409 -570 473 -498
rect 409 -622 415 -570
rect 467 -622 473 -570
rect 409 -694 473 -622
rect 409 -746 415 -694
rect 467 -746 473 -694
rect 577 -498 583 -446
rect 635 -498 801 -446
rect 853 -498 859 -446
rect 577 -570 859 -498
rect 577 -622 583 -570
rect 635 -622 801 -570
rect 853 -622 859 -570
rect 577 -694 859 -622
rect 577 -746 583 -694
rect 635 -746 801 -694
rect 853 -746 859 -694
rect 963 -498 969 -446
rect 1021 -498 1027 -446
rect 963 -570 1027 -498
rect 963 -622 969 -570
rect 1021 -622 1027 -570
rect 963 -694 1027 -622
rect 963 -746 969 -694
rect 1021 -746 1027 -694
rect 1357 -744 1377 -692
rect 1429 -744 1449 -692
rect 1743 -744 1763 -692
rect 1815 -744 1835 -692
rect 479 -836 499 -784
rect 551 -836 571 -784
rect 865 -836 885 -784
rect 937 -836 957 -784
rect 1287 -821 1351 -773
rect 1287 -873 1293 -821
rect 1345 -873 1351 -821
rect 1455 -821 1737 -773
rect 1455 -873 1461 -821
rect 1513 -873 1679 -821
rect 1731 -873 1737 -821
rect 1841 -821 1905 -773
rect 1841 -873 1847 -821
rect 1899 -873 1905 -821
rect 479 -944 499 -892
rect 551 -944 571 -892
rect 865 -944 885 -892
rect 937 -944 957 -892
rect 1357 -954 1377 -902
rect 1429 -954 1449 -902
rect 1743 -954 1763 -902
rect 1815 -954 1835 -902
rect 409 -1034 415 -982
rect 467 -1034 473 -982
rect 409 -1106 473 -1034
rect 409 -1158 415 -1106
rect 467 -1158 473 -1106
rect 409 -1230 473 -1158
rect 409 -1282 415 -1230
rect 467 -1282 473 -1230
rect 577 -1034 583 -982
rect 635 -1034 801 -982
rect 853 -1034 859 -982
rect 577 -1106 859 -1034
rect 577 -1158 583 -1106
rect 635 -1158 801 -1106
rect 853 -1158 859 -1106
rect 577 -1230 859 -1158
rect 577 -1282 583 -1230
rect 635 -1282 801 -1230
rect 853 -1282 859 -1230
rect 963 -1034 969 -982
rect 1021 -1034 1027 -982
rect 963 -1091 1027 -1034
rect 1357 -1062 1377 -1010
rect 1429 -1062 1449 -1010
rect 1743 -1062 1763 -1010
rect 1815 -1062 1835 -1010
rect 963 -1106 1351 -1091
rect 963 -1158 969 -1106
rect 1021 -1139 1351 -1106
rect 1021 -1158 1293 -1139
rect 963 -1191 1293 -1158
rect 1345 -1191 1351 -1139
rect 1455 -1139 1737 -1091
rect 1455 -1191 1461 -1139
rect 1513 -1191 1679 -1139
rect 1731 -1191 1737 -1139
rect 1841 -1139 1905 -1091
rect 1841 -1191 1847 -1139
rect 1899 -1191 1905 -1139
rect 963 -1230 1027 -1191
rect 963 -1282 969 -1230
rect 1021 -1282 1027 -1230
rect 1357 -1272 1377 -1220
rect 1429 -1272 1449 -1220
rect 1743 -1272 1763 -1220
rect 1815 -1272 1835 -1220
rect 479 -1372 499 -1320
rect 551 -1372 571 -1320
rect 865 -1372 885 -1320
rect 937 -1372 957 -1320
rect 1358 -1380 1377 -1328
rect 1429 -1380 1450 -1328
rect 1743 -1380 1763 -1328
rect 1815 -1380 1835 -1328
rect 479 -1480 499 -1428
rect 551 -1480 571 -1428
rect 865 -1480 885 -1428
rect 937 -1480 957 -1428
rect 1287 -1457 1351 -1409
rect 1287 -1509 1293 -1457
rect 1345 -1509 1351 -1457
rect 1455 -1457 1737 -1409
rect 1455 -1509 1461 -1457
rect 1513 -1509 1679 -1457
rect 1731 -1509 1737 -1457
rect 1841 -1457 1905 -1409
rect 1841 -1509 1847 -1457
rect 1899 -1509 1905 -1457
rect 409 -1570 415 -1518
rect 467 -1570 473 -1518
rect 409 -1642 473 -1570
rect 409 -1694 415 -1642
rect 467 -1694 473 -1642
rect 409 -1766 473 -1694
rect 409 -1818 415 -1766
rect 467 -1818 473 -1766
rect 577 -1570 583 -1518
rect 635 -1570 801 -1518
rect 853 -1570 859 -1518
rect 577 -1642 859 -1570
rect 577 -1694 583 -1642
rect 635 -1694 801 -1642
rect 853 -1694 859 -1642
rect 577 -1766 859 -1694
rect 577 -1818 583 -1766
rect 635 -1818 801 -1766
rect 853 -1818 859 -1766
rect 963 -1570 969 -1518
rect 1021 -1570 1027 -1518
rect 963 -1642 1027 -1570
rect 1357 -1590 1377 -1538
rect 1429 -1590 1449 -1538
rect 1743 -1590 1763 -1538
rect 1815 -1590 1835 -1538
rect 963 -1694 969 -1642
rect 1021 -1694 1027 -1642
rect 963 -1727 1027 -1694
rect 1357 -1698 1377 -1646
rect 1429 -1698 1449 -1646
rect 1742 -1698 1763 -1646
rect 1815 -1698 1834 -1646
rect 963 -1766 1351 -1727
rect 963 -1818 969 -1766
rect 1021 -1775 1351 -1766
rect 1021 -1818 1293 -1775
rect 963 -1827 1293 -1818
rect 1345 -1827 1351 -1775
rect 1455 -1775 1737 -1727
rect 1455 -1827 1461 -1775
rect 1513 -1827 1679 -1775
rect 1731 -1827 1737 -1775
rect 1841 -1775 1905 -1727
rect 1841 -1827 1847 -1775
rect 1899 -1827 1905 -1775
rect 479 -1908 499 -1856
rect 551 -1908 571 -1856
rect 865 -1908 885 -1856
rect 937 -1908 957 -1856
rect 1357 -1908 1377 -1856
rect 1429 -1908 1449 -1856
rect 1743 -1908 1763 -1856
rect 1815 -1908 1835 -1856
rect 493 -1988 499 -1936
rect 551 -1988 1763 -1936
rect 1815 -1988 1821 -1936
rect 279 -2043 415 -2037
rect 279 -2127 315 -2043
rect 349 -2127 415 -2043
rect 467 -2043 2035 -2037
rect 467 -2127 701 -2043
rect 735 -2127 1087 -2043
rect 1121 -2127 2035 -2043
rect 279 -2133 2035 -2127
rect 279 -2167 1847 -2161
rect 279 -2251 1193 -2167
rect 1227 -2251 1579 -2167
rect 1613 -2251 1847 -2167
rect 1899 -2167 2035 -2161
rect 1899 -2251 1965 -2167
rect 1999 -2251 2035 -2167
rect 279 -2257 2035 -2251
<< via1 >>
rect 499 128 551 180
rect 885 128 937 180
rect 415 38 467 90
rect 415 -86 467 -34
rect 415 -210 467 -158
rect 583 38 635 90
rect 801 38 853 90
rect 583 -86 635 -34
rect 801 -86 853 -34
rect 583 -210 635 -158
rect 801 -210 853 -158
rect 969 38 1021 90
rect 969 -86 1021 -34
rect 969 -210 1021 -158
rect 499 -300 551 -248
rect 885 -300 937 -248
rect 499 -408 551 -356
rect 885 -408 937 -356
rect 415 -498 467 -446
rect 415 -622 467 -570
rect 415 -746 467 -694
rect 583 -498 635 -446
rect 801 -498 853 -446
rect 583 -622 635 -570
rect 801 -622 853 -570
rect 583 -746 635 -694
rect 801 -746 853 -694
rect 969 -498 1021 -446
rect 969 -622 1021 -570
rect 969 -746 1021 -694
rect 1377 -744 1429 -692
rect 1763 -744 1815 -692
rect 499 -836 551 -784
rect 885 -836 937 -784
rect 1293 -873 1345 -821
rect 1461 -873 1513 -821
rect 1679 -873 1731 -821
rect 1847 -873 1899 -821
rect 499 -944 551 -892
rect 885 -944 937 -892
rect 1377 -954 1429 -902
rect 1763 -954 1815 -902
rect 415 -1034 467 -982
rect 415 -1158 467 -1106
rect 415 -1282 467 -1230
rect 583 -1034 635 -982
rect 801 -1034 853 -982
rect 583 -1158 635 -1106
rect 801 -1158 853 -1106
rect 583 -1282 635 -1230
rect 801 -1282 853 -1230
rect 969 -1034 1021 -982
rect 1377 -1062 1429 -1010
rect 1763 -1062 1815 -1010
rect 969 -1158 1021 -1106
rect 1293 -1191 1345 -1139
rect 1461 -1191 1513 -1139
rect 1679 -1191 1731 -1139
rect 1847 -1191 1899 -1139
rect 969 -1282 1021 -1230
rect 1377 -1272 1429 -1220
rect 1763 -1272 1815 -1220
rect 499 -1372 551 -1320
rect 885 -1372 937 -1320
rect 1377 -1380 1429 -1328
rect 1763 -1380 1815 -1328
rect 499 -1480 551 -1428
rect 885 -1480 937 -1428
rect 1293 -1509 1345 -1457
rect 1461 -1509 1513 -1457
rect 1679 -1509 1731 -1457
rect 1847 -1509 1899 -1457
rect 415 -1570 467 -1518
rect 415 -1694 467 -1642
rect 415 -1818 467 -1766
rect 583 -1570 635 -1518
rect 801 -1570 853 -1518
rect 583 -1694 635 -1642
rect 801 -1694 853 -1642
rect 583 -1818 635 -1766
rect 801 -1818 853 -1766
rect 969 -1570 1021 -1518
rect 1377 -1590 1429 -1538
rect 1763 -1590 1815 -1538
rect 969 -1694 1021 -1642
rect 1377 -1698 1429 -1646
rect 1763 -1698 1815 -1646
rect 969 -1818 1021 -1766
rect 1293 -1827 1345 -1775
rect 1461 -1827 1513 -1775
rect 1679 -1827 1731 -1775
rect 1847 -1827 1899 -1775
rect 499 -1908 551 -1856
rect 885 -1908 937 -1856
rect 1377 -1908 1429 -1856
rect 1763 -1908 1815 -1856
rect 499 -1988 551 -1936
rect 1763 -1988 1815 -1936
rect 415 -2127 467 -2037
rect 1847 -2251 1899 -2161
<< metal2 >>
rect 497 180 553 186
rect 497 128 499 180
rect 551 128 553 180
rect 413 90 469 96
rect 413 38 415 90
rect 467 38 469 90
rect 413 -34 469 38
rect 413 -86 415 -34
rect 467 -86 469 -34
rect 413 -158 469 -86
rect 413 -210 415 -158
rect 467 -210 469 -158
rect 413 -446 469 -210
rect 413 -498 415 -446
rect 467 -498 469 -446
rect 413 -570 469 -498
rect 413 -622 415 -570
rect 467 -622 469 -570
rect 413 -694 469 -622
rect 413 -746 415 -694
rect 467 -746 469 -694
rect 413 -982 469 -746
rect 413 -1034 415 -982
rect 467 -1034 469 -982
rect 413 -1106 469 -1034
rect 413 -1158 415 -1106
rect 467 -1158 469 -1106
rect 413 -1230 469 -1158
rect 413 -1282 415 -1230
rect 467 -1282 469 -1230
rect 413 -1518 469 -1282
rect 413 -1570 415 -1518
rect 467 -1570 469 -1518
rect 413 -1642 469 -1570
rect 413 -1694 415 -1642
rect 467 -1694 469 -1642
rect 413 -1766 469 -1694
rect 413 -1818 415 -1766
rect 467 -1818 469 -1766
rect 413 -2037 469 -1818
rect 497 -248 553 128
rect 883 180 939 186
rect 883 128 885 180
rect 937 128 939 180
rect 497 -300 499 -248
rect 551 -300 553 -248
rect 497 -356 553 -300
rect 497 -408 499 -356
rect 551 -408 553 -356
rect 497 -784 553 -408
rect 497 -836 499 -784
rect 551 -836 553 -784
rect 497 -892 553 -836
rect 497 -944 499 -892
rect 551 -944 553 -892
rect 497 -1320 553 -944
rect 497 -1372 499 -1320
rect 551 -1372 553 -1320
rect 497 -1428 553 -1372
rect 497 -1480 499 -1428
rect 551 -1480 553 -1428
rect 497 -1856 553 -1480
rect 581 90 637 96
rect 581 38 583 90
rect 635 38 637 90
rect 581 -34 637 38
rect 581 -86 583 -34
rect 635 -86 637 -34
rect 581 -158 637 -86
rect 581 -210 583 -158
rect 635 -210 637 -158
rect 581 -446 637 -210
rect 581 -498 583 -446
rect 635 -498 637 -446
rect 581 -570 637 -498
rect 581 -622 583 -570
rect 635 -622 637 -570
rect 581 -694 637 -622
rect 581 -746 583 -694
rect 635 -746 637 -694
rect 581 -982 637 -746
rect 581 -1034 583 -982
rect 635 -1034 637 -982
rect 581 -1106 637 -1034
rect 581 -1158 583 -1106
rect 635 -1158 637 -1106
rect 581 -1230 637 -1158
rect 581 -1282 583 -1230
rect 635 -1282 637 -1230
rect 581 -1518 637 -1282
rect 581 -1570 583 -1518
rect 635 -1570 637 -1518
rect 581 -1642 637 -1570
rect 581 -1694 583 -1642
rect 635 -1694 637 -1642
rect 581 -1766 637 -1694
rect 581 -1818 583 -1766
rect 635 -1818 637 -1766
rect 581 -1824 637 -1818
rect 799 90 855 96
rect 799 38 801 90
rect 853 38 855 90
rect 799 -34 855 38
rect 799 -86 801 -34
rect 853 -86 855 -34
rect 799 -158 855 -86
rect 799 -210 801 -158
rect 853 -210 855 -158
rect 799 -446 855 -210
rect 799 -498 801 -446
rect 853 -498 855 -446
rect 799 -570 855 -498
rect 799 -622 801 -570
rect 853 -622 855 -570
rect 799 -694 855 -622
rect 799 -746 801 -694
rect 853 -746 855 -694
rect 799 -982 855 -746
rect 799 -1034 801 -982
rect 853 -1034 855 -982
rect 799 -1106 855 -1034
rect 799 -1158 801 -1106
rect 853 -1158 855 -1106
rect 799 -1230 855 -1158
rect 799 -1282 801 -1230
rect 853 -1282 855 -1230
rect 799 -1518 855 -1282
rect 799 -1570 801 -1518
rect 853 -1570 855 -1518
rect 799 -1642 855 -1570
rect 799 -1694 801 -1642
rect 853 -1694 855 -1642
rect 799 -1766 855 -1694
rect 799 -1818 801 -1766
rect 853 -1818 855 -1766
rect 799 -1824 855 -1818
rect 883 -248 939 128
rect 883 -300 885 -248
rect 937 -300 939 -248
rect 883 -356 939 -300
rect 883 -408 885 -356
rect 937 -408 939 -356
rect 883 -784 939 -408
rect 883 -836 885 -784
rect 937 -836 939 -784
rect 883 -892 939 -836
rect 883 -944 885 -892
rect 937 -944 939 -892
rect 883 -1320 939 -944
rect 883 -1372 885 -1320
rect 937 -1372 939 -1320
rect 883 -1428 939 -1372
rect 883 -1480 885 -1428
rect 937 -1480 939 -1428
rect 497 -1908 499 -1856
rect 551 -1908 553 -1856
rect 497 -1936 553 -1908
rect 883 -1856 939 -1480
rect 967 90 1023 96
rect 967 38 969 90
rect 1021 38 1023 90
rect 967 -34 1023 38
rect 967 -86 969 -34
rect 1021 -86 1023 -34
rect 967 -158 1023 -86
rect 967 -210 969 -158
rect 1021 -210 1023 -158
rect 967 -446 1023 -210
rect 967 -498 969 -446
rect 1021 -498 1023 -446
rect 967 -570 1023 -498
rect 967 -622 969 -570
rect 1021 -622 1023 -570
rect 967 -694 1023 -622
rect 967 -746 969 -694
rect 1021 -746 1023 -694
rect 967 -982 1023 -746
rect 1375 -692 1431 -686
rect 1375 -744 1377 -692
rect 1429 -744 1431 -692
rect 967 -1034 969 -982
rect 1021 -1034 1023 -982
rect 967 -1106 1023 -1034
rect 967 -1158 969 -1106
rect 1021 -1158 1023 -1106
rect 967 -1230 1023 -1158
rect 967 -1282 969 -1230
rect 1021 -1282 1023 -1230
rect 967 -1518 1023 -1282
rect 967 -1570 969 -1518
rect 1021 -1570 1023 -1518
rect 967 -1642 1023 -1570
rect 967 -1694 969 -1642
rect 1021 -1694 1023 -1642
rect 967 -1766 1023 -1694
rect 967 -1818 969 -1766
rect 1021 -1818 1023 -1766
rect 967 -1824 1023 -1818
rect 1291 -821 1347 -767
rect 1291 -873 1293 -821
rect 1345 -873 1347 -821
rect 1291 -1139 1347 -873
rect 1291 -1191 1293 -1139
rect 1345 -1191 1347 -1139
rect 1291 -1457 1347 -1191
rect 1291 -1509 1293 -1457
rect 1345 -1509 1347 -1457
rect 1291 -1775 1347 -1509
rect 1291 -1827 1293 -1775
rect 1345 -1827 1347 -1775
rect 1291 -1833 1347 -1827
rect 1375 -902 1431 -744
rect 1761 -692 1817 -686
rect 1761 -744 1763 -692
rect 1815 -744 1817 -692
rect 1375 -954 1377 -902
rect 1429 -954 1431 -902
rect 1375 -1010 1431 -954
rect 1375 -1062 1377 -1010
rect 1429 -1062 1431 -1010
rect 1375 -1220 1431 -1062
rect 1375 -1272 1377 -1220
rect 1429 -1272 1431 -1220
rect 1375 -1328 1431 -1272
rect 1375 -1380 1377 -1328
rect 1429 -1380 1431 -1328
rect 1375 -1538 1431 -1380
rect 1375 -1590 1377 -1538
rect 1429 -1590 1431 -1538
rect 1375 -1646 1431 -1590
rect 1375 -1698 1377 -1646
rect 1429 -1698 1431 -1646
rect 883 -1908 885 -1856
rect 937 -1908 939 -1856
rect 883 -1914 939 -1908
rect 1375 -1856 1431 -1698
rect 1459 -821 1515 -767
rect 1459 -873 1461 -821
rect 1513 -873 1515 -821
rect 1459 -1139 1515 -873
rect 1459 -1191 1461 -1139
rect 1513 -1191 1515 -1139
rect 1459 -1457 1515 -1191
rect 1459 -1509 1461 -1457
rect 1513 -1509 1515 -1457
rect 1459 -1775 1515 -1509
rect 1459 -1827 1461 -1775
rect 1513 -1827 1515 -1775
rect 1459 -1833 1515 -1827
rect 1677 -821 1733 -767
rect 1677 -873 1679 -821
rect 1731 -873 1733 -821
rect 1677 -1139 1733 -873
rect 1677 -1191 1679 -1139
rect 1731 -1191 1733 -1139
rect 1677 -1457 1733 -1191
rect 1677 -1509 1679 -1457
rect 1731 -1509 1733 -1457
rect 1677 -1775 1733 -1509
rect 1677 -1827 1679 -1775
rect 1731 -1827 1733 -1775
rect 1677 -1833 1733 -1827
rect 1761 -902 1817 -744
rect 1761 -954 1763 -902
rect 1815 -954 1817 -902
rect 1761 -1010 1817 -954
rect 1761 -1062 1763 -1010
rect 1815 -1062 1817 -1010
rect 1761 -1220 1817 -1062
rect 1761 -1272 1763 -1220
rect 1815 -1272 1817 -1220
rect 1761 -1328 1817 -1272
rect 1761 -1380 1763 -1328
rect 1815 -1380 1817 -1328
rect 1761 -1538 1817 -1380
rect 1761 -1590 1763 -1538
rect 1815 -1590 1817 -1538
rect 1761 -1646 1817 -1590
rect 1761 -1698 1763 -1646
rect 1815 -1698 1817 -1646
rect 1375 -1908 1377 -1856
rect 1429 -1908 1431 -1856
rect 1375 -1914 1431 -1908
rect 1761 -1856 1817 -1698
rect 1761 -1908 1763 -1856
rect 1815 -1908 1817 -1856
rect 497 -1988 499 -1936
rect 551 -1988 553 -1936
rect 497 -1994 553 -1988
rect 1761 -1936 1817 -1908
rect 1761 -1988 1763 -1936
rect 1815 -1988 1817 -1936
rect 1761 -1994 1817 -1988
rect 1845 -821 1901 -767
rect 1845 -873 1847 -821
rect 1899 -873 1901 -821
rect 1845 -1139 1901 -873
rect 1845 -1191 1847 -1139
rect 1899 -1191 1901 -1139
rect 1845 -1457 1901 -1191
rect 1845 -1509 1847 -1457
rect 1899 -1509 1901 -1457
rect 1845 -1775 1901 -1509
rect 1845 -1827 1847 -1775
rect 1899 -1827 1901 -1775
rect 413 -2127 415 -2037
rect 467 -2127 469 -2037
rect 413 -2133 469 -2127
rect 1845 -2161 1901 -1827
rect 1845 -2251 1847 -2161
rect 1899 -2251 1901 -2161
rect 1845 -2257 1901 -2251
use sky130_fd_pr__pfet_01v8_TMY429  XM1
timestamp 1730624594
transform 1 0 525 0 1 -864
box -246 -1173 246 1173
use sky130_fd_pr__pfet_01v8_TMY429  XM2
timestamp 1730624594
transform 1 0 911 0 1 -864
box -246 -1173 246 1173
use sky130_fd_pr__nfet_01v8_XHGLWN  XM3
timestamp 1730624594
transform 1 0 1403 0 1 -1300
box -246 -737 246 737
use sky130_fd_pr__nfet_01v8_XHGLWN  XM4
timestamp 1730624594
transform 1 0 1789 0 1 -1300
box -246 -737 246 737
<< labels >>
flabel metal1 279 -2133 375 -2037 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel metal1 279 -2257 375 -2161 0 FreeSans 320 0 0 0 vssa
port 5 nsew
flabel via1 885 -1908 937 -1856 0 FreeSans 320 0 0 0 ckb
port 4 nsew
flabel via1 1377 -1908 1429 -1856 0 FreeSans 320 0 0 0 ck
port 3 nsew
flabel via1 1763 -744 1815 -692 0 FreeSans 320 0 0 0 in
port 2 nsew
flabel via1 969 38 1021 90 0 FreeSans 320 0 0 0 out
port 6 nsew
<< end >>
