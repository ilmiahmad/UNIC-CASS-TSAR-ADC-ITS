magic
tech sky130A
magscale 1 2
timestamp 1730612193
<< nwell >>
rect 11439 -2004 11665 -1778
rect 11162 -2840 11388 -2614
rect 1723 -3664 1949 -3438
<< pwell >>
rect -414 -2344 11406 -2248
rect -415 -3184 11168 -3088
<< psubdiff >>
rect -409 -2344 -385 -2310
rect 11425 -2344 11449 -2310
rect -410 -3184 -386 -3150
rect 11148 -3184 11172 -3150
rect 1953 -4024 1977 -3990
rect 3788 -4024 3812 -3990
<< nsubdiff >>
rect 11475 -1848 11535 -1814
rect 11569 -1848 11629 -1814
rect 11475 -1874 11509 -1848
rect 11475 -1934 11509 -1908
rect 11595 -1874 11629 -1848
rect 11595 -1934 11629 -1908
rect 11475 -1968 11535 -1934
rect 11569 -1968 11629 -1934
rect 11198 -2684 11258 -2650
rect 11292 -2684 11352 -2650
rect 11198 -2710 11232 -2684
rect 11198 -2770 11232 -2744
rect 11318 -2710 11352 -2684
rect 11318 -2770 11352 -2744
rect 11198 -2804 11258 -2770
rect 11292 -2804 11352 -2770
rect 1759 -3508 1819 -3474
rect 1853 -3508 1913 -3474
rect 1759 -3534 1793 -3508
rect 1759 -3594 1793 -3568
rect 1879 -3534 1913 -3508
rect 1879 -3594 1913 -3568
rect 1759 -3628 1819 -3594
rect 1853 -3628 1913 -3594
<< psubdiffcont >>
rect -385 -2344 11425 -2310
rect -386 -3184 11148 -3150
rect 1977 -4024 3788 -3990
<< nsubdiffcont >>
rect 11535 -1848 11569 -1814
rect 11475 -1908 11509 -1874
rect 11595 -1908 11629 -1874
rect 11535 -1968 11569 -1934
rect 11258 -2684 11292 -2650
rect 11198 -2744 11232 -2710
rect 11318 -2744 11352 -2710
rect 11258 -2804 11292 -2770
rect 1819 -3508 1853 -3474
rect 1759 -3568 1793 -3534
rect 1879 -3568 1913 -3534
rect 1819 -3628 1853 -3594
<< locali >>
rect 11475 -1848 11535 -1814
rect 11569 -1848 11629 -1814
rect 11475 -1874 11509 -1848
rect 11475 -1934 11509 -1908
rect 11595 -1874 11629 -1848
rect 11595 -1934 11629 -1908
rect 11475 -1968 11535 -1934
rect 11569 -1968 11629 -1934
rect -401 -2344 -385 -2310
rect 11425 -2344 11441 -2310
rect 11198 -2684 11258 -2650
rect 11292 -2684 11352 -2650
rect 11198 -2710 11232 -2684
rect 11198 -2770 11232 -2744
rect 11318 -2710 11352 -2684
rect 11318 -2770 11352 -2744
rect 11198 -2804 11258 -2770
rect 11292 -2804 11352 -2770
rect -402 -3184 -386 -3150
rect 11148 -3184 11164 -3150
rect 1759 -3508 1819 -3474
rect 1853 -3508 1913 -3474
rect 1759 -3534 1793 -3508
rect 1759 -3594 1793 -3568
rect 1879 -3534 1913 -3508
rect 1879 -3594 1913 -3568
rect 1759 -3628 1819 -3594
rect 1853 -3628 1913 -3594
rect 1961 -4024 1977 -3990
rect 3788 -4024 3804 -3990
<< viali >>
rect -385 -1769 -351 -1735
rect 1362 -1871 1396 -1837
rect 1820 -1871 1854 -1837
rect 3294 -1871 3328 -1837
rect 3752 -1871 3786 -1837
rect 5226 -1871 5260 -1837
rect 5684 -1871 5718 -1837
rect 7158 -1871 7192 -1837
rect 7616 -1871 7650 -1837
rect 9090 -1871 9124 -1837
rect 9548 -1871 9582 -1837
rect 11535 -1848 11569 -1814
rect -384 -2007 -350 -1973
rect 1548 -2007 1582 -1973
rect 3480 -2007 3514 -1973
rect 5412 -2007 5446 -1973
rect 7344 -2007 7378 -1973
rect 9276 -2007 9310 -1973
rect 11342 -2007 11376 -1973
rect 11033 -2081 11067 -2047
rect 11258 -2081 11292 -2047
rect -89 -2165 -55 -2131
rect 1067 -2143 1101 -2109
rect 2999 -2143 3033 -2109
rect 4931 -2143 4965 -2109
rect 6863 -2143 6897 -2109
rect 8795 -2143 8829 -2109
rect 10727 -2143 10761 -2109
rect -113 -2710 -79 -2676
rect 1361 -2711 1395 -2677
rect 1819 -2711 1853 -2677
rect 3293 -2711 3327 -2677
rect 3751 -2711 3785 -2677
rect 5225 -2711 5259 -2677
rect 5683 -2711 5717 -2677
rect 7157 -2711 7191 -2677
rect 7615 -2711 7649 -2677
rect 9089 -2711 9123 -2677
rect 9547 -2711 9581 -2677
rect 11258 -2684 11292 -2650
rect -385 -2847 -351 -2813
rect 1547 -2847 1581 -2813
rect 3479 -2847 3513 -2813
rect 5411 -2847 5445 -2813
rect 7343 -2847 7377 -2813
rect 9275 -2847 9309 -2813
rect 11021 -2847 11055 -2813
rect 1066 -2983 1100 -2949
rect 2998 -2983 3032 -2949
rect 4930 -2983 4964 -2949
rect 6862 -2983 6896 -2949
rect 8794 -2983 8828 -2949
rect 10726 -2983 10760 -2949
rect 1819 -3508 1853 -3474
rect 3705 -3687 3739 -3653
rect 2006 -3755 2040 -3721
rect 2114 -3755 2148 -3721
rect 2282 -3755 2316 -3721
rect 2650 -3755 2684 -3721
rect 2926 -3755 2960 -3721
rect 3478 -3755 3512 -3721
rect 3613 -3755 3647 -3721
<< metal1 >>
rect -769 -1735 11581 -1704
rect -769 -1769 -385 -1735
rect -351 -1769 11581 -1735
rect -769 -1800 11581 -1769
rect -769 -2544 -673 -1800
rect 11523 -1814 11581 -1800
rect 1350 -1837 1408 -1831
rect 1808 -1837 1866 -1831
rect 1350 -1871 1362 -1837
rect 1396 -1871 1820 -1837
rect 1854 -1871 1866 -1837
rect 1350 -1877 1408 -1871
rect 1808 -1877 1866 -1871
rect 3282 -1837 3340 -1831
rect 3740 -1837 3798 -1831
rect 3282 -1871 3294 -1837
rect 3328 -1871 3752 -1837
rect 3786 -1871 3798 -1837
rect 3282 -1877 3340 -1871
rect 3740 -1877 3798 -1871
rect 5214 -1837 5272 -1831
rect 5672 -1837 5730 -1831
rect 5214 -1871 5226 -1837
rect 5260 -1871 5684 -1837
rect 5718 -1871 5730 -1837
rect 5214 -1877 5272 -1871
rect 5672 -1877 5730 -1871
rect 7146 -1837 7204 -1831
rect 7604 -1837 7662 -1831
rect 7146 -1871 7158 -1837
rect 7192 -1871 7616 -1837
rect 7650 -1871 7662 -1837
rect 7146 -1877 7204 -1871
rect 7604 -1877 7662 -1871
rect 9078 -1837 9136 -1831
rect 9536 -1837 9594 -1831
rect 9078 -1871 9090 -1837
rect 9124 -1871 9548 -1837
rect 9582 -1871 9594 -1837
rect 11523 -1848 11535 -1814
rect 11569 -1848 11581 -1814
rect 11523 -1854 11581 -1848
rect 9078 -1877 9136 -1871
rect 9536 -1877 9594 -1871
rect -418 -2019 -408 -1967
rect -350 -2013 -338 -1967
rect -350 -2019 -340 -2013
rect 1514 -2019 1524 -1967
rect 1582 -2013 1594 -1967
rect 1582 -2019 1592 -2013
rect 3446 -2019 3456 -1967
rect 3514 -2013 3526 -1967
rect 3514 -2019 3524 -2013
rect 5378 -2019 5388 -1967
rect 5446 -2019 5458 -1967
rect 7310 -2019 7320 -1967
rect 7378 -2013 7390 -1967
rect 7378 -2019 7388 -2013
rect 9242 -2019 9252 -1967
rect 9310 -2019 9322 -1967
rect 11320 -2013 11330 -1961
rect 11388 -2013 11398 -1961
rect 11021 -2047 11079 -2041
rect 11246 -2047 11304 -2041
rect 11021 -2081 11033 -2047
rect 11067 -2081 11258 -2047
rect 11292 -2081 11304 -2047
rect 11021 -2087 11079 -2081
rect 11246 -2087 11304 -2081
rect 1045 -2109 1123 -2103
rect -111 -2177 -101 -2125
rect -43 -2177 -33 -2125
rect 1045 -2143 1067 -2109
rect 1101 -2143 1123 -2109
rect 1045 -2195 1055 -2143
rect 1113 -2195 1123 -2143
rect 2977 -2109 3055 -2103
rect 2977 -2143 2999 -2109
rect 3033 -2143 3055 -2109
rect 2977 -2195 2987 -2143
rect 3045 -2195 3055 -2143
rect 4909 -2109 4987 -2103
rect 4909 -2143 4931 -2109
rect 4965 -2143 4987 -2109
rect 4909 -2195 4919 -2143
rect 4977 -2195 4987 -2143
rect 6841 -2109 6919 -2103
rect 6841 -2143 6863 -2109
rect 6897 -2143 6919 -2109
rect 6841 -2195 6851 -2143
rect 6909 -2195 6919 -2143
rect 8773 -2109 8851 -2103
rect 8773 -2143 8795 -2109
rect 8829 -2143 8851 -2109
rect 8773 -2195 8783 -2143
rect 8841 -2195 8851 -2143
rect 10705 -2109 10783 -2103
rect 10705 -2143 10727 -2109
rect 10761 -2143 10783 -2109
rect 10705 -2195 10715 -2143
rect 10773 -2195 10783 -2143
rect -414 -2344 11778 -2248
rect -769 -2640 11453 -2544
rect -769 -3384 -673 -2640
rect 11246 -2650 11304 -2640
rect -135 -2720 -125 -2668
rect -67 -2720 -57 -2668
rect 1339 -2723 1349 -2671
rect 1407 -2677 1417 -2671
rect 1807 -2677 1865 -2671
rect 1407 -2711 1819 -2677
rect 1853 -2711 1865 -2677
rect 1407 -2723 1417 -2711
rect 1807 -2717 1865 -2711
rect 3281 -2677 3339 -2671
rect 3739 -2677 3797 -2671
rect 3281 -2711 3293 -2677
rect 3327 -2711 3751 -2677
rect 3785 -2711 3797 -2677
rect 3281 -2717 3339 -2711
rect 3739 -2717 3797 -2711
rect 5213 -2677 5271 -2671
rect 5671 -2677 5729 -2671
rect 5213 -2711 5225 -2677
rect 5259 -2711 5683 -2677
rect 5717 -2711 5729 -2677
rect 5213 -2717 5271 -2711
rect 5671 -2717 5729 -2711
rect 7145 -2677 7203 -2671
rect 7603 -2677 7661 -2671
rect 7145 -2711 7157 -2677
rect 7191 -2711 7615 -2677
rect 7649 -2711 7661 -2677
rect 7145 -2717 7203 -2711
rect 7603 -2717 7661 -2711
rect 9077 -2677 9135 -2671
rect 9535 -2677 9593 -2671
rect 9077 -2711 9089 -2677
rect 9123 -2711 9547 -2677
rect 9581 -2711 9593 -2677
rect 11246 -2684 11258 -2650
rect 11292 -2684 11304 -2650
rect 11246 -2690 11304 -2684
rect 9077 -2717 9135 -2711
rect 9535 -2717 9593 -2711
rect -407 -2859 -397 -2807
rect -339 -2859 -329 -2807
rect 1525 -2859 1535 -2807
rect 1593 -2859 1603 -2807
rect 3457 -2859 3467 -2807
rect 3525 -2859 3535 -2807
rect 5389 -2859 5399 -2807
rect 5457 -2859 5467 -2807
rect 7321 -2859 7331 -2807
rect 7389 -2859 7399 -2807
rect 9253 -2859 9263 -2807
rect 9321 -2859 9331 -2807
rect 10999 -2859 11009 -2807
rect 11067 -2859 11077 -2807
rect 1044 -2995 1054 -2943
rect 1112 -2995 1122 -2943
rect 2976 -2995 2986 -2943
rect 3044 -2995 3054 -2943
rect 4908 -2995 4918 -2943
rect 4976 -2995 4986 -2943
rect 6840 -2995 6850 -2943
rect 6908 -2995 6918 -2943
rect 8772 -2995 8782 -2943
rect 8840 -2995 8850 -2943
rect 10704 -2995 10714 -2943
rect 10772 -2995 10782 -2943
rect 11682 -3088 11778 -2344
rect -415 -3184 11778 -3088
rect -769 -3474 11453 -3384
rect -769 -3480 1819 -3474
rect 1807 -3508 1819 -3480
rect 1853 -3480 11453 -3474
rect 1853 -3508 1865 -3480
rect 1807 -3514 1865 -3508
rect 3683 -3699 3693 -3647
rect 3751 -3699 3761 -3647
rect 1984 -3761 1994 -3709
rect 2052 -3761 2062 -3709
rect 2102 -3721 2160 -3715
rect 2270 -3721 2328 -3715
rect 2102 -3755 2114 -3721
rect 2148 -3755 2282 -3721
rect 2316 -3755 2328 -3721
rect 2102 -3761 2160 -3755
rect 2270 -3761 2328 -3755
rect 2638 -3721 2696 -3715
rect 2914 -3721 2972 -3715
rect 2638 -3755 2650 -3721
rect 2684 -3755 2926 -3721
rect 2960 -3755 2972 -3721
rect 2638 -3761 2696 -3755
rect 2914 -3761 2972 -3755
rect 3456 -3721 3534 -3715
rect 3601 -3721 3659 -3715
rect 3456 -3755 3478 -3721
rect 3512 -3755 3613 -3721
rect 3647 -3755 3659 -3721
rect 3456 -3767 3534 -3755
rect 3601 -3761 3659 -3755
rect 3456 -3819 3466 -3767
rect 3524 -3819 3534 -3767
rect 11682 -3928 11778 -3184
rect -770 -4024 11778 -3928
<< via1 >>
rect -408 -1973 -350 -1967
rect -408 -2007 -384 -1973
rect -384 -2007 -350 -1973
rect -408 -2019 -350 -2007
rect 1524 -1973 1582 -1967
rect 1524 -2007 1548 -1973
rect 1548 -2007 1582 -1973
rect 1524 -2019 1582 -2007
rect 3456 -1973 3514 -1967
rect 3456 -2007 3480 -1973
rect 3480 -2007 3514 -1973
rect 3456 -2019 3514 -2007
rect 5388 -1973 5446 -1967
rect 5388 -2007 5412 -1973
rect 5412 -2007 5446 -1973
rect 5388 -2019 5446 -2007
rect 7320 -1973 7378 -1967
rect 7320 -2007 7344 -1973
rect 7344 -2007 7378 -1973
rect 7320 -2019 7378 -2007
rect 9252 -1973 9310 -1967
rect 9252 -2007 9276 -1973
rect 9276 -2007 9310 -1973
rect 9252 -2019 9310 -2007
rect 11330 -1973 11388 -1961
rect 11330 -2007 11342 -1973
rect 11342 -2007 11376 -1973
rect 11376 -2007 11388 -1973
rect 11330 -2013 11388 -2007
rect -101 -2131 -43 -2125
rect -101 -2165 -89 -2131
rect -89 -2165 -55 -2131
rect -55 -2165 -43 -2131
rect -101 -2177 -43 -2165
rect 1055 -2195 1113 -2143
rect 2987 -2195 3045 -2143
rect 4919 -2195 4977 -2143
rect 6851 -2195 6909 -2143
rect 8783 -2195 8841 -2143
rect 10715 -2195 10773 -2143
rect -125 -2676 -67 -2668
rect -125 -2710 -113 -2676
rect -113 -2710 -79 -2676
rect -79 -2710 -67 -2676
rect -125 -2720 -67 -2710
rect 1349 -2677 1407 -2671
rect 1349 -2711 1361 -2677
rect 1361 -2711 1395 -2677
rect 1395 -2711 1407 -2677
rect 1349 -2723 1407 -2711
rect -397 -2813 -339 -2807
rect -397 -2847 -385 -2813
rect -385 -2847 -351 -2813
rect -351 -2847 -339 -2813
rect -397 -2859 -339 -2847
rect 1535 -2813 1593 -2807
rect 1535 -2847 1547 -2813
rect 1547 -2847 1581 -2813
rect 1581 -2847 1593 -2813
rect 1535 -2859 1593 -2847
rect 3467 -2813 3525 -2807
rect 3467 -2847 3479 -2813
rect 3479 -2847 3513 -2813
rect 3513 -2847 3525 -2813
rect 3467 -2859 3525 -2847
rect 5399 -2813 5457 -2807
rect 5399 -2847 5411 -2813
rect 5411 -2847 5445 -2813
rect 5445 -2847 5457 -2813
rect 5399 -2859 5457 -2847
rect 7331 -2813 7389 -2807
rect 7331 -2847 7343 -2813
rect 7343 -2847 7377 -2813
rect 7377 -2847 7389 -2813
rect 7331 -2859 7389 -2847
rect 9263 -2813 9321 -2807
rect 9263 -2847 9275 -2813
rect 9275 -2847 9309 -2813
rect 9309 -2847 9321 -2813
rect 9263 -2859 9321 -2847
rect 11009 -2813 11067 -2807
rect 11009 -2847 11021 -2813
rect 11021 -2847 11055 -2813
rect 11055 -2847 11067 -2813
rect 11009 -2859 11067 -2847
rect 1054 -2949 1112 -2943
rect 1054 -2983 1066 -2949
rect 1066 -2983 1100 -2949
rect 1100 -2983 1112 -2949
rect 1054 -2995 1112 -2983
rect 2986 -2949 3044 -2943
rect 2986 -2983 2998 -2949
rect 2998 -2983 3032 -2949
rect 3032 -2983 3044 -2949
rect 2986 -2995 3044 -2983
rect 4918 -2949 4976 -2943
rect 4918 -2983 4930 -2949
rect 4930 -2983 4964 -2949
rect 4964 -2983 4976 -2949
rect 4918 -2995 4976 -2983
rect 6850 -2949 6908 -2943
rect 6850 -2983 6862 -2949
rect 6862 -2983 6896 -2949
rect 6896 -2983 6908 -2949
rect 6850 -2995 6908 -2983
rect 8782 -2949 8840 -2943
rect 8782 -2983 8794 -2949
rect 8794 -2983 8828 -2949
rect 8828 -2983 8840 -2949
rect 8782 -2995 8840 -2983
rect 10714 -2949 10772 -2943
rect 10714 -2983 10726 -2949
rect 10726 -2983 10760 -2949
rect 10760 -2983 10772 -2949
rect 10714 -2995 10772 -2983
rect 3693 -3653 3751 -3647
rect 3693 -3687 3705 -3653
rect 3705 -3687 3739 -3653
rect 3739 -3687 3751 -3653
rect 3693 -3699 3751 -3687
rect 1994 -3721 2052 -3709
rect 1994 -3755 2006 -3721
rect 2006 -3755 2040 -3721
rect 2040 -3755 2052 -3721
rect 1994 -3761 2052 -3755
rect 3466 -3819 3524 -3767
<< metal2 >>
rect -418 -1957 -340 -1947
rect 11320 -1951 11398 -1941
rect 1524 -1967 1582 -1957
rect 3456 -1967 3514 -1957
rect 5388 -1967 5446 -1957
rect 7320 -1967 7378 -1957
rect 9252 -1967 9310 -1957
rect -340 -2019 1524 -1967
rect 1582 -2019 3456 -1967
rect 3514 -2019 5388 -1967
rect 5446 -2019 7320 -1967
rect 7378 -2019 9252 -1967
rect 1524 -2029 1582 -2019
rect 3456 -2029 3514 -2019
rect 5388 -2029 5446 -2019
rect 7320 -2029 7378 -2019
rect 9252 -2029 9310 -2019
rect -418 -2039 -340 -2029
rect 11320 -2033 11398 -2023
rect -111 -2115 -33 -2105
rect 10705 -2133 10783 -2123
rect -111 -2197 -33 -2187
rect 1055 -2143 1113 -2133
rect 2987 -2143 3045 -2133
rect 4919 -2143 4977 -2133
rect 6851 -2143 6909 -2133
rect 8783 -2143 8841 -2133
rect 1113 -2195 2987 -2143
rect 3045 -2195 4919 -2143
rect 4977 -2195 6851 -2143
rect 6909 -2195 8783 -2143
rect 8841 -2195 10705 -2143
rect 1055 -2205 1113 -2195
rect 2987 -2205 3045 -2195
rect 4919 -2205 4977 -2195
rect 6851 -2205 6909 -2195
rect 8783 -2205 8841 -2195
rect 10705 -2215 10783 -2205
rect -135 -2436 -57 -2426
rect 11320 -2436 11398 -2426
rect -57 -2508 11320 -2436
rect -135 -2518 -57 -2508
rect 11320 -2518 11398 -2508
rect -135 -2658 -57 -2648
rect -135 -2740 -57 -2730
rect 1339 -2661 1417 -2651
rect 1339 -2743 1417 -2733
rect -407 -2797 -329 -2787
rect 11509 -2797 11587 -2787
rect 1535 -2807 1593 -2797
rect 3467 -2807 3525 -2797
rect 5399 -2807 5457 -2797
rect 7331 -2807 7389 -2797
rect 9263 -2807 9321 -2797
rect -884 -2859 -407 -2807
rect -329 -2859 1535 -2807
rect 1593 -2859 3467 -2807
rect 3525 -2859 5399 -2807
rect 5457 -2859 7331 -2807
rect 7389 -2859 9263 -2807
rect 1535 -2869 1593 -2859
rect 3467 -2869 3525 -2859
rect 5399 -2869 5457 -2859
rect 7331 -2869 7389 -2859
rect 9263 -2869 9321 -2859
rect 11009 -2807 11067 -2797
rect 11067 -2859 11509 -2807
rect 11009 -2869 11067 -2859
rect -407 -2879 -329 -2869
rect 11509 -2879 11587 -2869
rect 10704 -2933 10782 -2923
rect 1054 -2943 1112 -2933
rect 2986 -2943 3044 -2933
rect 4918 -2943 4976 -2933
rect 6850 -2943 6908 -2933
rect 8782 -2943 8840 -2933
rect -884 -2995 1054 -2943
rect 1112 -2995 2986 -2943
rect 3044 -2995 4918 -2943
rect 4976 -2995 6850 -2943
rect 6908 -2995 8782 -2943
rect 8840 -2995 10704 -2943
rect 1054 -3005 1112 -2995
rect 2986 -3005 3044 -2995
rect 4918 -3005 4976 -2995
rect 6850 -3005 6908 -2995
rect 8782 -3005 8840 -2995
rect 10704 -3015 10782 -3005
rect 3693 -3647 3751 -3637
rect 1339 -3698 1417 -3688
rect 3751 -3699 4084 -3647
rect 1994 -3709 2052 -3699
rect 3693 -3709 3751 -3699
rect 1417 -3761 1994 -3709
rect 1994 -3771 2052 -3761
rect 3466 -3767 3524 -3757
rect 1339 -3781 1417 -3771
rect 3524 -3819 4084 -3767
rect 3466 -3829 3524 -3819
<< via2 >>
rect -418 -1967 -340 -1957
rect -418 -2019 -408 -1967
rect -408 -2019 -350 -1967
rect -350 -2019 -340 -1967
rect -418 -2029 -340 -2019
rect 11320 -1961 11398 -1951
rect 11320 -2013 11330 -1961
rect 11330 -2013 11388 -1961
rect 11388 -2013 11398 -1961
rect 11320 -2023 11398 -2013
rect -111 -2125 -33 -2115
rect -111 -2177 -101 -2125
rect -101 -2177 -43 -2125
rect -43 -2177 -33 -2125
rect -111 -2187 -33 -2177
rect 10705 -2143 10783 -2133
rect 10705 -2195 10715 -2143
rect 10715 -2195 10773 -2143
rect 10773 -2195 10783 -2143
rect 10705 -2205 10783 -2195
rect -135 -2508 -57 -2436
rect 11320 -2508 11398 -2436
rect -135 -2668 -57 -2658
rect -135 -2720 -125 -2668
rect -125 -2720 -67 -2668
rect -67 -2720 -57 -2668
rect -135 -2730 -57 -2720
rect 1339 -2671 1417 -2661
rect 1339 -2723 1349 -2671
rect 1349 -2723 1407 -2671
rect 1407 -2723 1417 -2671
rect 1339 -2733 1417 -2723
rect -407 -2807 -329 -2797
rect -407 -2859 -397 -2807
rect -397 -2859 -339 -2807
rect -339 -2859 -329 -2807
rect -407 -2869 -329 -2859
rect 11509 -2869 11587 -2797
rect 10704 -2943 10782 -2933
rect 10704 -2995 10714 -2943
rect 10714 -2995 10772 -2943
rect 10772 -2995 10782 -2943
rect 10704 -3005 10782 -2995
rect 1339 -3771 1417 -3698
<< metal3 >>
rect 11310 -1951 11408 -1946
rect -428 -1957 -330 -1952
rect -428 -2029 -418 -1957
rect -340 -2029 -330 -1957
rect 11310 -2023 11320 -1951
rect 11398 -2023 11408 -1951
rect 11310 -2028 11408 -2023
rect -428 -2034 -330 -2029
rect -407 -2792 -340 -2034
rect -121 -2115 -23 -2110
rect -121 -2187 -111 -2115
rect -33 -2187 -23 -2115
rect -121 -2192 -23 -2187
rect 10695 -2133 10793 -2128
rect -111 -2295 -33 -2192
rect 10695 -2205 10705 -2133
rect 10783 -2205 10793 -2133
rect 10695 -2210 10793 -2205
rect -121 -2367 -111 -2295
rect -33 -2367 -23 -2295
rect -145 -2436 -47 -2431
rect -145 -2508 -135 -2436
rect -57 -2508 -47 -2436
rect -145 -2513 -47 -2508
rect -135 -2653 -57 -2513
rect -145 -2658 -47 -2653
rect -145 -2730 -135 -2658
rect -57 -2730 -47 -2658
rect -145 -2735 -47 -2730
rect 1329 -2661 1427 -2656
rect 1329 -2733 1339 -2661
rect 1417 -2733 1427 -2661
rect 1329 -2738 1427 -2733
rect -417 -2797 -319 -2792
rect -417 -2869 -407 -2797
rect -329 -2869 -319 -2797
rect -417 -2874 -319 -2869
rect 1339 -3693 1417 -2738
rect 10704 -2928 10783 -2210
rect 11320 -2431 11398 -2028
rect 11310 -2436 11408 -2431
rect 11310 -2508 11320 -2436
rect 11398 -2508 11408 -2436
rect 11499 -2437 11509 -2365
rect 11587 -2437 11597 -2365
rect 11310 -2513 11408 -2508
rect 11509 -2792 11587 -2437
rect 11499 -2797 11597 -2792
rect 11499 -2869 11509 -2797
rect 11587 -2869 11597 -2797
rect 11499 -2874 11597 -2869
rect 10694 -2933 10792 -2928
rect 10694 -3005 10704 -2933
rect 10782 -3005 10792 -2933
rect 10694 -3010 10792 -3005
rect 1329 -3698 1427 -3693
rect 1329 -3771 1339 -3698
rect 1417 -3771 1427 -3698
rect 1329 -3776 1427 -3771
<< via3 >>
rect -111 -2367 -33 -2295
rect 11509 -2437 11587 -2365
<< metal4 >>
rect -111 -2294 -33 -2293
rect -112 -2295 -32 -2294
rect -112 -2367 -111 -2295
rect -33 -2365 -32 -2295
rect 11508 -2365 11588 -2364
rect -33 -2367 11509 -2365
rect -112 -2368 11509 -2367
rect -111 -2437 11509 -2368
rect 11587 -2437 11588 -2365
rect 11508 -2438 11588 -2437
use sky130_fd_sc_hd__dfrtp_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform 1 0 1518 0 1 -2296
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2
timestamp 1730246015
transform 1 0 3450 0 1 -2296
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3
timestamp 1730246015
transform 1 0 5382 0 1 -2296
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform 1 0 11178 0 1 -2296
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  x5
timestamp 1730246015
transform 1 0 7314 0 1 -2296
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x7
timestamp 1730246015
transform 1 0 -414 0 1 -2296
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x11
timestamp 1730246015
transform 1 0 9246 0 1 -2296
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x12
timestamp 1730246015
transform 1 0 -415 0 1 -3136
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x13
timestamp 1730246015
transform 1 0 1517 0 1 -3136
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x14
timestamp 1730246015
transform 1 0 3449 0 1 -3136
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x15
timestamp 1730246015
transform 1 0 5381 0 1 -3136
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x16
timestamp 1730246015
transform 1 0 7313 0 1 -3136
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x21
timestamp 1730246015
transform 1 0 9245 0 1 -3136
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  x22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform 1 0 1977 0 1 -3976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform 1 0 2253 0 1 -3976
box -38 -48 498 592
use sky130_fd_sc_hd__inv_8  x24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform 1 0 2713 0 1 -3976
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  x25
timestamp 1730246015
transform 1 0 3541 0 1 -3976
box -38 -48 314 592
<< labels >>
flabel metal2 4055 -3687 4080 -3661 0 FreeSans 800 0 0 0 CLKSB
port 1 nsew
flabel metal2 4050 -3806 4076 -3781 0 FreeSans 800 0 0 0 CLKS
port 3 nsew
flabel metal2 -873 -2854 -845 -2819 0 FreeSans 800 0 0 0 CKC
port 4 nsew
flabel metal2 -870 -2983 -854 -2953 0 FreeSans 800 0 0 0 RST
port 11 nsew
flabel metal1 -744 -3999 -707 -3959 0 FreeSans 800 0 0 0 VSSD
port 12 nsew
flabel metal1 -733 -1771 -696 -1731 0 FreeSans 800 0 0 0 VDDD
port 14 nsew
<< end >>
