* PEX produced on Rab 06 Nov 2024 10:28:37  CST using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from sar.ext - technology: sky130A

.subckt sar CF[0] CF[1] CF[2] CF[3] CF[4] CF[5] CF[6] CF[7] CF[8] CF[9] CKO CLK CLKS
+ CLKSB COMP_N COMP_P DOUT[0] DOUT[1] DOUT[2] DOUT[3] DOUT[4] DOUT[5] DOUT[6] DOUT[7]
+ DOUT[8] DOUT[9] EN SWN[0] SWN[1] SWN[2] SWN[3] SWN[4] SWN[5] SWN[6] SWN[7] SWN[8]
+ SWN[9] SWP[0] SWP[1] SWP[2] SWP[3] SWP[4] SWP[5] SWP[6] SWP[7] SWP[8] SWP[9] VDDD
+ VSSD
X0 a_1835_9813.t1 a_2122_10091.t4 VDDD.t1358 VDDD.t1357 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1 VSSD.t722 a_4739_10625.t2 a_4700_10499.t1 VSSD.t721 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VDDD.t1179 a_6077_9813.t8 clknet_1_1__leaf_CLK.t15 VDDD.t1178 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VSSD.t914 a_5515_4159.t3 a_5449_4233.t1 VSSD.t913 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4 VDDD.t477 VSSD.t1852 VDDD.t476 VDDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5 a_10373_5487.t0 a_10329_5729.t4 a_10207_5487.t0 VSSD.t452 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X6 a_5515_4159.t1 CLKS.t16 VDDD.t284 VDDD.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VSSD.t1568 VDDD.t1979 VSSD.t1567 VSSD.t1566 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8 a_4463_8893.t1 CF[0].t4 VSSD.t1584 VSSD.t1583 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VDDD.t14 a_10667_9813.t3 a_10654_10205.t1 VDDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_4425_3861.t0 a_4259_3861.t2 VDDD.t826 VDDD.t825 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 a_3210_10927.t1 EN.t0 VSSD.t880 VSSD.t879 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X12 a_5037_4221.t1 a_4993_3829.t4 a_4871_4233.t0 VSSD.t1105 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X13 VDDD.t634 a_8008_10927.t4 a_8183_10901.t1 VDDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 VDDD.t1497 CLK.t0 a_6813_7093.t3 VDDD.t1496 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 VSSD.t1565 VDDD.t1980 VSSD.t1564 VSSD.t1563 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X16 a_2710_6031.t3 a_2584_6147.t2 a_2306_6163.t3 VSSD.t775 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X17 a_7321_6575.t0 a_6942_6941.t4 a_7249_6575.t0 VSSD.t499 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 CF[6].t1 a_10667_5247.t3 VDDD.t1343 VDDD.t1342 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X19 VSSD.t95 clknet_1_1__leaf_CLK.t32 a_8951_10927.t1 VSSD.t94 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 VSSD.t705 a_2411_4917.t4 a_2342_4943.t2 VSSD.t704 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X21 a_7331_9269.t5 COMP_N.t0 VSSD.t421 VSSD.t420 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 a_4619_4636.t0 a_4424_4667.t2 a_4929_4399.t0 VSSD.t706 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X23 a_5015_3009.t0 CF[4].t4 VDDD.t798 VDDD.t797 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 VDDD.t1187 a_4463_4541.t2 a_4424_4667.t0 VDDD.t1186 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X25 VDDD.t562 a_10207_10901.t3 a_10194_11293.t0 VDDD.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 a_6251_6549.t2 a_6538_6827.t4 VDDD.t655 VDDD.t654 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X27 a_4146_6827.t1 a_4424_6843.t2 a_4380_6941.t0 VDDD.t843 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 a_2905_4399.t0 a_2526_4765.t4 a_2833_4399.t0 VSSD.t935 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X29 a_2623_6273.t1 CF[8].t4 VSSD.t1637 VSSD.t1636 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X30 VSSD.t568 a_3031_10901.t3 a_2965_10927.t1 VSSD.t567 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X31 a_6541_8213.t1 a_6375_8213.t2 VSSD.t698 VSSD.t697 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X32 VDDD.t956 a_10943_6549.t3 CF[9].t1 VDDD.t955 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X33 a_2397_4399.t0 a_1835_4373.t3 VSSD.t332 VSSD.t331 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X34 a_6077_9813.t4 clknet_0_CLK.t32 VSSD.t462 VSSD.t461 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 a_5576_3677.t1 a_5055_3285.t3 VDDD.t1191 VDDD.t1190 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X36 VDDD.t1469 CF[2].t4 a_6743_4399.t0 VDDD.t1468 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X37 VSSD.t1562 VDDD.t1981 VSSD.t1561 VSSD.t1479 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X38 VDDD.t480 VSSD.t1853 VDDD.t479 VDDD.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X39 VDDD.t483 VSSD.t1854 VDDD.t482 VDDD.t481 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X40 a_5147_11989.t1 a_4972_12015.t4 a_5326_12015.t1 VSSD.t1155 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X41 a_4146_4651.t0 a_4463_4541.t3 a_4421_4399.t0 VSSD.t831 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X42 SWN[9].t3 a_3583_4917.t3 VSSD.t403 VSSD.t402 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X43 a_8638_4221.t0 CLKS.t17 VSSD.t233 VSSD.t232 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X44 a_10759_6335.t0 CLKS.t18 VDDD.t286 VDDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X45 a_4527_8181.t0 a_4371_8449.t2 a_4672_8207.t1 VDDD.t1939 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X46 VSSD.t417 a_10207_10901.t4 x2/net11.t3 VSSD.t416 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X47 VDDD.t486 VSSD.t1855 VDDD.t485 VDDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X48 VDDD.t489 VSSD.t1856 VDDD.t488 VDDD.t487 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X49 VSSD.t53 clknet_1_0__leaf_CLK.t32 a_9595_3311.t1 VSSD.t52 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X50 a_10203_6575.t1 a_9853_6575.t2 a_10108_6575.t0 VDDD.t1882 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X51 VDDD.t136 clknet_1_1__leaf_CLK.t33 a_8951_10927.t0 VDDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X52 a_10299_7423.t2 EN.t1 VDDD.t1226 VDDD.t1225 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X53 a_7494_2767.t2 a_7407_3009.t2 a_7090_2899.t3 VDDD.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X54 VDDD.t492 VSSD.t1857 VDDD.t491 VDDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X55 a_10676_3311.t1 a_9761_3311.t2 a_10329_3553.t0 VSSD.t855 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X56 a_9117_7663.t0 a_8951_7663.t2 VDDD.t1700 VDDD.t1699 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X57 a_3158_10205.t3 a_2400_10107.t2 a_2595_10076.t1 VDDD.t1532 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X58 a_7824_4399.t2 a_6743_4399.t2 a_7477_4641.t3 VDDD.t1537 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X59 VSSD.t1560 VDDD.t1982 VSSD.t1559 VSSD.t1558 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X60 SWP[3].t1 a_8459_4159.t3 VDDD.t246 VDDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X61 VDDD.t288 CLKS.t19 a_3859_8725.t0 VDDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X62 a_8275_6335.t0 CLKS.t20 VDDD.t290 VDDD.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X63 DOUT[4].t3 a_10207_7637.t3 VSSD.t948 VSSD.t947 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X64 VSSD.t1557 VDDD.t1983 VSSD.t1556 VSSD.t1555 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X65 VDDD.t1946 a_5515_4159.t4 a_5502_3855.t1 VDDD.t1945 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X66 a_10311_6941.t0 a_9687_6575.t2 a_10203_6575.t2 VDDD.t852 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X67 SWN[4].t3 a_4043_7637.t3 VSSD.t870 VSSD.t869 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X68 a_9577_4949.t0 a_9411_4949.t2 VDDD.t1457 VDDD.t1456 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X69 a_6855_6717.t0 CF[1].t4 VDDD.t570 VDDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X70 VSSD.t1554 VDDD.t1984 VSSD.t1553 VSSD.t1459 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X71 VSSD.t820 a_6077_9813.t9 clknet_1_1__leaf_CLK.t31 VSSD.t819 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X72 VSSD.t846 a_8435_8181.t6 x3/COMP_BUF_P.t15 VSSD.t845 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X73 VDDD.t754 a_7563_2741.t4 a_7494_2767.t0 VDDD.t753 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X74 VDDD.t357 a_10032_7663.t4 a_10207_7637.t0 VDDD.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X75 a_2158_8207.t1 a_2032_8323.t2 a_1754_8339.t2 VSSD.t549 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X76 VDDD.t1976 a_7654_4943.t8 clknet_1_0__leaf_CLK.t29 VDDD.t1975 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X77 a_4421_6575.t0 a_3859_6549.t3 VSSD.t812 VSSD.t811 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X78 a_6891_8585.t2 a_6541_8213.t2 a_6796_8573.t1 VDDD.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X79 a_7125_8751.t0 a_7090_9003.t4 a_6803_8725.t0 VSSD.t463 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X80 a_2309_10389.t0 a_2143_10389.t2 VDDD.t546 VDDD.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X81 VDDD.t495 VSSD.t1858 VDDD.t494 VDDD.t493 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X82 VDDD.t62 CF[3].t4 a_8126_2767.t0 VDDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X83 a_7348_10927.t1 x2/net3.t4 VSSD.t130 VSSD.t129 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X84 VSSD.t1851 a_7654_4943.t9 clknet_1_0__leaf_CLK.t30 VSSD.t1850 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X85 VSSD.t1552 VDDD.t1985 VSSD.t1551 VSSD.t1550 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X86 x2/net9.t1 a_3031_10901.t4 VDDD.t790 VDDD.t789 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X87 VDDD.t68 a_4411_6005.t3 SWN[2].t1 VDDD.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X88 VSSD.t1549 VDDD.t1986 VSSD.t1548 VSSD.t1547 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X89 VDDD.t292 CLKS.t21 a_5055_3285.t2 VDDD.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X90 a_2965_10927.t0 a_1775_10927.t2 a_2856_10927.t3 VSSD.t430 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X91 a_2840_11837.t1 x2/net9.t4 VDDD.t1177 VDDD.t1176 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X92 a_4653_5309.t0 a_4274_4943.t4 a_4581_5309.t1 VSSD.t613 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X93 VDDD.t1705 a_1651_4917.t3 SWP[8].t1 VDDD.t1704 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X94 VDDD.t1522 CKO.t4 a_6375_8213.t1 VDDD.t1521 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X95 a_2255_5185.t1 CF[8].t5 VSSD.t1639 VSSD.t1638 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X96 a_4145_5309.t0 a_3583_4917.t4 VSSD.t405 VSSD.t404 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X97 VSSD.t1546 VDDD.t1987 VSSD.t1545 VSSD.t1228 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X98 VDDD.t1272 a_2877_10357.t4 a_2767_10383.t0 VDDD.t1271 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X99 SWN[7].t1 a_1835_5461.t3 VDDD.t70 VDDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X100 VDDD.t498 VSSD.t1859 VDDD.t497 VDDD.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X101 a_2029_8573.t1 a_1467_8181.t3 VSSD.t767 VSSD.t675 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X102 VSSD.t1544 VDDD.t1988 VSSD.t1543 VSSD.t1542 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X103 CF[1].t3 a_5055_3285.t4 VSSD.t692 VSSD.t691 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X104 a_1789_8751.t0 a_1754_9003.t4 a_1467_8725.t0 VSSD.t1587 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X105 VDDD.t1545 a_7331_9269.t6 x3/COMP_BUF_N.t7 VDDD.t1544 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X106 VSSD.t1541 VDDD.t1989 VSSD.t1540 VSSD.t1254 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X107 a_5341_5487.t1 a_4779_5461.t3 VSSD.t836 VSSD.t835 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X108 VDDD.t1228 EN.t2 a_1467_8725.t2 VDDD.t1227 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X109 a_4895_10357.t0 a_4739_10625.t3 a_5040_10383.t1 VDDD.t1229 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X110 clknet_1_0__leaf_CLK.t31 a_7654_4943.t10 VDDD.t1978 VDDD.t1977 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X111 VSSD.t235 CLKS.t22 a_10281_4221.t1 VSSD.t234 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X112 VSSD.t134 a_6813_7093.t8 clknet_0_CLK.t31 VSSD.t133 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X113 a_2840_11837.t2 x2/net9.t5 VSSD.t818 VSSD.t817 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X114 VDDD.t501 VSSD.t1860 VDDD.t500 VDDD.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X115 a_6803_2741.t2 a_7090_2899.t4 VDDD.t1303 VDDD.t1302 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X116 VSSD.t1159 CKO.t5 a_8951_8751.t1 VSSD.t1158 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X117 a_4515_12381.t2 EN.t3 VDDD.t639 VDDD.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X118 SWN[2].t3 a_4411_6005.t4 VSSD.t38 VSSD.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X119 FINAL.t15 a_5307_7093.t6 VSSD.t910 VSSD.t909 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X120 a_9832_9661.t2 SWP[0].t4 VDDD.t1483 VDDD.t1482 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X121 VDDD.t312 CLKS.t23 a_5960_3677.t0 VDDD.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X122 VDDD.t1232 a_8275_6335.t3 a_8262_6031.t0 VDDD.t1231 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 SWN[5].t1 a_3767_8181.t3 VDDD.t8 VDDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X124 a_9372_10927.t2 x2/net5.t4 VSSD.t844 VSSD.t843 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X125 SWN[6].t3 a_3859_6549.t4 VSSD.t814 VSSD.t813 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X126 a_10032_8751.t1 a_9117_8751.t2 a_9685_8993.t0 VSSD.t723 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X127 a_10032_7663.t2 a_8951_7663.t3 a_9685_7905.t1 VDDD.t1701 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X128 a_3342_6031.t0 a_2623_6273.t2 a_2779_6005.t1 VSSD.t49 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X129 a_6081_7663.t1 a_5915_7663.t2 VSSD.t727 VSSD.t726 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X130 a_8008_10927.t0 a_7093_10927.t2 a_7661_11169.t3 VSSD.t194 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X131 a_9467_8751.t1 a_9117_8751.t3 a_9372_8751.t0 VDDD.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X132 a_4625_12257.t2 a_4407_12015.t4 VDDD.t1612 VDDD.t1611 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X133 VSSD.t962 a_3399_10687.t3 x2/net6.t3 VSSD.t961 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X134 VDDD.t1728 x3/COMP_BUF_P.t16 a_5734_2767.t0 VDDD.t1727 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X135 a_4343_4917.t1 a_4187_5185.t2 a_4488_4943.t2 VDDD.t1463 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X136 a_9274_10383.t0 a_8197_10389.t2 a_9112_10761.t3 VDDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X137 clknet_1_0__leaf_CLK.t23 a_7654_4943.t11 VSSD.t1603 VSSD.t1602 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X138 a_8459_4159.t1 a_8284_4233.t4 a_8638_4221.t1 VSSD.t964 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X139 a_6855_6717.t1 CF[1].t5 VSSD.t423 VSSD.t422 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X140 clknet_0_CLK.t15 a_6813_7093.t9 VDDD.t180 VDDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X141 VDDD.t407 a_2779_6005.t4 a_2710_6031.t0 VDDD.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X142 VSSD.t1539 VDDD.t1990 VSSD.t1538 VSSD.t1537 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X143 a_10111_5487.t3 a_9595_5487.t2 a_10016_5487.t3 VSSD.t1128 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X144 a_10676_5487.t2 a_9595_5487.t3 a_10329_5729.t3 VDDD.t1467 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X145 a_10877_6575.t0 a_9687_6575.t3 a_10768_6575.t0 VSSD.t683 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X146 VSSD.t1822 a_10667_9599.t3 DOUT[0].t3 VSSD.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X147 VDDD.t1198 a_8435_8181.t7 x3/COMP_BUF_P.t7 VDDD.t1197 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X148 VDDD.t1687 a_7824_4399.t4 a_7999_4373.t1 VDDD.t1686 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X149 a_9575_9117.t0 a_8951_8751.t2 a_9467_8751.t2 VDDD.t1961 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X150 VDDD.t1518 a_10237_6005.t4 a_10127_6031.t2 VDDD.t1517 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X151 VSSD.t1178 a_7331_9269.t7 x3/COMP_BUF_N.t15 VSSD.t1177 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X152 VSSD.t822 a_6077_9813.t10 clknet_1_1__leaf_CLK.t30 VSSD.t821 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X153 VSSD.t966 a_7631_8511.t3 a_7565_8585.t1 VSSD.t965 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X154 VSSD.t1536 VDDD.t1991 VSSD.t1535 VSSD.t1437 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X155 a_7090_9003.t1 a_7368_9019.t2 a_7324_9117.t1 VDDD.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X156 a_4906_4943.t3 a_4148_5059.t2 a_4343_4917.t0 VDDD.t582 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X157 a_2856_10927.t0 a_1941_10927.t2 a_2509_11169.t3 VSSD.t666 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X158 VSSD.t1619 a_2439_4541.t2 a_2400_4667.t1 VSSD.t1618 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X159 a_7153_8573.t1 a_7109_8181.t4 a_6987_8585.t1 VSSD.t1157 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X160 a_4764_4765.t2 a_4550_4765.t4 VDDD.t1408 VDDD.t1407 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X161 a_7348_5487.t1 x3/COMP_BUF_P.t17 VSSD.t1722 VSSD.t1721 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X162 VDDD.t1527 a_7948_7637.t4 clkload0.X.t7 VDDD.t1526 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X163 a_5481_11837.t1 a_5102_11471.t4 a_5409_11837.t0 VSSD.t110 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X164 VDDD.t831 x3/COMP_BUF_N.t16 a_3342_6031.t1 VDDD.t830 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X165 VDDD.t504 VSSD.t1861 VDDD.t503 VDDD.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X166 a_7827_3855.t1 CLKS.t24 VDDD.t314 VDDD.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X167 a_7093_3311.t1 a_6927_3311.t2 VSSD.t328 VSSD.t327 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X168 a_10207_3311.t0 a_9761_3311.t3 a_10111_3311.t0 VSSD.t856 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X169 a_6813_7093.t2 CLK.t1 VDDD.t1495 VDDD.t1494 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X170 a_4765_8573.t0 CLKS.t25 VSSD.t251 VSSD.t250 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X171 a_4411_2741.t2 a_4698_2899.t4 VDDD.t230 VDDD.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X172 VSSD.t826 a_3859_4373.t3 SWP[6].t3 VSSD.t825 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X173 VSSD.t253 CLKS.t26 a_4181_8751.t0 VSSD.t252 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X174 a_10584_6409.t1 a_9669_6037.t2 a_10237_6005.t0 VSSD.t394 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X175 VDDD.t1307 a_7631_8511.t4 DOUT[5].t1 VDDD.t1306 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X176 a_6251_10901.t2 EN.t4 VDDD.t641 VDDD.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X177 a_7164_4399.t0 x3/COMP_BUF_P.t18 VDDD.t1730 VDDD.t1729 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X178 VDDD.t709 a_2439_5629.t2 a_2400_5755.t0 VDDD.t708 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X179 a_5659_3453.t1 clknet_1_0__leaf_CLK.t33 VSSD.t55 VSSD.t54 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 a_9729_7663.t0 a_9685_7905.t4 a_9563_7663.t1 VSSD.t645 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X181 VSSD.t688 x2/net13.t8 CLKS.t5 VSSD.t687 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X182 VDDD.t643 EN.t5 a_1467_8181.t2 VDDD.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X183 a_4550_6941.t3 a_4463_6717.t2 a_4146_6827.t2 VDDD.t1682 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X184 a_10233_7497.t1 a_9043_7125.t2 a_10124_7497.t2 VSSD.t1720 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X185 a_4365_7663.t1 a_4330_7915.t4 a_4043_7637.t2 VSSD.t1759 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X186 VSSD.t997 a_10667_5247.t4 a_10601_5321.t1 VSSD.t996 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X187 VDDD.t507 VSSD.t1862 VDDD.t506 VDDD.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X188 VSSD.t1534 VDDD.t1992 VSSD.t1533 VSSD.t1532 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X189 a_2019_6005.t2 a_2306_6163.t4 VDDD.t879 VDDD.t878 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X190 VSSD.t255 CLKS.t27 a_2341_6397.t0 VSSD.t254 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X191 a_11030_3311.t0 CLKS.t28 VSSD.t257 VSSD.t256 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X192 DOUT[5].t3 a_7631_8511.t5 VSSD.t968 VSSD.t967 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X193 VSSD.t259 CLKS.t29 a_7521_4399.t1 VSSD.t258 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X194 VDDD.t1384 a_6251_6549.t3 SWN[1].t1 VDDD.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X195 a_7999_4373.t0 a_7824_4399.t5 a_8178_4399.t0 VSSD.t1693 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X196 VDDD.t857 a_5055_3285.t5 CF[1].t1 VDDD.t856 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X197 a_10189_5309.t1 a_10145_4917.t4 a_10023_5321.t0 VSSD.t861 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X198 a_2595_5724.t2 a_2400_5755.t2 a_2905_5487.t0 VSSD.t743 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X199 VDDD.t510 VSSD.t1863 VDDD.t509 VDDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X200 a_8100_6409.t3 a_7185_6037.t2 a_7753_6005.t1 VSSD.t708 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X201 VDDD.t316 CLKS.t30 a_7156_6941.t1 VDDD.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X202 VDDD.t170 a_5147_11989.t3 x2/TRIG1.t1 VDDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X203 clknet_1_1__leaf_CLK.t29 a_6077_9813.t11 VSSD.t824 VSSD.t823 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X204 a_10746_3855.t1 a_9669_3861.t2 a_10584_4233.t3 VDDD.t1928 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X205 a_10329_5729.t2 a_10111_5487.t4 VDDD.t1210 VDDD.t1209 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X206 a_7873_8751.t1 a_7494_9117.t4 a_7801_8751.t1 VSSD.t87 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X207 VDDD.t409 a_1835_4373.t4 SWP[7].t1 VDDD.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X208 a_7365_8751.t0 a_6803_8725.t3 VSSD.t290 VSSD.t289 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X209 CKO.t0 a_8615_7457.t3 VDDD.t242 VDDD.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X210 a_7551_5853.t0 CLKS.t31 VDDD.t392 VDDD.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X211 a_7624_4221.t0 x3/COMP_BUF_P.t19 VDDD.t1732 VDDD.t1731 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X212 x3/COMP_BUF_P.t14 a_8435_8181.t8 VSSD.t848 VSSD.t847 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X213 a_2122_5739.t0 a_2439_5629.t3 a_2397_5487.t1 VSSD.t540 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X214 a_7185_6037.t1 a_7019_6037.t2 VSSD.t842 VSSD.t841 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X215 a_9372_7663.t3 SWP[4].t4 VSSD.t840 VSSD.t839 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X216 VSSD.t668 x3/COMP_BUF_N.t17 a_5182_6941.t2 VSSD.t667 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X217 clknet_1_1__leaf_CLK.t14 a_6077_9813.t12 VDDD.t1181 VDDD.t1180 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X218 VDDD.t1950 x3/COMP_BUF_N.t18 a_5182_6941.t1 VDDD.t1949 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X219 a_3031_11849.t1 a_2585_11477.t2 a_2935_11849.t2 VSSD.t0 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X220 VDDD.t373 a_1467_8725.t3 DOUT[8].t1 VDDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X221 clknet_1_0__leaf_CLK.t24 a_7654_4943.t12 VDDD.t1608 VDDD.t1607 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X222 a_8701_7457.t1 FINAL.t16 a_8615_7457.t1 VSSD.t457 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X223 a_5729_11169.t3 a_5511_10927.t4 VSSD.t11 VSSD.t10 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X224 VDDD.t513 VSSD.t1864 VDDD.t512 VDDD.t511 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X225 a_4775_4233.t0 a_4259_3861.t3 a_4680_4221.t2 VSSD.t665 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X226 VDDD.t375 a_10759_4159.t3 CF[5].t1 VDDD.t374 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X227 VDDD.t516 VSSD.t1865 VDDD.t515 VDDD.t514 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X228 a_4380_4765.t0 a_3859_4373.t4 VDDD.t1183 VDDD.t1182 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X229 VSSD.t1531 VDDD.t1993 VSSD.t1530 VSSD.t1510 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X230 a_5377_3311.t1 a_5342_3563.t4 a_5055_3285.t0 VSSD.t155 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X231 a_2935_11849.t0 a_2419_11477.t2 a_2840_11837.t3 VSSD.t671 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X232 x2/net4.t1 a_8183_10901.t3 VDDD.t962 VDDD.t961 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X233 VSSD.t737 a_9287_10687.t3 x2/net5.t3 VSSD.t736 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X234 a_9577_9839.t0 a_9411_9839.t2 VDDD.t1925 VDDD.t1924 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X235 VSSD.t479 EN.t6 a_1789_8751.t1 VSSD.t478 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X236 VDDD.t519 VSSD.t1866 VDDD.t518 VDDD.t517 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X237 clknet_1_1__leaf_CLK.t28 a_6077_9813.t13 VSSD.t653 VSSD.t652 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X238 VDDD.t1378 a_7011_6812.t4 a_6942_6941.t0 VDDD.t1377 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X239 a_2767_10383.t1 a_2143_10389.t3 a_2659_10761.t1 VDDD.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X240 VDDD.t522 VSSD.t1867 VDDD.t521 VDDD.t520 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X241 a_8126_2767.t3 a_7407_3009.t3 a_7563_2741.t2 VSSD.t412 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X242 a_8183_5461.t0 CLKS.t32 VDDD.t394 VDDD.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X243 a_3859_6549.t2 a_4146_6827.t4 VDDD.t1642 VDDD.t1641 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X244 a_2399_11293.t0 a_1775_10927.t3 a_2291_10927.t1 VDDD.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X245 x2/net6.t2 a_3399_10687.t4 VSSD.t205 VSSD.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X246 a_10759_3071.t2 CLKS.t33 VDDD.t396 VDDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X247 VSSD.t1529 VDDD.t1994 VSSD.t1528 VSSD.t1527 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X248 a_2071_8893.t1 CKO.t6 VSSD.t1161 VSSD.t1160 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X249 VSSD.t1125 a_4187_5185.t3 a_4148_5059.t1 VSSD.t1124 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X250 VDDD.t846 a_4895_10357.t4 a_4826_10383.t2 VDDD.t845 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X251 clknet_1_0__leaf_CLK.t25 a_7654_4943.t13 VSSD.t1605 VSSD.t1604 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X252 a_9761_5487.t1 a_9595_5487.t4 VSSD.t1802 VSSD.t1801 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X253 a_4972_12015.t2 a_3891_12015.t2 a_4625_12257.t1 VDDD.t1346 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X254 a_6251_10901.t0 a_6076_10927.t4 a_6430_10927.t0 VSSD.t682 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X255 VSSD.t928 a_5383_5629.t2 a_5344_5755.t1 VSSD.t927 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X256 CF[7].t3 a_10851_5461.t3 VSSD.t686 VSSD.t685 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X257 VDDD.t1104 a_3859_6549.t5 SWN[6].t1 VDDD.t1103 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X258 VDDD.t525 VSSD.t1868 VDDD.t524 VDDD.t523 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X259 a_2856_10927.t2 a_1775_10927.t4 a_2509_11169.t2 VDDD.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X260 VDDD.t398 CLKS.t34 a_4764_6941.t0 VDDD.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X261 a_4458_8207.t3 a_4332_8323.t2 a_4054_8339.t2 VSSD.t1734 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X262 VDDD.t1803 VSSD.t1869 VDDD.t1802 VDDD.t1015 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X263 VDDD.t1938 a_7661_11169.t4 a_7551_11293.t0 VDDD.t1937 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X264 a_2595_7900.t1 a_2439_7805.t2 a_2740_8029.t1 VDDD.t1402 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X265 VDDD.t1806 VSSD.t1870 VDDD.t1805 VDDD.t1804 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X266 a_2905_9839.t1 a_2526_10205.t4 a_2833_9839.t1 VSSD.t581 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X267 VSSD.t348 a_7171_7637.t3 a_7105_7663.t1 VSSD.t347 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X268 VDDD.t1547 a_7331_9269.t8 x3/COMP_BUF_N.t6 VDDD.t1546 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X269 a_2397_9839.t0 a_1835_9813.t3 VSSD.t309 VSSD.t308 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X270 VDDD.t1809 VSSD.t1871 VDDD.t1808 VDDD.t1807 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X271 VSSD.t316 CLKS.t35 a_1973_5309.t0 VSSD.t315 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X272 VSSD.t1163 CKO.t7 a_5915_7663.t1 VSSD.t1162 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X273 DOUT[0].t1 a_10667_9599.t4 VDDD.t1948 VDDD.t1947 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X274 a_4733_3133.t1 a_4698_2899.t5 a_4411_2741.t1 VSSD.t182 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X275 DOUT[6].t1 a_7171_7637.t4 VDDD.t1557 VDDD.t1556 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X276 VSSD.t1526 VDDD.t1995 VSSD.t1525 VSSD.t1411 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X277 a_4330_7915.t2 a_4608_7931.t2 a_4564_8029.t1 VDDD.t1603 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X278 VDDD.t1610 a_7654_4943.t14 clknet_1_0__leaf_CLK.t26 VDDD.t1609 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X279 FINAL.t14 a_5307_7093.t7 VSSD.t912 VSSD.t911 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X280 VDDD.t1907 a_4463_8893.t2 a_4424_9019.t0 VDDD.t1906 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X281 VDDD.t1811 VSSD.t1872 VDDD.t1810 VDDD.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X282 VSSD.t1761 a_3675_11775.t3 x2/net10.t3 VSSD.t1760 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X283 VDDD.t1814 VSSD.t1873 VDDD.t1813 VDDD.t1812 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X284 VSSD.t1524 VDDD.t1996 VSSD.t1523 VSSD.t1522 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X285 a_2537_8573.t0 a_2158_8207.t4 a_2465_8573.t0 VSSD.t227 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X286 a_10667_5247.t0 CLKS.t36 VDDD.t400 VDDD.t399 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X287 VDDD.t1414 a_10299_7423.t3 DOUT[3].t1 VDDD.t1413 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X288 VSSD.t318 CLKS.t37 a_8425_6603.t0 VSSD.t317 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X289 VDDD.t402 CLKS.t38 a_3859_4373.t2 VDDD.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X290 a_3158_8029.t1 a_2400_7931.t2 a_2595_7900.t0 VDDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X291 VDDD.t752 a_4411_2741.t3 SWP[4].t1 VDDD.t751 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X292 a_7563_2741.t3 a_7407_3009.t4 a_7708_2767.t2 VDDD.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X293 a_10194_8029.t1 a_9117_7663.t2 a_10032_7663.t1 VDDD.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X294 VDDD.t441 a_4647_7805.t2 a_4608_7931.t0 VDDD.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X295 a_4619_8988.t0 a_4424_9019.t2 a_4929_8751.t0 VSSD.t1576 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X296 a_7109_8181.t1 a_6891_8585.t4 VSSD.t400 VSSD.t399 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X297 a_5734_2767.t2 a_5015_3009.t2 a_5171_2741.t0 VSSD.t740 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X298 VSSD.t1669 CLKS.t39 a_10373_5487.t1 VSSD.t1668 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X299 VSSD.t1521 VDDD.t1997 VSSD.t1520 VSSD.t1519 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X300 VSSD.t1518 VDDD.t1998 VSSD.t1517 VSSD.t1516 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X301 a_10851_3285.t1 a_10676_3311.t4 a_11030_3311.t1 VSSD.t725 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X302 a_7443_5487.t3 a_6927_5487.t2 a_7348_5487.t3 VSSD.t551 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X303 CLKS.t6 x2/net13.t9 VSSD.t690 VSSD.t689 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X304 VDDD.t1816 VSSD.t1874 VDDD.t1815 VDDD.t1790 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X305 CLKS.t7 x2/net13.t10 VDDD.t1352 VDDD.t1351 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X306 VSSD.t1515 VDDD.t1999 VSSD.t1514 VSSD.t1513 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X307 VDDD.t1927 a_8183_5461.t3 a_8170_5853.t1 VDDD.t1926 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X308 a_10115_6409.t0 a_9669_6037.t3 a_10019_6409.t1 VSSD.t395 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X309 DOUT[3].t3 a_10299_7423.t4 VSSD.t1078 VSSD.t1077 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X310 SWN[0].t1 a_3859_8725.t3 VDDD.t948 VDDD.t947 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X311 a_4775_4233.t2 a_4425_3861.t2 a_4680_4221.t3 VDDD.t1943 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X312 VDDD.t182 a_6813_7093.t10 clknet_0_CLK.t14 VDDD.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X313 DOUT[9].t3 a_1835_7637.t3 VSSD.t124 VSSD.t123 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X314 VSSD.t1512 VDDD.t2000 VSSD.t1511 VSSD.t1510 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X315 a_2291_10927.t0 a_1775_10927.t5 a_2196_10927.t2 VSSD.t527 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X316 a_8452_10749.t1 x2/net4.t4 VDDD.t692 VDDD.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X317 a_10127_3855.t1 a_9503_3861.t2 a_10019_4233.t1 VDDD.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X318 a_4181_4399.t0 a_4146_4651.t4 a_3859_4373.t0 VSSD.t986 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X319 VSSD.t1509 VDDD.t2001 VSSD.t1508 VSSD.t1405 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X320 a_4146_9003.t3 a_4463_8893.t3 a_4421_8751.t1 VSSD.t1794 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X321 VSSD.t369 a_8183_3285.t3 a_8117_3311.t1 VSSD.t368 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X322 VDDD.t865 a_5539_5724.t4 a_5470_5853.t2 VDDD.t864 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X323 a_7348_3311.t2 CF[1].t6 VDDD.t572 VDDD.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X324 VSSD.t1671 CLKS.t40 a_6573_6575.t0 VSSD.t1670 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X325 a_7661_3553.t0 a_7443_3311.t4 VDDD.t162 VDDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X326 VSSD.t57 clknet_1_0__leaf_CLK.t34 a_6927_3311.t1 VSSD.t56 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X327 SWP[0].t3 a_8275_6335.t4 VSSD.t884 VSSD.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X328 VSSD.t1673 CLKS.t41 a_7981_4221.t0 VSSD.t1672 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X329 clknet_1_1__leaf_CLK.t13 a_6077_9813.t14 VDDD.t820 VDDD.t819 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X330 a_7539_3311.t1 a_7093_3311.t2 a_7443_3311.t2 VSSD.t577 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X331 VSSD.t59 clknet_1_0__leaf_CLK.t35 a_9503_2773.t1 VSSD.t58 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X332 VSSD.t1675 CLKS.t42 a_7125_3133.t0 VSSD.t1674 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X333 VDDD.t102 a_2019_6005.t3 SWN[8].t1 VDDD.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X334 a_5171_6005.t3 a_5015_6273.t2 a_5316_6031.t2 VDDD.t1425 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X335 a_7494_9117.t0 a_7407_8893.t2 a_7090_9003.t0 VDDD.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X336 a_10667_5247.t1 a_10492_5321.t4 a_10846_5309.t1 VSSD.t378 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X337 a_5307_7093.t5 CF[0].t5 VSSD.t1586 VSSD.t1585 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X338 a_2740_5853.t2 a_2526_5853.t4 VDDD.t1427 VDDD.t1426 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X339 VDDD.t166 a_3675_11775.t4 a_3662_11471.t0 VDDD.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X340 a_8452_10749.t2 x2/net4.t5 VSSD.t531 VSSD.t530 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X341 VSSD.t82 a_10759_6335.t3 a_10693_6409.t1 VSSD.t81 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X342 VSSD.t768 a_1467_8181.t4 DOUT[7].t3 VSSD.t340 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X343 a_9575_9117.t1 EN.t7 VDDD.t645 VDDD.t644 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X344 a_4883_3855.t0 a_4259_3861.t4 a_4775_4233.t1 VDDD.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X345 VSSD.t136 a_6813_7093.t11 clknet_0_CLK.t30 VSSD.t135 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X346 a_5326_12015.t0 EN.t8 VSSD.t481 VSSD.t480 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X347 a_4089_8573.t1 a_4054_8339.t4 a_3767_8181.t1 VSSD.t1062 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X348 VDDD.t1620 a_10207_8725.t3 DOUT[2].t1 VDDD.t1619 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X349 VDDD.t1819 VSSD.t1875 VDDD.t1818 VDDD.t1817 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X350 SWN[8].t3 a_2019_6005.t4 VSSD.t76 VSSD.t75 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X351 VSSD.t1507 VDDD.t2002 VSSD.t1506 VSSD.t1505 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X352 a_5340_4233.t2 a_4425_3861.t3 a_4993_3829.t3 VSSD.t477 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X353 a_2309_10389.t1 a_2143_10389.t4 VSSD.t808 VSSD.t807 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X354 a_8008_3311.t0 a_6927_3311.t3 a_7661_3553.t2 VDDD.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X355 VDDD.t758 a_10851_3285.t3 a_10838_3677.t1 VDDD.t757 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X356 clknet_0_CLK.t13 a_6813_7093.t12 VDDD.t184 VDDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X357 VSSD.t181 a_7407_8893.t3 a_7368_9019.t0 VSSD.t180 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X358 a_2227_8988.t0 a_2032_9019.t2 a_2537_8751.t0 VSSD.t550 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X359 VSSD.t126 a_5147_11989.t4 a_5081_12015.t1 VSSD.t125 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X360 VDDD.t64 CF[3].t5 a_7203_3861.t0 VDDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X361 VDDD.t1345 a_10667_5247.t5 a_10654_4943.t0 VDDD.t1344 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X362 VSSD.t483 EN.t9 a_4669_12015.t1 VSSD.t482 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X363 a_5734_6031.t2 a_4976_6147.t2 a_5171_6005.t0 VDDD.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X364 VDDD.t1694 x2/TRIG1.t4 a_5734_11471.t2 VDDD.t1693 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X365 a_4343_4917.t3 a_4148_5059.t3 a_4653_5309.t1 VSSD.t941 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X366 VSSD.t886 a_8275_6335.t5 a_8209_6409.t0 VSSD.t885 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X367 VDDD.t1200 a_8435_8181.t9 x3/COMP_BUF_P.t6 VDDD.t1199 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X368 a_5090_8207.t0 a_4371_8449.t3 a_4527_8181.t1 VSSD.t1818 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X369 VDDD.t1821 VSSD.t1876 VDDD.t1820 VDDD.t1750 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X370 clknet_1_0__leaf_CLK.t27 a_7654_4943.t15 VSSD.t1607 VSSD.t1606 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X371 VDDD.t1952 x3/COMP_BUF_N.t19 a_8126_9117.t1 VDDD.t1951 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X372 VDDD.t384 a_10237_2741.t4 a_10127_2767.t1 VDDD.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X373 a_7535_6409.t2 a_7185_6037.t3 a_7440_6397.t3 VDDD.t868 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X374 SWP[5].t3 a_5515_4159.t5 VSSD.t1821 VSSD.t1820 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X375 a_5383_5629.t0 CF[9].t4 VDDD.t1222 VDDD.t1221 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X376 VSSD.t655 a_6077_9813.t15 clknet_1_1__leaf_CLK.t27 VSSD.t654 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X377 a_5409_6397.t0 CLKS.t43 VSSD.t1677 VSSD.t1676 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X378 a_8183_10901.t0 a_8008_10927.t5 a_8362_10927.t0 VSSD.t475 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X379 a_7011_6812.t3 a_6855_6717.t2 a_7156_6941.t2 VDDD.t611 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X380 VDDD.t1529 a_7948_7637.t5 clkload0.X.t6 VDDD.t1528 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X381 a_7331_9269.t4 COMP_N.t1 VSSD.t566 VSSD.t565 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X382 a_7551_11293.t1 EN.t10 VDDD.t1586 VDDD.t1585 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X383 VDDD.t1930 a_10851_5461.t4 CF[7].t1 VDDD.t1929 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X384 a_3158_8029.t0 a_2439_7805.t3 a_2595_7900.t2 VSSD.t1063 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X385 VDDD.t1824 VSSD.t1877 VDDD.t1823 VDDD.t1822 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X386 a_4425_3861.t1 a_4259_3861.t5 VSSD.t397 VSSD.t396 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X387 VSSD.t1679 CLKS.t44 a_4733_3133.t0 VSSD.t1678 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X388 a_6891_8585.t0 a_6375_8213.t3 a_6796_8573.t0 VSSD.t699 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X389 a_9685_7905.t2 a_9467_7663.t4 VDDD.t1902 VDDD.t1901 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X390 a_5458_10383.t2 a_4739_10625.t4 a_4895_10357.t1 VSSD.t720 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X391 VDDD.t76 x2/net11.t4 x2/TRIG2.t0 VDDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X392 a_9685_11169.t2 a_9467_10927.t4 VSSD.t1792 VSSD.t1791 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X393 a_2439_7805.t0 CKO.t8 VDDD.t1524 VDDD.t1523 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X394 a_7657_11849.t1 a_6467_11477.t2 a_7548_11849.t0 VSSD.t960 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X395 a_7551_11293.t2 a_6927_10927.t2 a_7443_10927.t1 VDDD.t1905 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X396 a_7643_6031.t2 a_7019_6037.t3 a_7535_6409.t1 VDDD.t1194 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X397 x2/TRIG1.t3 a_5147_11989.t5 VSSD.t128 VSSD.t127 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X398 a_5015_3009.t1 CF[4].t5 VSSD.t626 VSSD.t625 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X399 a_10111_5487.t1 a_9761_5487.t2 a_10016_5487.t0 VDDD.t701 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X400 clknet_0_CLK.t29 a_6813_7093.t13 VSSD.t138 VSSD.t137 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X401 a_10023_9839.t1 a_9577_9839.t2 a_9927_9839.t3 VSSD.t532 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X402 a_9924_4221.t1 CF[6].t4 VDDD.t1630 VDDD.t1629 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X403 CF[2].t0 a_6803_2741.t3 VDDD.t1277 VDDD.t1276 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X404 VSSD.t1706 SWP[9].t4 a_3158_8029.t2 VSSD.t1705 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X405 VSSD.t1504 VDDD.t2003 VSSD.t1503 VSSD.t1502 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X406 a_9467_8751.t3 a_8951_8751.t3 a_9372_8751.t1 VSSD.t1833 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X407 a_6803_8725.t1 a_7090_9003.t5 VDDD.t439 VDDD.t438 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X408 a_7574_6941.t2 a_6816_6843.t2 a_7011_6812.t0 VDDD.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X409 a_7171_7637.t0 a_6996_7663.t4 a_7350_7663.t0 VSSD.t197 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X410 a_6185_10927.t1 a_4995_10927.t2 a_6076_10927.t2 VSSD.t664 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X411 a_6077_9813.t0 clknet_0_CLK.t33 VDDD.t22 VDDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X412 VDDD.t1588 EN.t11 a_1835_9813.t2 VDDD.t1587 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X413 clknet_1_1__leaf_CLK.t26 a_6077_9813.t16 VSSD.t657 VSSD.t656 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X414 VSSD.t1609 a_7654_4943.t16 clknet_1_0__leaf_CLK.t28 VSSD.t1608 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X415 VDDD.t1614 x2/net6.t4 x2/net12.t1 VDDD.t1613 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X416 a_8446_3855.t1 a_7369_3861.t2 a_8284_4233.t2 VDDD.t895 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X417 VDDD.t232 a_10145_4917.t5 a_10035_4943.t2 VDDD.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X418 VDDD.t1341 a_5515_4159.t6 SWP[5].t1 VDDD.t1340 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X419 a_2399_11293.t2 EN.t12 VDDD.t1590 VDDD.t1589 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X420 VSSD.t521 a_2439_9981.t2 a_2400_10107.t0 VSSD.t520 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X421 VSSD.t9 a_10667_9813.t4 DOUT[1].t3 VSSD.t8 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X422 VDDD.t1250 a_5307_7093.t8 FINAL.t7 VDDD.t1249 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X423 VSSD.t357 a_10851_3285.t4 CF[4].t2 VSSD.t356 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X424 VDDD.t1541 a_10768_6575.t4 a_10943_6549.t1 VDDD.t1540 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X425 a_9575_11293.t1 EN.t13 VDDD.t1592 VDDD.t1591 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X426 VDDD.t1424 a_7477_4641.t4 a_7367_4765.t0 VDDD.t1423 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X427 VDDD.t1826 VSSD.t1878 VDDD.t1825 VDDD.t1755 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X428 a_3017_6397.t1 CLKS.t45 VSSD.t1681 VSSD.t1680 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X429 a_7705_10927.t0 a_7661_11169.t5 a_7539_10927.t0 VSSD.t1813 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X430 a_4929_4399.t1 a_4550_4765.t5 a_4857_4399.t1 VSSD.t1068 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X431 VSSD.t1501 VDDD.t2004 VSSD.t1500 VSSD.t1499 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X432 VSSD.t1498 VDDD.t2005 VSSD.t1497 VSSD.t1496 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X433 SWP[4].t3 a_4411_2741.t4 VSSD.t587 VSSD.t586 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X434 a_7011_6812.t1 a_6816_6843.t3 a_7321_6575.t1 VSSD.t101 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X435 VSSD.t1100 COMP_P.t0 a_8435_8181.t2 VSSD.t1099 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X436 VSSD.t345 a_2071_8449.t2 a_2032_8323.t0 VSSD.t344 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X437 CF[9].t3 a_10943_6549.t4 VSSD.t792 VSSD.t791 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X438 a_10219_3677.t0 CLKS.t46 VDDD.t1673 VDDD.t1672 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X439 a_9209_7125.t0 a_9043_7125.t3 VDDD.t1723 VDDD.t1722 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X440 a_7948_7637.t1 clknet_1_0__leaf_CLK.t36 VDDD.t360 VDDD.t359 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X441 a_4312_12015.t2 x2/net10.t4 VDDD.t1878 VDDD.t1877 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X442 x2/net7.t1 a_4135_10357.t3 VDDD.t116 VDDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X443 a_9577_4949.t1 a_9411_4949.t3 VSSD.t1115 VSSD.t1114 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X444 a_4734_8029.t1 a_4647_7805.t3 a_4330_7915.t0 VDDD.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X445 VDDD.t120 a_10492_9839.t4 a_10667_9813.t0 VDDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X446 VDDD.t1594 EN.t14 a_2740_8029.t2 VDDD.t1593 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X447 a_1938_5075.t3 a_2216_5059.t2 a_2172_4943.t1 VDDD.t1373 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X448 a_2924_6031.t0 a_2710_6031.t4 VDDD.t1543 VDDD.t1542 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X449 VSSD.t1495 VDDD.t2006 VSSD.t1494 VSSD.t1493 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X450 a_10237_3829.t2 a_10019_4233.t4 VSSD.t447 VSSD.t446 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X451 VDDD.t745 a_2595_10076.t4 a_2526_10205.t1 VDDD.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X452 a_4330_7915.t3 a_4647_7805.t4 a_4605_7663.t1 VSSD.t1742 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X453 VDDD.t249 a_3399_10687.t5 a_3386_10383.t1 VDDD.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X454 a_10019_6409.t3 a_9503_6037.t2 a_9924_6397.t3 VSSD.t776 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X455 a_7407_8893.t0 CF[3].t6 VDDD.t66 VDDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X456 a_9577_9301.t0 a_9411_9301.t2 VDDD.t186 VDDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X457 a_6538_6827.t0 a_6855_6717.t3 a_6813_6575.t1 VSSD.t450 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X458 a_8183_3285.t1 a_8008_3311.t4 a_8362_3311.t0 VSSD.t516 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X459 VDDD.t792 a_3031_10901.t5 a_3018_11293.t0 VDDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X460 VSSD.t750 a_2227_8181.t4 a_2158_8207.t3 VSSD.t293 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X461 VDDD.t1268 a_2595_7900.t4 a_2526_8029.t1 VDDD.t1267 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X462 VSSD.t774 a_3859_8725.t4 SWN[0].t3 VSSD.t773 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X463 VDDD.t386 a_7456_8585.t4 a_7631_8511.t0 VDDD.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X464 VDDD.t1364 a_7937_3829.t4 a_7827_3855.t2 VDDD.t1363 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X465 VDDD.t1366 a_10032_10927.t4 a_10207_10901.t0 VDDD.t1365 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X466 a_2553_10927.t0 a_2509_11169.t4 a_2387_10927.t1 VSSD.t275 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X467 a_7548_11849.t2 a_6633_11477.t2 a_7201_11445.t2 VSSD.t1737 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X468 VSSD.t261 CLKS.t47 a_4089_8573.t0 VSSD.t260 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X469 a_2227_8181.t1 a_2032_8323.t3 a_2537_8573.t1 VSSD.t550 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X470 VDDD.t1829 VSSD.t1879 VDDD.t1828 VDDD.t1827 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X471 VSSD.t1492 VDDD.t2007 VSSD.t1491 VSSD.t1490 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X472 a_10851_3285.t0 CLKS.t48 VDDD.t318 VDDD.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X473 VDDD.t1832 VSSD.t1880 VDDD.t1831 VDDD.t1830 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X474 VDDD.t320 CLKS.t49 a_3583_4917.t0 VDDD.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 a_4288_8207.t0 a_3767_8181.t4 VDDD.t10 VDDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X476 VDDD.t1570 CF[0].t6 a_5307_7093.t2 VDDD.t1569 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X477 a_4837_8573.t0 a_4458_8207.t4 a_4765_8573.t1 VSSD.t335 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X478 VSSD.t620 a_3031_10901.t6 x2/net9.t3 VSSD.t619 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X479 a_5815_3548.t2 a_5620_3579.t2 a_6125_3311.t1 VSSD.t795 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X480 VSSD.t659 a_6077_9813.t17 clknet_1_1__leaf_CLK.t25 VSSD.t658 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X481 VDDD.t1954 x3/COMP_BUF_N.t20 a_5366_8029.t2 VDDD.t1953 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X482 VDDD.t1835 VSSD.t1881 VDDD.t1834 VDDD.t1833 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X483 VDDD.t474 COMP_N.t2 a_7331_9269.t2 VDDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X484 x2/net3.t2 a_7723_11775.t3 VSSD.t1815 VSSD.t1814 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X485 a_6076_10927.t1 a_5161_10927.t2 a_5729_11169.t0 VSSD.t65 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X486 a_6796_8573.t2 SWP[5].t4 VDDD.t818 VDDD.t817 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X487 VDDD.t1531 a_7948_7637.t6 clkload0.X.t5 VDDD.t1530 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X488 a_9372_7663.t2 SWP[4].t5 VDDD.t1193 VDDD.t1192 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X489 VDDD.t1838 VSSD.t1882 VDDD.t1837 VDDD.t1836 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X490 a_5342_3563.t0 a_5659_3453.t2 a_5617_3311.t0 VSSD.t631 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X491 a_2306_6163.t2 a_2584_6147.t3 a_2540_6031.t1 VDDD.t949 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X492 VSSD.t1599 a_10667_5247.t6 CF[6].t3 VSSD.t1598 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X493 a_10016_5487.t1 CF[8].t6 VDDD.t1643 VDDD.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X494 VDDD.t1840 VSSD.t1883 VDDD.t1839 VDDD.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X495 a_8275_6335.t1 a_8100_6409.t4 a_8454_6397.t1 VSSD.t1810 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X496 a_6539_8029.t0 a_5915_7663.t3 a_6431_7663.t1 VDDD.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X497 a_10145_10081.t3 a_9927_9839.t4 VSSD.t1812 VSSD.t853 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X498 a_4135_10357.t0 a_4422_10515.t4 VDDD.t620 VDDD.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X499 VDDD.t322 CLKS.t50 a_4488_4943.t0 VDDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X500 a_4274_4943.t2 a_4148_5059.t4 a_3870_5075.t3 VSSD.t942 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X501 clknet_0_CLK.t28 a_6813_7093.t14 VSSD.t187 VSSD.t186 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X502 a_1651_4917.t1 a_1938_5075.t4 VDDD.t1873 VDDD.t1872 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X503 VDDD.t699 a_2071_8893.t2 a_2032_9019.t0 VDDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X504 CLKS.t8 x2/net13.t11 VSSD.t1011 VSSD.t1010 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X505 VDDD.t1663 a_10584_4233.t4 a_10759_4159.t2 VDDD.t1662 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X506 a_7109_8181.t0 a_6891_8585.t5 VDDD.t932 VDDD.t931 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X507 a_4973_6397.t0 a_4411_6005.t5 VSSD.t40 VSSD.t39 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X508 VSSD.t1597 EN.t15 a_7705_10927.t1 VSSD.t1596 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X509 VSSD.t633 a_5659_3453.t3 a_5620_3579.t1 VSSD.t632 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X510 a_2122_4651.t1 a_2400_4667.t2 a_2356_4765.t0 VDDD.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X511 a_10785_5487.t0 a_9595_5487.t5 a_10676_5487.t3 VSSD.t1803 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X512 a_9927_9839.t2 a_9577_9839.t3 a_9832_9839.t3 VDDD.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X513 VSSD.t1489 VDDD.t2008 VSSD.t1488 VSSD.t1462 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X514 a_10693_3145.t1 a_9503_2773.t2 a_10584_3145.t2 VSSD.t1694 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X515 a_8170_3677.t0 a_7093_3311.t3 a_8008_3311.t3 VDDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X516 a_3333_10761.t0 a_2143_10389.t5 a_3224_10761.t1 VSSD.t809 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X517 a_6077_9813.t1 clknet_0_CLK.t34 VDDD.t24 VDDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X518 VDDD.t234 a_6813_7093.t15 clknet_0_CLK.t12 VDDD.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X519 CLKSB.t0 CLKS.t51 VDDD.t324 VDDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X520 VDDD.t1956 a_8435_8181.t10 x3/COMP_BUF_P.t5 VDDD.t1955 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X521 VSSD.t5 a_3767_8181.t5 SWN[5].t3 VSSD.t4 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X522 VDDD.t1624 a_4625_12257.t4 a_4515_12381.t1 VDDD.t1623 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X523 VSSD.t1487 VDDD.t2009 VSSD.t1486 VSSD.t1485 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X524 VSSD.t143 CKO.t9 a_9043_7125.t1 VSSD.t142 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X525 a_9467_10927.t0 a_9117_10927.t2 a_9372_10927.t0 VDDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X526 VDDD.t362 clknet_1_0__leaf_CLK.t37 a_9595_5487.t0 VDDD.t361 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X527 VDDD.t608 a_6251_10901.t3 x2/net2.t1 VDDD.t607 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X528 VSSD.t281 a_7654_4943.t17 clknet_1_0__leaf_CLK.t5 VSSD.t280 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X529 VDDD.t592 a_10329_5729.t5 a_10219_5853.t0 VDDD.t591 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X530 VSSD.t1573 a_7171_7637.t5 DOUT[6].t3 VSSD.t1572 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X531 a_4698_11603.t1 a_4976_11587.t2 a_4932_11471.t0 VDDD.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X532 VSSD.t1039 a_7011_6812.t5 a_6942_6941.t1 VSSD.t1038 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X533 VDDD.t1264 a_8183_5461.t4 SWP[1].t1 VDDD.t1263 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X534 VDDD.t1842 VSSD.t1884 VDDD.t1841 VDDD.t1796 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X535 a_7456_8585.t1 a_6375_8213.t4 a_7109_8181.t2 VDDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X536 a_7710_11471.t0 a_6633_11477.t3 a_7548_11849.t3 VDDD.t1874 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X537 VSSD.t145 CKO.t10 a_9411_9301.t1 VSSD.t144 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X538 a_5171_2741.t1 a_5015_3009.t3 a_5316_2767.t2 VDDD.t734 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X539 a_2356_8029.t0 a_1835_7637.t4 VDDD.t1934 VDDD.t1933 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X540 clknet_1_1__leaf_CLK.t24 a_6077_9813.t18 VSSD.t661 VSSD.t660 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X541 VDDD.t364 clknet_1_0__leaf_CLK.t38 a_9503_3861.t0 VDDD.t363 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X542 clkload0.X.t4 a_7948_7637.t7 VDDD.t431 VDDD.t430 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X543 VSSD.t1170 a_3675_11775.t5 a_3609_11849.t1 VSSD.t1169 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X544 VSSD.t189 a_6813_7093.t16 clknet_0_CLK.t27 VSSD.t188 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X545 a_5458_10383.t3 a_4700_10499.t2 a_4895_10357.t3 VDDD.t418 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X546 a_7443_5487.t0 a_7093_5487.t2 a_7348_5487.t2 VDDD.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X547 a_4698_6163.t3 a_5015_6273.t3 a_4973_6397.t1 VSSD.t1090 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X548 VDDD.t1511 a_7201_11445.t4 a_7091_11471.t0 VDDD.t1510 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X549 VDDD.t901 a_9287_10687.t4 a_9274_10383.t1 VDDD.t900 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X550 a_10237_3829.t1 a_10019_4233.t5 VDDD.t603 VDDD.t602 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X551 x3/COMP_BUF_P.t13 a_8435_8181.t11 VSSD.t1828 VSSD.t1827 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X552 CF[5].t0 a_10759_4159.t4 VDDD.t833 VDDD.t832 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X553 VDDD.t1845 VSSD.t1885 VDDD.t1844 VDDD.t1843 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X554 a_10667_9599.t2 EN.t16 VDDD.t1596 VDDD.t1595 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X555 VSSD.t1728 EN.t17 a_9729_10927.t0 VSSD.t1727 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X556 VSSD.t1484 VDDD.t2010 VSSD.t1483 VSSD.t1482 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X557 a_10667_9813.t2 EN.t18 VDDD.t1865 VDDD.t1864 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X558 a_4187_5185.t0 CF[9].t5 VDDD.t1224 VDDD.t1223 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X559 VSSD.t184 a_10207_8725.t4 a_10141_8751.t0 VSSD.t183 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X560 a_3386_10383.t0 a_2309_10389.t2 a_3224_10761.t3 VDDD.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X561 a_10601_5321.t0 a_9411_4949.t4 a_10492_5321.t1 VSSD.t1116 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X562 VDDD.t1295 a_7661_3553.t4 a_7551_3677.t0 VDDD.t1294 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X563 a_5734_2767.t3 a_4976_2883.t2 a_5171_2741.t2 VDDD.t1484 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X564 VDDD.t1847 VSSD.t1886 VDDD.t1846 VDDD.t1050 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X565 VDDD.t1850 VSSD.t1887 VDDD.t1849 VDDD.t1848 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X566 VDDD.t1852 VSSD.t1888 VDDD.t1851 VDDD.t1787 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X567 VSSD.t1481 VDDD.t2011 VSSD.t1480 VSSD.t1479 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X568 a_7643_6031.t0 CLKS.t52 VDDD.t326 VDDD.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X569 VDDD.t1855 VSSD.t1889 VDDD.t1854 VDDD.t1853 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X570 a_10207_10901.t2 EN.t19 VDDD.t1867 VDDD.t1866 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X571 clknet_1_0__leaf_CLK.t6 a_7654_4943.t18 VSSD.t283 VSSD.t282 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X572 VSSD.t449 a_6251_10901.t4 a_6185_10927.t0 VSSD.t448 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X573 VDDD.t1858 VSSD.t1890 VDDD.t1857 VDDD.t1856 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X574 a_6076_10927.t3 a_4995_10927.t3 a_5729_11169.t1 VDDD.t823 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X575 VSSD.t146 CKO.t11 a_9411_9839.t1 VSSD.t144 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X576 a_9761_3311.t0 a_9595_3311.t2 VDDD.t1392 VDDD.t1391 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X577 VSSD.t501 a_8183_3285.t4 CF[0].t0 VSSD.t500 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X578 a_7551_5853.t1 a_6927_5487.t3 a_7443_5487.t2 VDDD.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X579 VSSD.t1708 x2/net12.t4 x2/net13.t4 VSSD.t1707 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X580 VSSD.t663 a_6077_9813.t19 clknet_1_1__leaf_CLK.t23 VSSD.t662 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X581 a_7801_3133.t1 CLKS.t53 VSSD.t263 VSSD.t262 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X582 a_10584_4233.t0 a_9503_3861.t3 a_10237_3829.t0 VDDD.t454 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X583 a_7563_8988.t1 a_7407_8893.t4 a_7708_9117.t1 VDDD.t1690 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X584 VSSD.t1478 VDDD.t2012 VSSD.t1477 VSSD.t1476 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X585 VDDD.t226 a_5015_6273.t4 a_4976_6147.t0 VDDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X586 a_5066_5739.t3 a_5344_5755.t2 a_5300_5853.t0 VDDD.t1291 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X587 a_10492_9839.t2 a_9577_9839.t4 a_10145_10081.t1 VSSD.t156 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X588 a_9924_6397.t1 CF[9].t6 VSSD.t874 VSSD.t873 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X589 VSSD.t1475 VDDD.t2013 VSSD.t1474 VSSD.t1473 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X590 x2/net9.t2 a_3031_10901.t7 VSSD.t622 VSSD.t621 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X591 a_10035_10205.t2 EN.t20 VDDD.t1869 VDDD.t1868 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X592 VSSD.t1472 VDDD.t2014 VSSD.t1471 VSSD.t1470 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X593 VDDD.t1861 VSSD.t1891 VDDD.t1860 VDDD.t1859 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X594 a_9669_6037.t1 a_9503_6037.t3 VSSD.t778 VSSD.t777 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X595 a_2779_6005.t2 a_2584_6147.t4 a_3089_6397.t1 VSSD.t790 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X596 VSSD.t850 a_4619_6812.t4 a_4550_6941.t1 VSSD.t849 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X597 VDDD.t1718 a_2255_5185.t2 a_2216_5059.t0 VDDD.t1717 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X598 a_6649_7905.t3 a_6431_7663.t4 VSSD.t61 VSSD.t60 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X599 VSSD.t833 a_4463_4541.t4 a_4424_4667.t1 VSSD.t832 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X600 VSSD.t1469 VDDD.t2015 VSSD.t1468 VSSD.t1448 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X601 a_4181_8751.t1 a_4146_9003.t4 a_3859_8725.t2 VSSD.t987 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X602 VSSD.t1467 VDDD.t2016 VSSD.t1466 VSSD.t1465 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X603 VSSD.t1464 VDDD.t2017 VSSD.t1463 VSSD.t1462 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X604 VSSD.t1461 VDDD.t2018 VSSD.t1460 VSSD.t1459 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X605 a_4932_6031.t1 a_4411_6005.t6 VDDD.t695 VDDD.t694 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X606 VDDD.t1871 EN.t21 a_1835_7637.t2 VDDD.t1870 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X607 a_9655_7497.t0 a_9209_7125.t2 a_9559_7497.t3 VSSD.t1711 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X608 a_5102_6031.t1 a_5015_6273.t5 a_4698_6163.t2 VDDD.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X609 VSSD.t1130 CF[2].t5 a_6743_4399.t1 VSSD.t1129 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X610 VSSD.t1824 x3/COMP_BUF_N.t21 a_4906_4943.t2 VSSD.t1823 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X611 a_2306_6163.t0 a_2623_6273.t3 a_2581_6397.t1 VSSD.t50 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X612 VDDD.t366 clknet_1_0__leaf_CLK.t39 a_7948_7637.t0 VDDD.t365 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X613 SWP[2].t1 a_7999_4373.t3 VDDD.t741 VDDD.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X614 VDDD.t1354 x2/net13.t12 CLKS.t9 VDDD.t1353 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X615 a_5409_11837.t1 EN.t22 VSSD.t1730 VSSD.t1729 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X616 a_2341_6397.t1 a_2306_6163.t5 a_2019_6005.t1 VSSD.t718 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X617 SWN[1].t3 a_6251_6549.t4 VSSD.t1043 VSSD.t1042 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X618 clkload0.X.t15 a_7948_7637.t8 VSSD.t351 VSSD.t350 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1134 ps=1.38 w=0.42 l=0.15
X619 a_7355_4399.t1 a_6909_4399.t2 a_7259_4399.t2 VSSD.t470 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X620 a_2905_5487.t1 a_2526_5853.t5 a_2833_5487.t1 VSSD.t1091 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X621 a_4973_11837.t0 a_4411_11445.t3 VSSD.t1798 VSSD.t1797 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X622 a_2342_4943.t3 a_2255_5185.t3 a_1938_5075.t0 VDDD.t1719 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X623 a_8178_4399.t1 CLKS.t54 VSSD.t265 VSSD.t264 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X624 a_2397_5487.t0 a_1835_5461.t4 VSSD.t42 VSSD.t41 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X625 a_5307_7093.t1 CF[0].t7 VDDD.t1572 VDDD.t1571 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X626 VDDD.t1321 a_10667_9599.t5 a_10654_9295.t0 VDDD.t1320 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X627 SWP[7].t3 a_1835_4373.t5 VSSD.t312 VSSD.t311 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X628 a_4550_6941.t0 a_4424_6843.t3 a_4146_6827.t0 VSSD.t677 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X629 VSSD.t1776 a_4371_8449.t4 a_4332_8323.t1 VSSD.t1775 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X630 VSSD.t1458 VDDD.t2019 VSSD.t1457 VSSD.t1351 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X631 clknet_1_1__leaf_CLK.t12 a_6077_9813.t20 VDDD.t822 VDDD.t821 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X632 VDDD.t1038 VSSD.t1892 VDDD.t1037 VDDD.t1036 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X633 clknet_1_1__leaf_CLK.t11 a_6077_9813.t21 VDDD.t126 VDDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X634 a_7654_4943.t3 clknet_0_CLK.t35 VDDD.t26 VDDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X635 a_2974_4943.t2 a_2255_5185.t4 a_2411_4917.t2 VSSD.t1717 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X636 VSSD.t116 a_5539_5724.t5 a_5470_5853.t3 VSSD.t115 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X637 VDDD.t1429 a_5171_6005.t4 a_5102_6031.t2 VDDD.t1428 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X638 a_10207_7637.t1 a_10032_7663.t5 a_10386_7663.t1 VSSD.t288 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X639 x2/net2.t0 a_6251_10901.t5 VDDD.t610 VDDD.t609 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X640 a_7661_3553.t1 a_7443_3311.t5 VSSD.t118 VSSD.t117 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X641 VDDD.t1040 VSSD.t1893 VDDD.t1039 VDDD.t1003 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X642 VDDD.t861 a_2623_6273.t4 a_2584_6147.t0 VDDD.t860 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X643 a_9669_2773.t0 a_9503_2773.t3 VDDD.t1689 VDDD.t1688 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X644 VDDD.t667 a_2411_4917.t5 a_2342_4943.t1 VDDD.t666 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X645 VDDD.t107 a_10759_6335.t4 a_10746_6031.t1 VDDD.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X646 VDDD.t1043 VSSD.t1894 VDDD.t1042 VDDD.t1041 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X647 VSSD.t1166 a_4527_8181.t4 a_4458_8207.t1 VSSD.t1165 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X648 a_4407_12015.t2 a_3891_12015.t3 a_4312_12015.t0 VSSD.t998 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X649 VDDD.t556 a_7407_3009.t5 a_7368_2883.t0 VDDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X650 VDDD.t46 a_8183_10901.t4 x2/net4.t0 VDDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X651 VDDD.t1734 x3/COMP_BUF_P.t20 a_2974_4943.t0 VDDD.t1733 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X652 a_6772_6941.t0 a_6251_6549.t5 VDDD.t1386 VDDD.t1385 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X653 VDDD.t1416 a_10299_7423.t5 a_10286_7119.t0 VDDD.t1415 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X654 clkload0.X.t3 a_7948_7637.t9 VDDD.t433 VDDD.t432 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X655 DOUT[2].t3 a_10207_8725.t5 VSSD.t1770 VSSD.t1769 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X656 a_2465_8751.t1 EN.t23 VSSD.t1731 VSSD.t514 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X657 a_2439_9981.t0 clknet_1_1__leaf_CLK.t34 VDDD.t138 VDDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X658 VSSD.t1826 x3/COMP_BUF_N.t22 a_5734_6031.t1 VSSD.t1825 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X659 a_4527_8181.t3 a_4332_8323.t3 a_4837_8573.t1 VSSD.t1735 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X660 VSSD.t1456 VDDD.t2020 VSSD.t1455 VSSD.t1454 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X661 VSSD.t1180 a_7331_9269.t9 x3/COMP_BUF_N.t14 VSSD.t1179 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X662 a_7937_3829.t2 a_7719_4233.t4 VSSD.t1724 VSSD.t1723 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X663 VDDD.t332 CLKS.t55 a_7708_2767.t1 VDDD.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X664 a_5470_5853.t1 a_5344_5755.t3 a_5066_5739.t2 VSSD.t951 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X665 a_2710_6031.t2 a_2623_6273.t5 a_2306_6163.t1 VDDD.t862 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X666 a_2526_4765.t3 a_2439_4541.t3 a_2122_4651.t2 VDDD.t1625 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X667 a_7494_2767.t1 a_7368_2883.t2 a_7090_2899.t1 VSSD.t984 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X668 a_7093_5487.t0 a_6927_5487.t4 VDDD.t159 VDDD.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X669 VDDD.t1208 a_10032_8751.t4 a_10207_8725.t2 VDDD.t1207 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X670 a_5515_4159.t0 a_5340_4233.t4 a_5694_4221.t1 VSSD.t80 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X671 CLKS.t10 x2/net13.t13 VSSD.t1013 VSSD.t1012 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X672 a_10421_6817.t3 a_10203_6575.t4 VSSD.t1701 VSSD.t1700 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X673 VDDD.t368 clknet_1_0__leaf_CLK.t40 a_9687_6575.t0 VDDD.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X674 VSSD.t191 a_6813_7093.t17 clknet_0_CLK.t26 VSSD.t190 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X675 VSSD.t1453 VDDD.t2021 VSSD.t1452 VSSD.t1451 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X676 CF[4].t3 a_10851_3285.t5 VDDD.t1412 VDDD.t1411 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X677 a_6539_8029.t2 EN.t24 VDDD.t669 VDDD.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X678 VSSD.t1450 VDDD.t2022 VSSD.t1449 VSSD.t1448 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X679 a_5960_3677.t2 a_5746_3677.t4 VDDD.t1339 VDDD.t1338 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X680 VSSD.t1447 VDDD.t2023 VSSD.t1446 VSSD.t1422 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X681 VDDD.t334 CLKS.t56 a_5316_6031.t0 VDDD.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X682 a_7705_5487.t1 a_7661_5729.t4 a_7539_5487.t1 VSSD.t618 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X683 VSSD.t84 a_10759_6335.t5 CF[8].t0 VSSD.t83 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X684 a_6996_7663.t3 a_6081_7663.t2 a_6649_7905.t1 VSSD.t333 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X685 VDDD.t1046 VSSD.t1895 VDDD.t1045 VDDD.t1044 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X686 clknet_1_0__leaf_CLK.t7 a_7654_4943.t19 VSSD.t285 VSSD.t284 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X687 a_10838_3677.t0 a_9761_3311.t4 a_10676_3311.t0 VDDD.t1203 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X688 VDDD.t330 a_10145_9269.t4 a_10035_9295.t1 VDDD.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X689 a_8362_10927.t1 EN.t25 VSSD.t505 VSSD.t504 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X690 VDDD.t687 x2/net7.t4 a_3158_10205.t1 VDDD.t686 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X691 VSSD.t1445 VDDD.t2024 VSSD.t1444 VSSD.t1443 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X692 a_7618_8207.t0 a_6541_8213.t3 a_7456_8585.t2 VDDD.t1102 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X693 VDDD.t172 a_5147_11989.t6 a_5134_12381.t0 VDDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X694 a_8339_6603.t2 FINAL.t17 VDDD.t622 VDDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X695 a_4146_9003.t1 a_4424_9019.t3 a_4380_9117.t1 VDDD.t1560 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X696 VDDD.t336 CLKS.t57 a_2556_4943.t2 VDDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X697 SWP[9].t3 a_4779_5461.t4 VSSD.t838 VSSD.t837 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X698 a_9464_7485.t3 SWP[3].t4 VSSD.t109 VSSD.t108 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X699 a_3158_4765.t3 a_2439_4541.t4 a_2595_4636.t3 VSSD.t1620 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X700 VDDD.t876 a_5340_4233.t5 a_5515_4159.t2 VDDD.t875 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X701 a_2372_9117.t1 a_2158_9117.t4 VDDD.t270 VDDD.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X702 a_7563_2741.t1 a_7368_2883.t3 a_7873_3133.t1 VSSD.t985 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X703 a_9832_9661.t3 SWP[0].t5 VSSD.t1133 VSSD.t901 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X704 VSSD.t1442 VDDD.t2025 VSSD.t1441 VSSD.t1440 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X705 VSSD.t1439 VDDD.t2026 VSSD.t1438 VSSD.t1437 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X706 VDDD.t1049 VSSD.t1896 VDDD.t1048 VDDD.t1047 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X707 VDDD.t1052 VSSD.t1897 VDDD.t1051 VDDD.t1050 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X708 a_7171_7637.t2 EN.t26 VDDD.t671 VDDD.t670 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X709 x2/net10.t1 a_3675_11775.t6 VDDD.t897 VDDD.t896 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X710 VSSD.t1436 VDDD.t2027 VSSD.t1435 VSSD.t1434 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X711 a_3500_11849.t2 a_2585_11477.t3 a_3153_11445.t1 VSSD.t1 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X712 a_6888_11837.t2 x2/net2.t4 VDDD.t93 VDDD.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X713 a_4929_8751.t1 a_4550_9117.t4 a_4857_8751.t1 VSSD.t1647 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X714 VDDD.t128 a_6077_9813.t22 clknet_1_1__leaf_CLK.t10 VDDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X715 VSSD.t1107 x3/COMP_BUF_P.t21 a_3158_4765.t2 VSSD.t1106 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X716 VDDD.t1451 x3/COMP_BUF_P.t22 a_3158_4765.t1 VDDD.t1450 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X717 VDDD.t636 a_10421_6817.t4 a_10311_6941.t2 VDDD.t635 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X718 VDDD.t338 CLKS.t58 a_6251_6549.t0 VDDD.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X719 clknet_0_CLK.t25 a_6813_7093.t18 VSSD.t193 VSSD.t192 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X720 x3/COMP_BUF_P.t12 a_8435_8181.t12 VSSD.t1830 VSSD.t1829 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X721 VDDD.t1305 a_8284_4233.t5 a_8459_4159.t2 VDDD.t1304 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X722 a_8170_11293.t1 a_7093_10927.t3 a_8008_10927.t1 VDDD.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X723 a_10032_8751.t3 a_8951_8751.t4 a_9685_8993.t2 VDDD.t1962 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X724 a_10601_9673.t0 a_9411_9301.t3 a_10492_9673.t1 VSSD.t139 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X725 a_6909_4399.t0 a_6743_4399.t3 VDDD.t1539 VDDD.t1538 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X726 a_8008_3311.t2 a_7093_3311.t4 a_7661_3553.t3 VSSD.t122 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X727 VSSD.t507 EN.t27 a_2157_7663.t1 VSSD.t506 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X728 a_7477_4641.t1 a_7259_4399.t4 VDDD.t771 VDDD.t770 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X729 x2/net13.t5 x2/net12.t5 VDDD.t1709 VDDD.t1708 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X730 VSSD.t407 a_3583_4917.t5 SWN[9].t2 VSSD.t406 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X731 VDDD.t236 a_6813_7093.t19 clknet_0_CLK.t11 VDDD.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X732 VSSD.t991 a_7563_8988.t4 a_7494_9117.t1 VSSD.t990 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X733 a_10016_3311.t2 CF[5].t4 VSSD.t31 VSSD.t30 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X734 a_5041_7663.t1 CLKS.t59 VSSD.t270 VSSD.t269 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X735 clknet_1_0__leaf_CLK.t8 a_7654_4943.t20 VDDD.t353 VDDD.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X736 VSSD.t36 CF[3].t7 a_7203_3861.t1 VSSD.t35 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X737 VDDD.t340 CLKS.t60 a_2924_6031.t1 VDDD.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X738 a_6573_6575.t1 a_6538_6827.t5 a_6251_6549.t1 VSSD.t488 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X739 VDDD.t1054 VSSD.t1898 VDDD.t1053 VDDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X740 a_7249_6575.t1 CLKS.t61 VSSD.t272 VSSD.t271 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X741 x2/net4.t3 a_8183_10901.t5 VSSD.t322 VSSD.t321 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X742 a_2564_10749.t2 x2/TRIG2.t2 VDDD.t1462 VDDD.t1461 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X743 VDDD.t812 a_9685_7905.t5 a_9575_8029.t0 VDDD.t811 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X744 a_1835_4373.t1 a_2122_4651.t4 VDDD.t1863 VDDD.t1862 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X745 VSSD.t1433 VDDD.t2028 VSSD.t1432 VSSD.t1431 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X746 VSSD.t287 a_7654_4943.t21 clknet_1_0__leaf_CLK.t9 VSSD.t286 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X747 VSSD.t1710 x2/net12.t6 x2/net13.t6 VSSD.t1709 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X748 a_2196_10927.t0 x2/net8.t4 VDDD.t588 VDDD.t587 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X749 a_9832_9839.t0 SWP[1].t4 VSSD.t902 VSSD.t901 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X750 a_5182_6941.t3 a_4463_6717.t3 a_4619_6812.t2 VSSD.t1690 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X751 VSSD.t465 clknet_1_0__leaf_CLK.t41 a_9687_6575.t1 VSSD.t464 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X752 VDDD.t1057 VSSD.t1899 VDDD.t1056 VDDD.t1055 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X753 a_9117_8751.t0 a_8951_8751.t5 VDDD.t1360 VDDD.t1359 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X754 a_7125_3133.t1 a_7090_2899.t5 a_6803_2741.t1 VSSD.t963 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X755 a_9117_7663.t1 a_8951_7663.t4 VSSD.t1703 VSSD.t1702 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X756 a_9559_7497.t2 a_9209_7125.t3 a_9464_7485.t1 VDDD.t1712 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X757 a_10846_5309.t0 CLKS.t62 VSSD.t274 VSSD.t273 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X758 a_5470_5853.t0 a_5383_5629.t3 a_5066_5739.t0 VDDD.t1265 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X759 VSSD.t1430 VDDD.t2029 VSSD.t1429 VSSD.t1428 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X760 VDDD.t1932 a_8100_6409.t5 a_8275_6335.t2 VDDD.t1931 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X761 a_10768_6575.t2 a_9853_6575.t3 a_10421_6817.t1 VSSD.t1757 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X762 VSSD.t950 a_10207_7637.t4 DOUT[4].t2 VSSD.t949 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X763 FINAL.t6 a_5307_7093.t9 VDDD.t147 VDDD.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X764 a_3197_11837.t0 a_3153_11445.t4 a_3031_11849.t0 VSSD.t1646 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X765 VSSD.t1427 VDDD.t2030 VSSD.t1426 VSSD.t1425 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X766 a_6633_11477.t0 a_6467_11477.t3 VDDD.t1301 VDDD.t1300 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X767 VSSD.t1424 VDDD.t2031 VSSD.t1423 VSSD.t1422 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X768 a_2564_10749.t3 x2/TRIG2.t3 VSSD.t1123 VSSD.t1122 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X769 a_5171_2741.t3 a_4976_2883.t3 a_5481_3133.t1 VSSD.t1134 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X770 VSSD.t542 a_2439_5629.t4 a_2400_5755.t1 VSSD.t541 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X771 a_4948_8029.t0 a_4734_8029.t4 VDDD.t145 VDDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X772 VSSD.t1763 a_4043_7637.t4 SWN[4].t2 VSSD.t1762 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X773 x2/net12.t0 x2/net6.t5 VDDD.t1616 VDDD.t1615 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X774 SWP[8].t3 a_1651_4917.t4 VSSD.t930 VSSD.t929 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X775 VSSD.t993 a_4411_11445.t4 x2/net1.t3 VSSD.t992 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X776 a_7937_3829.t3 a_7719_4233.t5 VDDD.t1736 VDDD.t1735 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X777 VSSD.t739 a_9287_10687.t5 a_9221_10761.t1 VSSD.t738 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X778 a_8435_8181.t3 COMP_P.t1 VSSD.t1102 VSSD.t1101 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X779 VSSD.t509 EN.t28 a_8809_10749.t1 VSSD.t508 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X780 VDDD.t681 a_2439_9981.t3 a_2400_10107.t1 VDDD.t680 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X781 SWN[9].t1 a_3583_4917.t6 VDDD.t548 VDDD.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X782 VSSD.t1756 a_10759_3071.t3 a_10693_3145.t0 VSSD.t1755 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X783 VDDD.t1559 a_7171_7637.t6 a_7158_8029.t1 VDDD.t1558 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X784 a_2372_8207.t0 a_2158_8207.t5 VDDD.t1917 VDDD.t1916 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X785 a_4826_10383.t1 a_4700_10499.t3 a_4422_10515.t2 VSSD.t1031 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X786 a_5090_8207.t1 a_4332_8323.t4 a_4527_8181.t2 VDDD.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X787 VSSD.t172 a_2595_7900.t5 a_2526_8029.t2 VSSD.t171 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X788 a_9667_7119.t0 a_9043_7125.t4 a_9559_7497.t1 VDDD.t1724 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X789 a_2029_8751.t1 a_1467_8725.t4 VSSD.t676 VSSD.t675 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X790 a_6053_3311.t0 CLKS.t63 VSSD.t890 VSSD.t889 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X791 a_9729_8751.t1 a_9685_8993.t4 a_9563_8751.t1 VSSD.t862 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X792 VSSD.t1109 x3/COMP_BUF_P.t23 a_6102_5853.t1 VSSD.t1108 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X793 VDDD.t1453 x3/COMP_BUF_P.t24 a_6102_5853.t0 VDDD.t1452 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X794 VDDD.t342 a_10676_5487.t4 a_10851_5461.t2 VDDD.t341 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X795 VDDD.t1059 VSSD.t1900 VDDD.t1058 VDDD.t1041 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X796 VSSD.t1421 VDDD.t2032 VSSD.t1420 VSSD.t1419 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X797 a_10219_3677.t2 a_9595_3311.t3 a_10111_3311.t2 VDDD.t1393 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X798 a_7105_7663.t0 a_5915_7663.t4 a_6996_7663.t0 VSSD.t728 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X799 a_8284_4233.t3 a_7203_3861.t2 a_7937_3829.t1 VDDD.t1432 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X800 VDDD.t28 clknet_0_CLK.t36 a_7654_4943.t2 VDDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X801 a_4857_6575.t0 CLKS.t64 VSSD.t892 VSSD.t891 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X802 a_4669_12015.t0 a_4625_12257.t5 a_4503_12015.t0 VSSD.t202 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X803 a_5619_11293.t2 a_4995_10927.t4 a_5511_10927.t2 VDDD.t824 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X804 FINAL.t5 a_5307_7093.t10 VDDD.t149 VDDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X805 VSSD.t1009 SWP[7].t4 a_2790_8207.t3 VSSD.t751 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X806 VSSD.t1418 VDDD.t2033 VSSD.t1417 VSSD.t1393 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X807 VDDD.t72 a_1835_5461.t5 SWN[7].t0 VDDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X808 VDDD.t1062 VSSD.t1901 VDDD.t1061 VDDD.t1060 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X809 a_3018_11293.t1 a_1941_10927.t3 a_2856_10927.t1 VDDD.t827 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X810 a_5409_3133.t1 CLKS.t65 VSSD.t894 VSSD.t893 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X811 a_2526_8029.t3 a_2400_7931.t3 a_2122_7915.t3 VSSD.t441 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X812 VSSD.t694 a_5055_3285.t6 CF[1].t2 VSSD.t693 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X813 VSSD.t1416 VDDD.t2034 VSSD.t1415 VSSD.t1414 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X814 x3/COMP_BUF_N.t5 a_7331_9269.t10 VDDD.t1549 VDDD.t1548 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X815 a_4779_5461.t1 a_5066_5739.t4 VDDD.t922 VDDD.t921 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X816 a_6527_7663.t1 a_6081_7663.t3 a_6431_7663.t2 VSSD.t334 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X817 SWN[3].t3 a_6803_8725.t4 VSSD.t292 VSSD.t291 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X818 a_4932_2767.t0 a_4411_2741.t5 VDDD.t703 VDDD.t702 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X819 VDDD.t574 CF[1].t7 a_6927_5487.t0 VDDD.t573 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X820 VSSD.t545 a_5147_11989.t7 x2/TRIG1.t2 VSSD.t544 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X821 a_9372_8751.t2 SWP[2].t4 VSSD.t1037 VSSD.t1036 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X822 a_5205_10749.t0 a_4826_10383.t4 a_5133_10749.t0 VSSD.t952 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X823 a_5102_2767.t0 a_5015_3009.t4 a_4698_2899.t0 VDDD.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X824 VSSD.t105 a_5307_7093.t11 FINAL.t13 VSSD.t104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X825 VDDD.t435 a_7948_7637.t10 clkload0.X.t2 VDDD.t434 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X826 VDDD.t1065 VSSD.t1902 VDDD.t1064 VDDD.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X827 VDDD.t536 a_4779_5461.t5 SWP[9].t1 VDDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X828 VDDD.t1068 VSSD.t1903 VDDD.t1067 VDDD.t1066 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X829 VDDD.t344 a_2509_11169.t5 a_2399_11293.t1 VDDD.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X830 VSSD.t1413 VDDD.t2035 VSSD.t1412 VSSD.t1411 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X831 VDDD.t1238 CLKS.t66 a_5684_5853.t1 VDDD.t1237 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X832 a_2439_4541.t0 CF[7].t4 VDDD.t903 VDDD.t902 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X833 a_7631_8511.t1 a_7456_8585.t5 a_7810_8573.t0 VSSD.t310 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X834 a_4932_11471.t1 a_4411_11445.t5 VDDD.t1335 VDDD.t1334 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X835 a_7350_7663.t1 EN.t29 VSSD.t511 VSSD.t510 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X836 VSSD.t896 CLKS.t67 a_5037_4221.t0 VSSD.t895 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X837 VDDD.t679 a_9685_11169.t4 a_9575_11293.t2 VDDD.t678 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X838 VDDD.t1070 VSSD.t1904 VDDD.t1069 VDDD.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X839 a_4463_6717.t0 CF[6].t5 VDDD.t1632 VDDD.t1631 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X840 a_8117_3311.t0 a_6927_3311.t4 a_8008_3311.t1 VSSD.t1773 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X841 a_10759_4159.t0 CLKS.t68 VDDD.t1240 VDDD.t1239 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X842 VDDD.t1574 CF[0].t8 a_7019_6037.t0 VDDD.t1573 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X843 VSSD.t513 EN.t30 a_3197_11837.t1 VSSD.t512 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X844 VDDD.t1711 x2/net12.t7 x2/net13.t7 VDDD.t1710 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X845 VDDD.t224 a_5171_2741.t4 a_5102_2767.t1 VDDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X846 VSSD.t1410 VDDD.t2036 VSSD.t1409 VSSD.t1408 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X847 a_4422_10515.t1 a_4739_10625.t5 a_4697_10749.t1 VSSD.t719 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X848 a_3153_11445.t2 a_2935_11849.t4 VDDD.t1286 VDDD.t1285 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X849 a_6983_11849.t2 a_6467_11477.t4 a_6888_11837.t1 VSSD.t517 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X850 VDDD.t1073 VSSD.t1905 VDDD.t1072 VDDD.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X851 VDDD.t1388 a_10759_3071.t4 a_10746_2767.t0 VDDD.t1387 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X852 VSSD.t749 a_4343_4917.t4 a_4274_4943.t1 VSSD.t748 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X853 a_4605_7663.t0 a_4043_7637.t5 VSSD.t1765 VSSD.t1764 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X854 a_4550_9117.t3 a_4463_8893.t4 a_4146_9003.t2 VDDD.t1552 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X855 clknet_1_1__leaf_CLK.t22 a_6077_9813.t23 VSSD.t89 VSSD.t88 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X856 VSSD.t1407 VDDD.t2037 VSSD.t1406 VSSD.t1405 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X857 a_2122_10091.t0 a_2400_10107.t3 a_2356_10205.t1 VDDD.t1533 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X858 a_9927_9839.t0 a_9411_9839.t3 a_9832_9839.t2 VSSD.t1023 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X859 VDDD.t118 a_4135_10357.t4 x2/net7.t0 VDDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X860 clkload0.X.t1 a_7948_7637.t11 VDDD.t437 VDDD.t436 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X861 VSSD.t1182 a_7331_9269.t11 x3/COMP_BUF_N.t13 VSSD.t1181 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X862 VSSD.t572 a_7999_4373.t4 SWP[2].t3 VSSD.t571 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X863 VSSD.t1404 VDDD.t2038 VSSD.t1403 VSSD.t1402 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X864 VSSD.t1401 VDDD.t2039 VSSD.t1400 VSSD.t1399 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X865 a_5511_10927.t3 a_4995_10927.t5 a_5416_10927.t2 VSSD.t1845 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X866 VSSD.t1398 VDDD.t2040 VSSD.t1397 VSSD.t1396 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X867 a_2411_4917.t3 a_2255_5185.t5 a_2556_4943.t1 VDDD.t1881 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X868 a_4503_12015.t1 a_4057_12015.t2 a_4407_12015.t3 VSSD.t1164 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X869 VDDD.t888 clknet_1_1__leaf_CLK.t35 a_6467_11477.t0 VDDD.t887 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X870 VDDD.t1076 VSSD.t1906 VDDD.t1075 VDDD.t1074 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X871 a_8362_3311.t1 CLKS.t69 VSSD.t898 VSSD.t897 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X872 x2/net8.t3 a_1835_9813.t4 VSSD.t307 VSSD.t306 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X873 VDDD.t1078 VSSD.t1907 VDDD.t1077 VDDD.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X874 VSSD.t148 CKO.t12 a_6375_8213.t0 VSSD.t147 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X875 VSSD.t1570 a_4463_8893.t5 a_4424_9019.t1 VSSD.t1569 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X876 CKO.t1 a_8339_6603.t3 VDDD.t829 VDDD.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X877 VDDD.t40 CF[5].t5 a_4259_3861.t0 VDDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X878 VDDD.t1081 VSSD.t1908 VDDD.t1080 VDDD.t1079 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X879 a_7873_3133.t0 a_7494_2767.t4 a_7801_3133.t0 VSSD.t635 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X880 a_8126_9117.t0 a_7407_8893.t5 a_7563_8988.t0 VSSD.t1695 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X881 VSSD.t1395 VDDD.t2041 VSSD.t1394 VSSD.t1393 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X882 a_10299_6575.t0 a_9853_6575.t4 a_10203_6575.t0 VSSD.t1758 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X883 a_7661_5729.t1 a_7443_5487.t4 VDDD.t1876 VDDD.t1875 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X884 a_10281_6397.t1 a_10237_6005.t5 a_10115_6409.t1 VSSD.t1156 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X885 VDDD.t1242 CLKS.t70 a_5316_2767.t1 VDDD.t1241 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X886 a_7365_3133.t1 a_6803_2741.t4 VSSD.t938 VSSD.t937 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X887 VSSD.t940 a_6803_2741.t5 CF[2].t1 VSSD.t939 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X888 a_5102_2767.t3 a_4976_2883.t4 a_4698_2899.t2 VSSD.t1746 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X889 VDDD.t940 x3/COMP_BUF_N.t23 a_5182_9117.t1 VDDD.t939 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X890 VDDD.t355 a_7654_4943.t22 clknet_1_0__leaf_CLK.t10 VDDD.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X891 a_3675_11775.t2 EN.t31 VDDD.t1471 VDDD.t1470 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X892 a_5746_3677.t0 a_5659_3453.t4 a_5342_3563.t1 VDDD.t805 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X893 a_10194_9117.t0 a_9117_8751.t4 a_10032_8751.t0 VDDD.t881 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X894 a_7348_10927.t0 x2/net3.t5 VDDD.t174 VDDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X895 VSSD.t1392 VDDD.t2042 VSSD.t1391 VSSD.t1390 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X896 a_10938_6397.t0 CLKS.t71 VSSD.t553 VSSD.t552 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X897 a_2974_4943.t3 a_2216_5059.t3 a_2411_4917.t1 VDDD.t1374 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X898 a_2071_8449.t0 CKO.t13 VDDD.t189 VDDD.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X899 VSSD.t1389 VDDD.t2043 VSSD.t1388 VSSD.t1387 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X900 a_5617_3311.t1 a_5055_3285.t7 VSSD.t696 VSSD.t695 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X901 VDDD.t1084 VSSD.t1909 VDDD.t1083 VDDD.t1082 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X902 VSSD.t1817 a_7723_11775.t4 x2/net3.t3 VSSD.t1816 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X903 VSSD.t764 x3/COMP_BUF_N.t24 a_8126_9117.t2 VSSD.t763 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X904 a_4463_6717.t1 CF[6].t6 VSSD.t1622 VSSD.t1621 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X905 VDDD.t1958 a_8435_8181.t13 x3/COMP_BUF_P.t4 VDDD.t1957 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X906 a_3859_8725.t1 a_4146_9003.t5 VDDD.t605 VDDD.t604 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X907 VDDD.t1520 a_7109_8181.t5 a_6999_8207.t2 VDDD.t1519 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X908 a_8454_6397.t0 CLKS.t72 VSSD.t555 VSSD.t554 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X909 VDDD.t1473 EN.t32 a_4135_10357.t2 VDDD.t1472 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X910 a_3043_11471.t2 EN.t33 VDDD.t1475 VDDD.t1474 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X911 VSSD.t557 CLKS.t73 a_8701_7457.t0 VSSD.t556 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X912 x3/COMP_BUF_P.t11 a_8435_8181.t14 VSSD.t1832 VSSD.t1831 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X913 VDDD.t191 CKO.t14 a_8951_7663.t0 VDDD.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X914 VSSD.t467 clknet_1_0__leaf_CLK.t42 a_9503_3861.t1 VSSD.t466 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X915 a_4146_4651.t3 a_4424_4667.t3 a_4380_4765.t1 VDDD.t866 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X916 a_7477_4641.t2 a_7259_4399.t5 VSSD.t612 VSSD.t611 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X917 VDDD.t1087 VSSD.t1910 VDDD.t1086 VDDD.t1085 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X918 a_10207_7637.t2 EN.t34 VDDD.t1477 VDDD.t1476 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X919 VDDD.t729 CLKS.t74 a_4764_9117.t0 VDDD.t728 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X920 VSSD.t559 CLKS.t75 a_3905_5309.t0 VSSD.t558 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X921 a_3675_11775.t0 a_3500_11849.t4 a_3854_11837.t0 VSSD.t379 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X922 a_4733_11837.t0 a_4698_11603.t4 a_4411_11445.t0 VSSD.t434 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X923 VDDD.t1090 VSSD.t1911 VDDD.t1089 VDDD.t1088 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X924 VDDD.t560 a_8008_5487.t4 a_8183_5461.t1 VDDD.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X925 VDDD.t1726 a_6855_6717.t4 a_6816_6843.t0 VDDD.t1725 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X926 a_4187_5185.t1 CF[9].t7 VSSD.t876 VSSD.t875 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X927 VDDD.t1370 a_5015_11713.t2 a_4976_11587.t0 VDDD.t1369 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X928 a_4973_3133.t1 a_4411_2741.t6 VSSD.t537 VSSD.t536 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X929 a_7654_4943.t1 clknet_0_CLK.t37 VDDD.t30 VDDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X930 VSSD.t1386 VDDD.t2044 VSSD.t1385 VSSD.t1384 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X931 VDDD.t1093 VSSD.t1912 VDDD.t1092 VDDD.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X932 VDDD.t920 SWP[8].t4 a_2790_9117.t2 VDDD.t919 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X933 a_3158_10205.t0 a_2439_9981.t4 a_2595_10076.t0 VSSD.t522 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X934 VDDD.t731 CLKS.t76 a_7708_9117.t0 VDDD.t730 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X935 SWP[1].t3 a_8183_5461.t5 VSSD.t922 VSSD.t921 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X936 a_5383_5629.t1 CF[9].t8 VSSD.t878 VSSD.t877 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X937 a_7753_6005.t3 a_7535_6409.t4 VSSD.t1616 VSSD.t1615 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X938 VDDD.t1919 a_7723_11775.t5 a_7710_11471.t1 VDDD.t1918 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X939 VDDD.t238 a_6813_7093.t20 clknet_0_CLK.t10 VDDD.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X940 a_9667_7119.t1 EN.t35 VDDD.t1479 VDDD.t1478 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X941 a_10492_9839.t1 a_9411_9839.t4 a_10145_10081.t0 VDDD.t1261 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X942 a_2537_8751.t1 a_2158_9117.t5 a_2465_8751.t0 VSSD.t227 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X943 VDDD.t1095 VSSD.t1913 VDDD.t1094 VDDD.t1033 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X944 a_4672_8207.t2 a_4458_8207.t5 VDDD.t714 VDDD.t713 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X945 FINAL.t4 a_5307_7093.t12 VDDD.t151 VDDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X946 SWN[2].t0 a_4411_6005.t7 VDDD.t697 VDDD.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X947 VDDD.t78 a_10237_3829.t4 a_10127_3855.t0 VDDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X948 VSSD.t1383 VDDD.t2045 VSSD.t1382 VSSD.t1381 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X949 a_9575_11293.t0 a_8951_10927.t2 a_9467_10927.t2 VDDD.t1508 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X950 a_2877_10357.t3 a_2659_10761.t4 VDDD.t842 VDDD.t841 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X951 VSSD.t526 x2/net7.t5 a_3158_10205.t2 VSSD.t525 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X952 VDDD.t1098 VSSD.t1914 VDDD.t1097 VDDD.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X953 a_10032_10927.t1 a_8951_10927.t3 a_9685_11169.t0 VDDD.t1509 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X954 a_2356_10205.t0 a_1835_9813.t5 VDDD.t1218 VDDD.t1217 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X955 VSSD.t1080 a_10299_7423.t6 a_10233_7497.t0 VSSD.t1079 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X956 x3/COMP_BUF_N.t4 a_7331_9269.t12 VDDD.t1551 VDDD.t1550 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X957 a_1467_8725.t1 a_1754_9003.t5 VDDD.t427 VDDD.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X958 a_5619_11293.t1 EN.t36 VDDD.t1481 VDDD.t1480 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X959 clknet_1_1__leaf_CLK.t21 a_6077_9813.t24 VSSD.t91 VSSD.t90 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X960 VSSD.t1750 a_2255_5185.t6 a_2216_5059.t1 VSSD.t1749 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X961 VDDD.t1738 VSSD.t1915 VDDD.t1737 VDDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X962 a_10023_5321.t1 a_9577_4949.t2 a_9927_5321.t2 VSSD.t604 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X963 VSSD.t107 a_5307_7093.t13 FINAL.t12 VSSD.t106 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X964 a_2833_7663.t1 EN.t37 VSSD.t1132 VSSD.t1131 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X965 VSSD.t561 CLKS.t77 a_7705_5487.t0 VSSD.t560 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X966 VSSD.t981 a_10667_9599.t6 a_10601_9673.t1 VSSD.t980 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X967 a_4421_4399.t1 a_3859_4373.t5 VSSD.t828 VSSD.t827 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X968 a_5134_12381.t1 a_4057_12015.t3 a_4972_12015.t3 VDDD.t1525 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X969 VDDD.t1741 VSSD.t1916 VDDD.t1740 VDDD.t1739 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X970 a_10189_9661.t0 a_10145_9269.t5 a_10023_9673.t1 VSSD.t268 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X971 a_10141_10927.t0 a_8951_10927.t4 a_10032_10927.t0 VSSD.t1149 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X972 a_7443_10927.t0 a_6927_10927.t3 a_7348_10927.t3 VSSD.t1793 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X973 a_5316_11471.t0 a_5102_11471.t5 VDDD.t157 VDDD.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X974 VSSD.t1380 VDDD.t2046 VSSD.t1379 VSSD.t1378 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X975 VDDD.t1288 a_10207_7637.t5 a_10194_8029.t0 VDDD.t1287 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X976 a_4647_7805.t0 CF[4].t6 VDDD.t800 VDDD.t799 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X977 VDDD.t95 a_10145_10081.t4 a_10035_10205.t1 VDDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X978 VSSD.t1047 a_10759_3071.t5 CF[3].t3 VSSD.t1046 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X979 VDDD.t1743 VSSD.t1917 VDDD.t1742 VDDD.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X980 a_10108_6575.t2 EN.t38 VDDD.t214 VDDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X981 VSSD.t163 EN.t39 a_7153_8573.t0 VSSD.t162 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X982 VSSD.t1744 a_4647_7805.t5 a_4608_7931.t1 VSSD.t1743 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X983 a_9927_5321.t3 a_9577_4949.t3 a_9832_5309.t3 VDDD.t345 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X984 a_5171_11445.t1 a_4976_11587.t3 a_5481_11837.t0 VSSD.t433 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X985 VDDD.t1912 a_9112_10761.t4 a_9287_10687.t1 VDDD.t1911 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X986 a_10759_6335.t1 a_10584_6409.t4 a_10938_6397.t1 VSSD.t1008 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X987 a_9729_10927.t1 a_9685_11169.t5 a_9563_10927.t1 VSSD.t185 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X988 a_5539_5724.t1 a_5383_5629.t4 a_5684_5853.t2 VDDD.t206 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X989 a_2740_8029.t0 a_2526_8029.t4 VDDD.t122 VDDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X990 clknet_0_CLK.t24 a_6813_7093.t21 VSSD.t798 VSSD.t797 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X991 VSSD.t1173 a_1835_7637.t5 DOUT[9].t2 VSSD.t1172 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X992 a_4329_8573.t1 a_3767_8181.t6 VSSD.t7 VSSD.t6 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X993 VSSD.t1754 a_7563_2741.t5 a_7494_2767.t3 VSSD.t1753 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X994 CF[8].t1 a_10759_6335.t6 VSSD.t86 VSSD.t85 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X995 a_7824_4399.t0 a_6909_4399.t3 a_7477_4641.t0 VSSD.t471 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X996 a_10943_6549.t2 a_10768_6575.t5 a_11122_6575.t1 VSSD.t1175 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X997 a_3031_10901.t2 EN.t40 VDDD.t216 VDDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X998 VDDD.t870 a_6251_10901.t6 a_6238_11293.t0 VDDD.t869 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X999 clknet_0_CLK.t9 a_6813_7093.t22 VDDD.t964 VDDD.t963 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1000 VSSD.t1377 VDDD.t2047 VSSD.t1376 VSSD.t1301 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1001 a_7999_4373.t2 CLKS.t78 VDDD.t733 VDDD.t732 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1002 a_6431_7663.t3 a_6081_7663.t4 a_6336_7663.t1 VDDD.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1003 VSSD.t1136 a_6855_6717.t5 a_6816_6843.t1 VSSD.t1135 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1004 VDDD.t1214 SWP[7].t5 a_2790_8207.t2 VDDD.t1213 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1005 VDDD.t1746 VSSD.t1918 VDDD.t1745 VDDD.t1744 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1006 VSSD.t888 a_8275_6335.t6 SWP[0].t2 VSSD.t887 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1007 clknet_0_CLK.t23 a_6813_7093.t23 VSSD.t800 VSSD.t799 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1008 VSSD.t1644 a_10667_9813.t5 a_10601_9839.t1 VSSD.t980 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1009 a_9924_3133.t1 CF[4].t7 VSSD.t628 VSSD.t627 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1010 a_5773_10927.t0 a_5729_11169.t4 a_5607_10927.t0 VSSD.t12 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1011 VDDD.t1749 VSSD.t1919 VDDD.t1748 VDDD.t1747 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1012 VSSD.t353 a_10851_3285.t6 a_10785_3311.t1 VSSD.t352 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1013 a_9669_2773.t1 a_9503_2773.t4 VSSD.t1767 VSSD.t1766 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1014 VSSD.t1375 VDDD.t2048 VSSD.t1374 VSSD.t1373 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1015 a_10189_9839.t0 a_10145_10081.t5 a_10023_9839.t0 VSSD.t268 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1016 VSSD.t1628 a_7331_9269.t13 x3/COMP_BUF_N.t12 VSSD.t1627 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1017 VDDD.t1752 VSSD.t1920 VDDD.t1751 VDDD.t1750 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1018 VDDD.t1754 VSSD.t1921 VDDD.t1753 VDDD.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1019 VDDD.t1564 a_6803_8725.t5 SWN[3].t1 VDDD.t1563 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1020 VSSD.t1372 VDDD.t2049 VSSD.t1371 VSSD.t1370 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1021 VSSD.t165 EN.t41 a_9729_7663.t1 VSSD.t164 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1022 VSSD.t414 a_7407_3009.t6 a_7368_2883.t1 VSSD.t413 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1023 a_5102_11471.t1 a_5015_11713.t3 a_4698_11603.t2 VDDD.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1024 a_10373_3311.t1 a_10329_3553.t4 a_10207_3311.t1 VSSD.t979 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1025 a_10141_7663.t1 a_8951_7663.t5 a_10032_7663.t3 VSSD.t881 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1026 DOUT[0].t2 a_10667_9599.t7 VSSD.t983 VSSD.t982 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1027 a_10329_5729.t0 a_10111_5487.t5 VSSD.t456 VSSD.t455 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1028 VSSD.t715 a_6251_10901.t7 x2/net2.t3 VSSD.t714 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1029 a_6633_11477.t1 a_6467_11477.t5 VSSD.t519 VSSD.t518 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1030 a_8126_2767.t2 a_7368_2883.t4 a_7563_2741.t0 VDDD.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1031 SWP[6].t2 a_3859_4373.t6 VSSD.t830 VSSD.t829 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1032 DOUT[5].t0 a_7631_8511.t6 VDDD.t1309 VDDD.t1308 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1033 VSSD.t1661 CLKS.t79 a_2157_4399.t0 VSSD.t1660 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1034 VSSD.t1663 CLKS.t80 a_10189_5309.t0 VSSD.t1662 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1035 a_1467_8181.t1 a_1754_8339.t4 VDDD.t1580 VDDD.t1579 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1036 DOUT[4].t1 a_10207_7637.t6 VDDD.t1290 VDDD.t1289 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1037 VSSD.t1369 VDDD.t2050 VSSD.t1368 VSSD.t1367 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1038 VDDD.t859 a_4619_8988.t4 a_4550_9117.t1 VDDD.t858 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1039 a_8459_4159.t0 CLKS.t81 VDDD.t1665 VDDD.t1664 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1040 a_4043_7637.t1 a_4330_7915.t5 VDDD.t452 VDDD.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1041 a_7407_8893.t1 CF[3].t8 VSSD.t711 VSSD.t710 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1042 a_10386_7663.t0 EN.t42 VSSD.t167 VSSD.t166 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1043 a_7369_3861.t0 a_7203_3861.t3 VDDD.t1434 VDDD.t1433 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1044 SWN[4].t1 a_4043_7637.t6 VDDD.t1885 VDDD.t1884 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1045 VSSD.t1366 VDDD.t2051 VSSD.t1365 VSSD.t1364 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1046 x3/COMP_BUF_P.t3 a_8435_8181.t15 VDDD.t1960 VDDD.t1959 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1047 VDDD.t130 a_6077_9813.t25 clknet_1_1__leaf_CLK.t9 VDDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1048 CLKS.t11 x2/net13.t14 VSSD.t1015 VSSD.t1014 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1049 a_10676_3311.t3 a_9595_3311.t4 a_10329_3553.t3 VDDD.t1460 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1050 a_4488_4943.t1 a_4274_4943.t5 VDDD.t773 VDDD.t772 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1051 a_5539_5724.t3 a_5344_5755.t4 a_5849_5487.t1 VSSD.t580 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1052 x2/net1.t2 a_4411_11445.t6 VSSD.t995 VSSD.t994 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1053 a_2387_10927.t0 a_1941_10927.t4 a_2291_10927.t3 VSSD.t1819 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1054 a_10032_10927.t2 a_9117_10927.t3 a_9685_11169.t3 VSSD.t1028 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1055 a_9559_7497.t0 a_9043_7125.t5 a_9464_7485.t0 VSSD.t636 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1056 VDDD.t1331 a_7563_8988.t5 a_7494_9117.t2 VDDD.t1330 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1057 VDDD.t132 a_6077_9813.t26 clknet_1_1__leaf_CLK.t8 VDDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1058 VSSD.t1363 VDDD.t2052 VSSD.t1362 VSSD.t1272 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1059 a_8765_10357.t2 a_8547_10761.t4 VDDD.t1329 VDDD.t1328 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1060 VSSD.t1361 VDDD.t2053 VSSD.t1360 VSSD.t1263 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1061 a_7259_4399.t1 a_6743_4399.t4 a_7164_4399.t3 VSSD.t1174 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1062 VDDD.t558 a_4803_7900.t4 a_4734_8029.t0 VDDD.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1063 a_8547_10761.t3 a_8031_10389.t2 a_8452_10749.t3 VSSD.t1811 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1064 DOUT[8].t0 a_1467_8725.t5 VDDD.t840 VDDD.t839 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1065 a_2158_9117.t1 a_2071_8893.t3 a_1754_9003.t0 VDDD.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1066 VDDD.t1667 CLKS.t82 a_3767_8181.t0 VDDD.t1666 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1067 a_4371_8449.t1 CF[5].t6 VDDD.t42 VDDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1068 a_1754_9003.t2 a_2071_8893.t4 a_2029_8751.t0 VSSD.t523 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1069 a_5694_4221.t0 CLKS.t83 VSSD.t1665 VSSD.t1664 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1070 VSSD.t1667 CLKS.t84 a_4181_6575.t0 VSSD.t1666 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1071 VSSD.t199 a_8459_4159.t4 SWP[3].t3 VSSD.t198 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1072 a_7654_4943.t7 clknet_0_CLK.t38 VSSD.t15 VSSD.t14 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1073 a_9372_8751.t3 SWP[2].t5 VDDD.t1376 VDDD.t1375 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1074 VSSD.t772 a_2595_4636.t4 a_2526_4765.t1 VSSD.t771 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1075 a_9685_8993.t1 a_9467_8751.t4 VDDD.t466 VDDD.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1076 VSSD.t1111 x3/COMP_BUF_P.t25 a_5734_2767.t1 VSSD.t1110 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1077 a_2411_4917.t0 a_2216_5059.t4 a_2721_5309.t1 VSSD.t119 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1078 VDDD.t1757 VSSD.t1922 VDDD.t1756 VDDD.t1755 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1079 a_4550_4765.t2 a_4463_4541.t5 a_4146_4651.t1 VDDD.t1188 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1080 VSSD.t1359 VDDD.t2054 VSSD.t1358 VSSD.t1357 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1081 a_2439_7805.t1 CKO.t15 VSSD.t1835 VSSD.t1834 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1082 a_2779_6005.t0 a_2623_6273.t6 a_2924_6031.t2 VDDD.t863 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1083 a_2595_4636.t2 a_2439_4541.t5 a_2740_4765.t2 VDDD.t1626 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1084 VDDD.t765 a_7654_4943.t23 clknet_1_0__leaf_CLK.t17 VDDD.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1085 VSSD.t681 a_2071_8893.t5 a_2032_9019.t1 VSSD.t344 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1086 VSSD.t169 EN.t43 a_5773_10927.t1 VSSD.t168 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1087 a_3870_5075.t0 a_4187_5185.t4 a_4145_5309.t1 VSSD.t1126 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1088 SWP[5].t0 a_5515_4159.t7 VDDD.t707 VDDD.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1089 VSSD.t469 clknet_1_0__leaf_CLK.t43 a_9595_5487.t1 VSSD.t468 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1090 a_10299_7423.t0 a_10124_7497.t4 a_10478_7485.t0 VSSD.t346 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1091 a_2921_10749.t0 a_2877_10357.t5 a_2755_10761.t0 VSSD.t936 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1092 a_9287_10687.t2 EN.t44 VDDD.t218 VDDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1093 a_2122_5739.t2 a_2400_5755.t3 a_2356_5853.t1 VDDD.t908 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1094 a_10693_4233.t0 a_9503_3861.t4 a_10584_4233.t1 VSSD.t1577 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1095 VDDD.t36 clknet_0_CLK.t39 a_7654_4943.t0 VDDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1096 SWN[6].t0 a_3859_6549.t6 VDDD.t1106 VDDD.t1105 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1097 VDDD.t890 clknet_1_1__leaf_CLK.t36 a_2419_11477.t0 VDDD.t889 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1098 a_10676_5487.t1 a_9761_5487.t3 a_10329_5729.t1 VSSD.t535 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1099 a_10584_3145.t0 a_9669_2773.t2 a_10237_2741.t0 VSSD.t472 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1100 a_10667_9599.t0 a_10492_9673.t4 a_10846_9661.t0 VSSD.t435 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1101 a_2526_4765.t0 a_2400_4667.t3 a_2122_4651.t0 VSSD.t225 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1102 a_7551_3677.t1 CLKS.t85 VDDD.t1669 VDDD.t1668 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1103 a_4104_4943.t0 a_3583_4917.t7 VDDD.t550 VDDD.t549 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1104 clknet_0_CLK.t8 a_6813_7093.t24 VDDD.t966 VDDD.t965 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1105 VDDD.t1760 VSSD.t1923 VDDD.t1759 VDDD.t1758 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1106 VSSD.t1356 VDDD.t2055 VSSD.t1355 VSSD.t1354 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1107 FINAL.t3 a_5307_7093.t14 VDDD.t153 VDDD.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1108 VDDD.t899 a_3675_11775.t7 x2/net10.t0 VDDD.t898 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1109 a_10035_10205.t0 a_9411_9839.t5 a_9927_9839.t1 VDDD.t1262 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1110 a_3342_6031.t3 a_2584_6147.t5 a_2779_6005.t3 VDDD.t954 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1111 VSSD.t746 x3/COMP_BUF_P.t26 a_5182_4765.t1 VSSD.t745 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1112 VDDD.t911 x3/COMP_BUF_P.t27 a_5182_4765.t0 VDDD.t910 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1113 a_3158_4765.t0 a_2400_4667.t4 a_2595_4636.t1 VDDD.t268 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1114 x3/COMP_BUF_N.t3 a_7331_9269.t14 VDDD.t1636 VDDD.t1635 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1115 VDDD.t1516 a_4972_12015.t5 a_5147_11989.t2 VDDD.t1515 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1116 VDDD.t1763 VSSD.t1924 VDDD.t1762 VDDD.t1761 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1117 a_8435_8181.t4 COMP_P.t2 VSSD.t1104 VSSD.t1103 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1118 VDDD.t1445 a_8183_10901.t6 a_8170_11293.t0 VDDD.t1444 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1119 VDDD.t1766 VSSD.t1925 VDDD.t1765 VDDD.t1764 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1120 x2/net13.t0 x2/net12.t8 VDDD.t814 VDDD.t813 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1121 VSSD.t794 a_10943_6549.t5 CF[9].t2 VSSD.t793 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1122 VDDD.t1769 VSSD.t1926 VDDD.t1768 VDDD.t1767 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1123 a_10023_9673.t0 a_9577_9301.t2 a_9927_9673.t2 VSSD.t532 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1124 x2/net2.t2 a_6251_10901.t8 VSSD.t717 VSSD.t716 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1125 VSSD.t48 x2/net11.t5 x2/TRIG2.t1 VSSD.t47 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1126 VDDD.t38 clknet_0_CLK.t40 a_6077_9813.t2 VDDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1127 a_2157_7663.t0 a_2122_7915.t4 a_1835_7637.t0 VSSD.t13 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1128 VSSD.t732 clknet_1_1__leaf_CLK.t37 a_6467_11477.t1 VSSD.t731 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1129 VDDD.t816 x2/net12.t9 x2/net13.t1 VDDD.t815 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1130 VDDD.t1772 VSSD.t1927 VDDD.t1771 VDDD.t1770 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1131 a_4619_6812.t3 a_4463_6717.t4 a_4764_6941.t1 VDDD.t1683 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1132 DOUT[3].t0 a_10299_7423.t7 VDDD.t1418 VDDD.t1417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1133 a_8183_3285.t0 CLKS.t86 VDDD.t1671 VDDD.t1670 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1134 a_3859_4373.t1 a_4146_4651.t5 VDDD.t1212 VDDD.t1211 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1135 a_8615_7457.t2 FINAL.t18 VDDD.t624 VDDD.t623 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1136 a_2158_8207.t0 a_2071_8449.t3 a_1754_8339.t0 VDDD.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1137 VSSD.t409 a_8183_10901.t7 x2/net4.t2 VSSD.t408 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1138 a_6336_7663.t3 SWP[6].t4 VSSD.t624 VSSD.t623 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1139 a_9287_10687.t0 a_9112_10761.t5 a_9466_10749.t0 VSSD.t871 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1140 a_8209_6409.t1 a_7019_6037.t4 a_8100_6409.t0 VSSD.t2 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1141 a_10667_9813.t1 a_10492_9839.t5 a_10846_9839.t0 VSSD.t435 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1142 VDDD.t718 x2/net13.t15 CLKS.t0 VDDD.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1143 VDDD.t1774 VSSD.t1928 VDDD.t1773 VDDD.t1147 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1144 VDDD.t1185 a_3859_4373.t7 SWP[6].t1 VDDD.t1184 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1145 SWP[0].t1 a_8275_6335.t7 VDDD.t1234 VDDD.t1233 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1146 VDDD.t968 a_6813_7093.t25 clknet_0_CLK.t7 VDDD.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1147 a_3609_11849.t0 a_2419_11477.t3 a_3500_11849.t1 VSSD.t672 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1148 x2/net5.t0 a_9287_10687.t6 VDDD.t836 VDDD.t835 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1149 a_10492_5321.t3 a_9577_4949.t4 a_10145_4917.t3 VSSD.t451 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1150 VDDD.t1777 VSSD.t1929 VDDD.t1776 VDDD.t1775 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1151 VDDD.t272 CLKS.t87 a_4764_4765.t0 VDDD.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1152 VSSD.t1353 VDDD.t2056 VSSD.t1352 VSSD.t1351 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1153 VSSD.t802 a_6813_7093.t26 clknet_0_CLK.t22 VSSD.t801 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1154 SWP[4].t0 a_4411_2741.t7 VDDD.t705 VDDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1155 a_5307_7093.t0 CF[0].t9 VDDD.t1576 VDDD.t1575 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1156 VSSD.t804 a_6813_7093.t27 clknet_0_CLK.t21 VSSD.t803 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1157 VDDD.t1653 a_10667_9813.t6 DOUT[1].t1 VDDD.t1652 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1158 a_5182_6941.t0 a_4424_6843.t4 a_4619_6812.t0 VDDD.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1159 VDDD.t944 a_1467_8181.t5 DOUT[7].t1 VDDD.t943 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1160 VDDD.t618 a_2227_8181.t5 a_2158_8207.t2 VDDD.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1161 a_10111_3311.t3 a_9595_3311.t5 a_10016_3311.t3 VSSD.t1118 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1162 VDDD.t594 a_10943_6549.t6 a_10930_6941.t0 VDDD.t593 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1163 VSSD.t150 a_5307_7093.t15 FINAL.t11 VSSD.t149 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1164 clknet_1_1__leaf_CLK.t20 a_6077_9813.t27 VSSD.t93 VSSD.t92 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1165 a_4993_3829.t2 a_4775_4233.t4 VSSD.t735 VSSD.t734 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1166 VSSD.t229 CLKS.t88 a_10281_6397.t0 VSSD.t228 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1167 SWN[8].t0 a_2019_6005.t5 VDDD.t1970 VDDD.t1969 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1168 VDDD.t1618 x2/net6.t6 a_5458_10383.t0 VDDD.t1617 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1169 VDDD.t1780 VSSD.t1930 VDDD.t1779 VDDD.t1778 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1170 VSSD.t207 a_3399_10687.t6 a_3333_10761.t1 VSSD.t206 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1171 a_7631_6409.t1 a_7185_6037.t4 a_7535_6409.t3 VSSD.t709 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1172 VDDD.t274 CLKS.t89 a_4411_6005.t0 VDDD.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1173 VSSD.t1053 EN.t45 a_2921_10749.t1 VSSD.t1052 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1174 DOUT[7].t2 a_1467_8181.t6 VSSD.t769 VSSD.t342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1175 clknet_1_0__leaf_CLK.t18 a_7654_4943.t24 VSSD.t606 VSSD.t605 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1176 VSSD.t1350 VDDD.t2057 VSSD.t1349 VSSD.t1348 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1177 a_7348_3311.t3 CF[1].t8 VSSD.t425 VSSD.t424 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1178 a_1754_8339.t3 a_2071_8449.t4 a_2029_8573.t0 VSSD.t523 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1179 x2/net7.t3 a_4135_10357.t5 VSSD.t1713 VSSD.t1712 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1180 a_9821_7485.t0 a_9777_7093.t4 a_9655_7497.t1 VSSD.t1796 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1181 a_4619_6812.t1 a_4424_6843.t5 a_4929_6575.t0 VSSD.t678 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1182 VDDD.t1783 VSSD.t1931 VDDD.t1782 VDDD.t1781 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1183 VDDD.t1786 VSSD.t1932 VDDD.t1785 VDDD.t1784 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1184 a_8809_10749.t0 a_8765_10357.t4 a_8643_10761.t1 VSSD.t779 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1185 VDDD.t630 clknet_1_0__leaf_CLK.t44 a_9503_6037.t0 VDDD.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1186 VDDD.t663 a_8183_3285.t5 a_8170_3677.t1 VDDD.t662 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1187 x2/net11.t1 a_10207_10901.t5 VDDD.t564 VDDD.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1188 a_5481_6397.t0 a_5102_6031.t4 a_5409_6397.t1 VSSD.t761 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1189 SWN[7].t3 a_1835_5461.t6 VSSD.t44 VSSD.t43 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1190 VSSD.t1033 a_5015_11713.t4 a_4976_11587.t1 VSSD.t1032 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1191 a_7708_2767.t0 a_7494_2767.t5 VDDD.t809 VDDD.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1192 a_2342_4943.t0 a_2216_5059.t5 a_1938_5075.t2 VSSD.t120 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1193 VSSD.t1347 VDDD.t2058 VSSD.t1346 VSSD.t1231 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1194 a_5734_11471.t1 a_5015_11713.t5 a_5171_11445.t3 VSSD.t1034 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1195 VSSD.t1345 VDDD.t2059 VSSD.t1344 VSSD.t1343 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1196 a_4146_6827.t3 a_4463_6717.t5 a_4421_6575.t1 VSSD.t1691 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1197 a_9209_7125.t1 a_9043_7125.t6 VSSD.t638 VSSD.t637 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1198 a_10145_10081.t2 a_9927_9839.t5 VDDD.t1936 VDDD.t1935 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1199 a_4883_3855.t1 CLKS.t90 VDDD.t276 VDDD.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1200 a_10207_8725.t1 a_10032_8751.t5 a_10386_8751.t1 VSSD.t863 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1201 VSSD.t341 a_1467_8725.t6 DOUT[8].t3 VSSD.t340 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1202 a_9685_7905.t3 a_9467_7663.t5 VSSD.t1790 VSSD.t1789 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1203 VDDD.t1789 VSSD.t1933 VDDD.t1788 VDDD.t1787 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1204 VDDD.t1606 a_10667_5247.t7 CF[6].t0 VDDD.t1605 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1205 a_9577_9301.t1 a_9411_9301.t4 VSSD.t1022 VSSD.t919 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1206 VDDD.t1792 VSSD.t1934 VDDD.t1791 VDDD.t1790 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1207 VSSD.t381 COMP_N.t3 a_7331_9269.t3 VSSD.t380 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1208 VSSD.t1342 VDDD.t2060 VSSD.t1341 VSSD.t1340 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1209 a_9669_3861.t0 a_9503_3861.t5 VDDD.t1562 VDDD.t1561 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1210 a_4463_4541.t0 CF[6].t7 VDDD.t1634 VDDD.t1633 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1211 VSSD.t1339 VDDD.t2061 VSSD.t1338 VSSD.t1337 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1212 CF[7].t0 a_10851_5461.t5 VDDD.t1293 VDDD.t1292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1213 a_5147_11989.t0 EN.t46 VDDD.t1397 VDDD.t1396 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1214 a_7093_10927.t0 a_6927_10927.t4 VSSD.t1095 VSSD.t1094 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1215 a_7093_5487.t1 a_6927_5487.t5 VSSD.t112 VSSD.t111 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1216 a_10207_5487.t1 a_9761_5487.t4 a_10111_5487.t0 VSSD.t159 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1217 a_3854_11837.t1 EN.t47 VSSD.t1055 VSSD.t1054 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1218 a_10115_3145.t1 a_9669_2773.t3 a_10019_3145.t2 VSSD.t473 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1219 VDDD.t1399 EN.t48 a_2740_10205.t1 VDDD.t1398 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1220 a_7810_8573.t1 EN.t49 VSSD.t1057 VSSD.t1056 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1221 VDDD.t104 a_2439_7805.t4 a_2400_7931.t0 VDDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1222 VSSD.t1336 VDDD.t2062 VSSD.t1335 VSSD.t1334 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1223 VSSD.t23 clknet_0_CLK.t41 a_7654_4943.t6 VSSD.t22 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1224 a_2935_11849.t3 a_2585_11477.t4 a_2840_11837.t0 VDDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1225 a_4697_10749.t0 a_4135_10357.t6 VSSD.t1715 VSSD.t1714 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1226 a_2526_5853.t2 a_2439_5629.t5 a_2122_5739.t1 VDDD.t710 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1227 a_6888_11837.t3 x2/net2.t5 VSSD.t71 VSSD.t70 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1228 clknet_1_1__leaf_CLK.t7 a_6077_9813.t28 VDDD.t134 VDDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1229 a_10127_6031.t0 CLKS.t91 VDDD.t278 VDDD.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1230 VSSD.t33 CF[5].t7 a_4259_3861.t1 VSSD.t32 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1231 a_4421_8751.t0 a_3859_8725.t5 VSSD.t615 VSSD.t614 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1232 a_9927_9673.t3 a_9577_9301.t3 a_9832_9661.t0 VDDD.t1189 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1233 a_5066_5739.t1 a_5383_5629.t5 a_5341_5487.t0 VSSD.t160 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1234 a_7090_2899.t2 a_7407_3009.t7 a_7365_3133.t0 VSSD.t415 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1235 a_11030_5487.t0 CLKS.t92 VSSD.t231 VSSD.t230 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1236 a_4680_4221.t0 x3/COMP_BUF_P.t28 VDDD.t913 VDDD.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1237 clknet_1_0__leaf_CLK.t19 a_7654_4943.t25 VDDD.t767 VDDD.t766 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1238 a_10019_6409.t0 a_9669_6037.t4 a_9924_6397.t2 VDDD.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1239 a_5342_3563.t2 a_5620_3579.t3 a_5576_3677.t0 VDDD.t959 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1240 a_10311_6941.t1 CLKS.t93 VDDD.t280 VDDD.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1241 a_7093_10927.t1 a_6927_10927.t5 VDDD.t1438 VDDD.t1437 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1242 VSSD.t1059 EN.t50 a_4457_10749.t0 VSSD.t1058 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1243 x2/net8.t1 a_1835_9813.t6 VDDD.t1216 VDDD.t1215 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1244 VSSD.t1333 VDDD.t2063 VSSD.t1332 VSSD.t1321 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1245 a_6430_10927.t1 EN.t51 VSSD.t1061 VSSD.t1060 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1246 a_4993_3829.t0 a_4775_4233.t5 VDDD.t20 VDDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1247 a_9577_9839.t1 a_9411_9839.t6 VSSD.t920 VSSD.t919 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1248 VDDD.t1795 VSSD.t1935 VDDD.t1794 VDDD.t1793 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1249 VDDD.t1443 COMP_P.t3 a_8435_8181.t5 VDDD.t1442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1250 a_9761_3311.t1 a_9595_3311.t6 VSSD.t1120 VSSD.t1119 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1251 a_7324_2767.t1 a_6803_2741.t6 VDDD.t1279 VDDD.t1278 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1252 a_2581_6397.t0 a_2019_6005.t6 VSSD.t1842 VSSD.t1841 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1253 a_5015_6273.t0 CF[2].t6 VDDD.t1297 VDDD.t1296 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1254 VSSD.t1144 CLK.t2 a_6813_7093.t7 VSSD.t1143 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1255 VDDD.t282 CLKS.t94 a_2740_4765.t1 VDDD.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1256 VSSD.t1070 a_7948_7637.t12 clkload0.X.t14 VSSD.t1069 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1257 VDDD.t1649 a_4619_4636.t4 a_4550_4765.t0 VDDD.t1648 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1258 CF[4].t0 a_10851_3285.t7 VSSD.t355 VSSD.t354 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1259 VDDD.t1431 a_10124_7497.t5 a_10299_7423.t1 VDDD.t1430 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1260 a_3500_11849.t0 a_2419_11477.t4 a_3153_11445.t0 VDDD.t834 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1261 VDDD.t1499 a_6813_7093.t28 clknet_0_CLK.t6 VDDD.t1498 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1262 a_6431_7663.t0 a_5915_7663.t5 a_6336_7663.t0 VSSD.t729 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1263 VSSD.t490 EN.t52 a_2157_9839.t1 VSSD.t489 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1264 a_2833_4399.t1 CLKS.t95 VSSD.t237 VSSD.t236 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1265 a_3158_5853.t0 a_2439_5629.t6 a_2595_5724.t1 VSSD.t543 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1266 DOUT[9].t1 a_1835_7637.t6 VDDD.t1536 VDDD.t1535 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1267 DOUT[1].t2 a_10667_9813.t7 VSSD.t1645 VSSD.t982 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1268 a_5416_10927.t0 x2/net1.t4 VDDD.t1923 VDDD.t1922 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1269 a_8643_10761.t0 a_8197_10389.t3 a_8547_10761.t1 VSSD.t131 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1270 a_5340_4233.t1 a_4259_3861.t6 a_4993_3829.t1 VDDD.t542 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1271 a_5449_4233.t0 a_4259_3861.t7 a_5340_4233.t0 VSSD.t398 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1272 a_7156_6941.t0 a_6942_6941.t5 VDDD.t661 VDDD.t660 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1273 VDDD.t1798 VSSD.t1936 VDDD.t1797 VDDD.t1796 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1274 a_6909_4399.t1 a_6743_4399.t5 VSSD.t444 VSSD.t443 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1275 VDDD.t472 a_3500_11849.t5 a_3675_11775.t1 VDDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1276 a_7494_9117.t3 a_7368_9019.t3 a_7090_9003.t2 VSSD.t266 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1277 VDDD.t942 x3/COMP_BUF_N.t25 a_4906_4943.t1 VDDD.t941 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1278 a_10111_3311.t1 a_9761_3311.t5 a_10016_3311.t0 VDDD.t1204 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1279 x3/COMP_BUF_N.t2 a_7331_9269.t15 VDDD.t1638 VDDD.t1637 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1280 VSSD.t766 x3/COMP_BUF_N.t26 a_3158_5853.t3 VSSD.t765 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1281 VDDD.t1422 x3/COMP_BUF_N.t27 a_3158_5853.t2 VDDD.t1421 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1282 VSSD.t1045 a_6251_6549.t6 SWN[1].t2 VSSD.t1044 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1283 a_4312_12015.t3 x2/net10.t5 VSSD.t1741 VSSD.t1740 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1284 a_6102_5853.t2 a_5383_5629.t6 a_5539_5724.t0 VSSD.t161 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1285 a_10124_7497.t0 a_9209_7125.t4 a_9777_7093.t3 VSSD.t203 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1286 SWN[0].t2 a_3859_8725.t6 VSSD.t617 VSSD.t616 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1287 VDDD.t720 x2/net13.t16 CLKS.t1 VDDD.t719 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1288 a_10281_3133.t1 a_10237_2741.t5 a_10115_3145.t0 VSSD.t303 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1289 VSSD.t314 a_1835_4373.t6 SWP[7].t2 VSSD.t313 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1290 a_8393_4233.t1 a_7203_3861.t4 a_8284_4233.t1 VSSD.t297 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1291 a_8126_9117.t3 a_7368_9019.t4 a_7563_8988.t3 VDDD.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1292 a_7440_6397.t0 x3/COMP_BUF_P.t29 VDDD.t914 VDDD.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1293 VDDD.t1801 VSSD.t1937 VDDD.t1800 VDDD.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1294 a_6813_7093.t6 CLK.t3 VSSD.t359 VSSD.t358 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1295 VDDD.t468 a_3153_11445.t5 a_3043_11471.t1 VDDD.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1296 VSSD.t1331 VDDD.t2064 VSSD.t1330 VSSD.t1213 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1297 a_7259_4399.t3 a_6909_4399.t4 a_7164_4399.t2 VDDD.t1332 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1298 CF[3].t0 a_10759_3071.t6 VSSD.t1041 VSSD.t1040 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1299 x2/net3.t1 a_7723_11775.t6 VDDD.t1921 VDDD.t1920 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1300 a_10492_9673.t2 a_9577_9301.t4 a_10145_9269.t1 VSSD.t156 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1301 a_10938_3133.t0 CLKS.t96 VSSD.t239 VSSD.t238 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1302 VSSD.t1329 VDDD.t2065 VSSD.t1328 VSSD.t1327 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1303 VSSD.t241 CLKS.t97 a_10373_3311.t0 VSSD.t240 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1304 a_7753_6005.t2 a_7535_6409.t5 VDDD.t1436 VDDD.t1435 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1305 clknet_0_CLK.t5 a_6813_7093.t29 VDDD.t1501 VDDD.t1500 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1306 VDDD.t892 clknet_1_1__leaf_CLK.t38 a_8031_10389.t0 VDDD.t891 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1307 a_7443_3311.t0 a_6927_3311.t5 a_7348_3311.t0 VSSD.t1774 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1308 VDDD.t1206 a_9685_8993.t5 a_9575_9117.t2 VDDD.t1205 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1309 a_1835_5461.t1 a_2122_5739.t4 VDDD.t590 VDDD.t589 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1310 VDDD.t973 VSSD.t1938 VDDD.t972 VDDD.t971 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1311 VSSD.t1326 VDDD.t2066 VSSD.t1325 VSSD.t1324 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1312 clknet_0_CLK.t20 a_6813_7093.t30 VSSD.t1146 VSSD.t1145 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1313 VDDD.t975 VSSD.t1939 VDDD.t974 VDDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1314 a_2623_6273.t0 CF[8].t7 VDDD.t1645 VDDD.t1644 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1315 a_4458_8207.t2 a_4371_8449.t5 a_4054_8339.t0 VDDD.t1896 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1316 a_7815_4233.t1 a_7369_3861.t3 a_7719_4233.t0 VSSD.t733 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1317 a_10035_4943.t0 a_9411_4949.t5 a_9927_5321.t0 VDDD.t1458 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1318 a_6541_8213.t0 a_6375_8213.t5 VDDD.t221 VDDD.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1319 VSSD.t579 a_2595_10076.t5 a_2526_10205.t2 VSSD.t578 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1320 VDDD.t978 VSSD.t1940 VDDD.t977 VDDD.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1321 VDDD.t294 CLKS.t98 a_6803_2741.t0 VDDD.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1322 a_9117_8751.t1 a_8951_8751.t6 VSSD.t1020 VSSD.t1019 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1323 a_7407_3009.t0 clknet_1_0__leaf_CLK.t45 VDDD.t632 VDDD.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1324 VSSD.t534 a_4411_6005.t8 SWN[2].t2 VSSD.t533 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1325 a_7563_8988.t2 a_7368_9019.t5 a_7873_8751.t0 VSSD.t267 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1326 a_6538_6827.t2 a_6816_6843.t4 a_6772_6941.t1 VDDD.t1908 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1327 VSSD.t608 a_7654_4943.t26 clknet_1_0__leaf_CLK.t20 VSSD.t607 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1328 VSSD.t371 a_6077_9813.t29 clknet_1_1__leaf_CLK.t19 VSSD.t370 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1329 VSSD.t1772 a_10207_8725.t6 DOUT[2].t2 VSSD.t1771 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1330 a_7367_4765.t2 a_6743_4399.t6 a_7259_4399.t0 VDDD.t601 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1331 a_3905_5309.t1 a_3870_5075.t4 a_3583_4917.t1 VSSD.t1154 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1332 VSSD.t1323 VDDD.t2067 VSSD.t1322 VSSD.t1321 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1333 a_2721_5309.t0 a_2342_4943.t4 a_2649_5309.t0 VSSD.t114 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1334 a_10207_10901.t1 a_10032_10927.t5 a_10386_10927.t0 VSSD.t1026 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1335 VDDD.t894 clknet_1_1__leaf_CLK.t39 a_3891_12015.t0 VDDD.t893 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1336 a_8100_6409.t1 a_7019_6037.t5 a_7753_6005.t0 VDDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1337 VSSD.t1320 VDDD.t2068 VSSD.t1319 VSSD.t1318 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1338 a_7331_9269.t1 COMP_N.t4 VDDD.t210 VDDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1339 VDDD.t980 VSSD.t1941 VDDD.t979 VDDD.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1340 a_5015_11713.t0 clknet_1_1__leaf_CLK.t40 VDDD.t953 VDDD.t952 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1341 a_4764_6941.t2 a_4550_6941.t4 VDDD.t1696 VDDD.t1695 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1342 a_2213_5309.t1 a_1651_4917.t5 VSSD.t932 VSSD.t931 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1343 a_5777_5487.t1 CLKS.t99 VSSD.t243 VSSD.t242 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1344 a_7079_11849.t0 a_6633_11477.t4 a_6983_11849.t0 VSSD.t1027 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1345 a_4422_10515.t3 a_4700_10499.t4 a_4656_10383.t1 VDDD.t528 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1346 VSSD.t178 a_5015_6273.t6 a_4976_6147.t1 VSSD.t177 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1347 VDDD.t12 a_3767_8181.t7 SWN[5].t0 VDDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1348 VSSD.t547 x2/net13.t17 CLKS.t2 VSSD.t546 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1349 VSSD.t670 a_10759_4159.t5 a_10693_4233.t1 VSSD.t669 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1350 VDDD.t1941 a_4527_8181.t5 a_4458_8207.t0 VDDD.t1940 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1351 a_2740_10205.t2 a_2526_10205.t5 VDDD.t748 VDDD.t747 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1352 clknet_1_1__leaf_CLK.t6 a_6077_9813.t30 VDDD.t456 VDDD.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1353 VDDD.t382 a_2595_5724.t4 a_2526_5853.t0 VDDD.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1354 VSSD.t816 a_3859_6549.t7 SWN[6].t2 VSSD.t815 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1355 a_2540_6031.t0 a_2019_6005.t7 VDDD.t1972 VDDD.t1971 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1356 a_2526_10205.t0 a_2400_10107.t4 a_2122_10091.t1 VSSD.t1167 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1357 CF[0].t1 a_8183_3285.t6 VDDD.t665 VDDD.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1358 a_2356_4765.t1 a_1835_4373.t7 VDDD.t388 VDDD.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1359 CF[6].t2 a_10667_5247.t8 VSSD.t1601 VSSD.t1600 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1360 VSSD.t1317 VDDD.t2069 VSSD.t1316 VSSD.t1298 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1361 a_10851_5461.t1 a_10676_5487.t5 a_11030_5487.t1 VSSD.t401 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1362 VSSD.t1315 VDDD.t2070 VSSD.t1314 VSSD.t1313 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1363 VSSD.t789 a_4803_7900.t5 a_4734_8029.t2 VSSD.t788 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1364 a_8655_10383.t2 EN.t53 VDDD.t657 VDDD.t656 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1365 VDDD.t983 VSSD.t1942 VDDD.t982 VDDD.t981 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1366 a_2291_10927.t2 a_1941_10927.t5 a_2196_10927.t3 VDDD.t1942 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1367 VDDD.t16 a_5729_11169.t5 a_5619_11293.t0 VDDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1368 SWN[5].t2 a_3767_8181.t8 VSSD.t1840 VSSD.t1839 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1369 VDDD.t296 CLKS.t100 a_8339_6603.t0 VDDD.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1370 VSSD.t1312 VDDD.t2071 VSSD.t1311 VSSD.t1310 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1371 VSSD.t924 a_8183_5461.t6 a_8117_5487.t1 VSSD.t923 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1372 a_4054_8339.t1 a_4371_8449.t6 a_4329_8573.t0 VSSD.t1777 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1373 a_2595_7900.t3 a_2400_7931.t4 a_2905_7663.t1 VSSD.t1171 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1374 VSSD.t781 clknet_1_1__leaf_CLK.t41 a_2419_11477.t1 VSSD.t780 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1375 VSSD.t427 CF[1].t9 a_6927_5487.t1 VSSD.t426 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1376 DOUT[6].t2 a_7171_7637.t7 VSSD.t1575 VSSD.t1574 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1377 VDDD.t985 VSSD.t1943 VDDD.t984 VDDD.t511 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1378 a_10019_3145.t1 a_9503_2773.t5 a_9924_3133.t2 VSSD.t1768 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1379 VSSD.t1309 VDDD.t2072 VSSD.t1308 VSSD.t1307 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1380 VDDD.t659 EN.t54 a_5316_11471.t1 VDDD.t658 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1381 x3/COMP_BUF_P.t2 a_8435_8181.t16 VDDD.t924 VDDD.t923 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1382 VDDD.t946 a_2595_4636.t5 a_2526_4765.t2 VDDD.t945 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1383 a_7539_5487.t0 a_7093_5487.t3 a_7443_5487.t1 VSSD.t208 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1384 VDDD.t298 CLKS.t101 a_4411_2741.t0 VDDD.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1385 a_6813_6575.t0 a_6251_6549.t7 VSSD.t570 VSSD.t569 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1386 a_3224_10761.t0 a_2143_10389.t6 a_2877_10357.t1 VDDD.t1100 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1387 VDDD.t769 a_7654_4943.t27 clknet_1_0__leaf_CLK.t21 VDDD.t768 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1388 VDDD.t988 VSSD.t1944 VDDD.t987 VDDD.t986 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1389 a_7654_4943.t5 clknet_0_CLK.t42 VSSD.t25 VSSD.t24 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1390 a_10016_3311.t1 CF[5].t8 VDDD.t34 VDDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1391 VDDD.t244 a_6996_7663.t5 a_7171_7637.t1 VDDD.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1392 a_2526_10205.t3 a_2439_9981.t5 a_2122_10091.t2 VDDD.t1621 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1393 a_2439_4541.t1 CF[7].t5 VSSD.t742 VSSD.t741 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1394 a_2122_7915.t1 a_2439_7805.t5 a_2397_7663.t1 VSSD.t77 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1395 VSSD.t1084 x3/COMP_BUF_N.t28 a_5182_9117.t2 VSSD.t1083 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1396 a_4803_7900.t0 a_4647_7805.t6 a_4948_8029.t2 VDDD.t1879 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1397 a_7981_4221.t1 a_7937_3829.t5 a_7815_4233.t0 VSSD.t1025 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1398 VSSD.t1306 VDDD.t2073 VSSD.t1305 VSSD.t1304 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1399 VSSD.t755 a_8435_8181.t17 x3/COMP_BUF_P.t10 VSSD.t754 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1400 VDDD.t737 a_5015_3009.t5 a_4976_2883.t0 VDDD.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1401 SWP[3].t2 a_8459_4159.t5 VSSD.t201 VSSD.t200 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1402 a_4380_6941.t1 a_3859_6549.t8 VDDD.t1108 VDDD.t1107 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1403 VSSD.t703 a_2623_6273.t7 a_2584_6147.t1 VSSD.t702 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1404 VDDD.t85 a_3224_10761.t4 a_3399_10687.t0 VDDD.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1405 a_2439_5629.t1 CF[7].t6 VDDD.t905 VDDD.t904 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1406 CF[9].t0 a_10943_6549.t7 VDDD.t596 VDDD.t595 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1407 VSSD.t1086 x3/COMP_BUF_N.t29 a_3342_6031.t2 VSSD.t1085 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1408 VDDD.t938 a_2856_10927.t4 a_3031_10901.t0 VDDD.t937 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1409 a_6336_7663.t2 SWP[6].t5 VDDD.t796 VDDD.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1410 a_7624_4221.t1 x3/COMP_BUF_P.t30 VSSD.t363 VSSD.t362 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1411 VDDD.t991 VSSD.t1945 VDDD.t990 VDDD.t989 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1412 a_11122_6575.t0 CLKS.t102 VSSD.t245 VSSD.t244 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1413 VSSD.t783 clknet_1_1__leaf_CLK.t42 a_3891_12015.t1 VSSD.t782 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1414 a_7369_3861.t1 a_7203_3861.t5 VSSD.t299 VSSD.t298 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1415 VDDD.t300 CLKS.t103 a_2019_6005.t0 VDDD.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1416 a_10759_3071.t0 a_10584_3145.t4 a_10938_3133.t1 VSSD.t67 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1417 VDDD.t576 clknet_1_0__leaf_CLK.t46 a_9595_3311.t0 VDDD.t575 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1418 VDDD.t302 CLKS.t104 a_1835_4373.t0 VDDD.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1419 VSSD.t970 a_7631_8511.t7 DOUT[5].t2 VSSD.t969 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1420 a_5366_8029.t1 a_4608_7931.t3 a_4803_7900.t2 VDDD.t1604 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1421 VDDD.t1319 a_10329_3553.t5 a_10219_3677.t1 VDDD.t1318 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1422 a_9927_5321.t1 a_9411_4949.t6 a_9832_5309.t0 VSSD.t1117 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1423 a_5133_10749.t1 EN.t55 VSSD.t492 VSSD.t491 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1424 a_3089_6397.t0 a_2710_6031.t5 a_3017_6397.t0 VSSD.t1176 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1425 a_9563_7663.t0 a_9117_7663.t3 a_9467_7663.t1 VSSD.t431 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1426 VSSD.t574 a_7999_4373.t5 a_7933_4399.t0 VSSD.t573 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1427 VDDD.t32 a_10759_4159.t6 a_10746_3855.t0 VDDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1428 a_2790_9117.t1 a_2071_8893.t6 a_2227_8988.t3 VSSD.t524 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1429 a_9832_9839.t1 SWP[1].t5 VDDD.t1244 VDDD.t1243 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1430 VSSD.t1303 VDDD.t2074 VSSD.t1302 VSSD.t1301 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1431 VSSD.t1300 VDDD.t2075 VSSD.t1299 VSSD.t1298 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1432 VSSD.t494 EN.t56 a_7245_11837.t1 VSSD.t493 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1433 a_3043_11471.t0 a_2419_11477.t5 a_2935_11849.t1 VDDD.t1282 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1434 a_2157_4399.t1 a_2122_4651.t5 a_1835_4373.t2 VSSD.t1726 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1435 a_1754_9003.t1 a_2032_9019.t3 a_1988_9117.t0 VDDD.t807 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1436 a_7443_3311.t3 a_7093_3311.t5 a_7348_3311.t1 VDDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1437 a_5734_6031.t3 a_5015_6273.t7 a_5171_6005.t2 VSSD.t179 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1438 VSSD.t934 a_1651_4917.t6 SWP[8].t2 VSSD.t933 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1439 VSSD.t1297 VDDD.t2076 VSSD.t1296 VSSD.t1295 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1440 a_7661_11169.t0 a_7443_10927.t4 VDDD.t240 VDDD.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1441 a_7565_8585.t0 a_6375_8213.t6 a_7456_8585.t0 VSSD.t170 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1442 a_9466_10749.t1 EN.t57 VSSD.t496 VSSD.t495 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1443 a_9372_10927.t1 x2/net5.t5 VDDD.t1196 VDDD.t1195 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1444 a_7201_11445.t0 a_6983_11849.t4 VDDD.t404 VDDD.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1445 VDDD.t552 a_3583_4917.t8 SWN[9].t0 VDDD.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1446 VSSD.t752 SWP[8].t5 a_2790_9117.t3 VSSD.t751 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1447 VDDD.t1441 a_5171_11445.t4 a_5102_11471.t2 VDDD.t1440 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1448 a_5502_3855.t0 a_4425_3861.t4 a_5340_4233.t3 VDDD.t1944 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1449 VSSD.t1698 a_5171_6005.t5 a_5102_6031.t3 VSSD.t1697 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1450 VDDD.t578 clknet_1_0__leaf_CLK.t47 a_9411_4949.t0 VDDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1451 VDDD.t1299 CF[2].t7 a_6378_3677.t0 VDDD.t1298 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1452 a_10127_2767.t0 CLKS.t105 VDDD.t304 VDDD.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1453 CKO.t2 a_8615_7457.t4 VSSD.t959 VSSD.t958 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1454 DOUT[1].t0 a_10667_9813.t8 VDDD.t1655 VDDD.t1654 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1455 a_4656_10383.t0 a_4135_10357.t7 VDDD.t1714 VDDD.t1713 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1456 VDDD.t993 VSSD.t1946 VDDD.t992 VDDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1457 clknet_1_1__leaf_CLK.t18 a_6077_9813.t31 VSSD.t373 VSSD.t372 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1458 a_8547_10761.t2 a_8197_10389.t4 a_8452_10749.t0 VDDD.t178 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1459 a_10019_3145.t3 a_9669_2773.t4 a_9924_3133.t3 VDDD.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1460 VDDD.t251 a_3399_10687.t7 x2/net6.t1 VDDD.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1461 VSSD.t1294 VDDD.t2077 VSSD.t1293 VSSD.t1292 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1462 a_6987_8585.t0 a_6541_8213.t4 a_6891_8585.t3 VSSD.t98 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1463 a_9221_10761.t0 a_8031_10389.t3 a_9112_10761.t0 VSSD.t100 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1464 VDDD.t306 CLKS.t106 a_3859_6549.t0 VDDD.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1465 a_7164_4399.t1 x3/COMP_BUF_P.t31 VSSD.t365 VSSD.t364 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1466 a_7551_3677.t2 a_6927_3311.t6 a_7443_3311.t1 VDDD.t1893 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1467 a_4698_2899.t1 a_5015_3009.t6 a_4973_3133.t0 VSSD.t562 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1468 VSSD.t644 CLK.t4 a_6813_7093.t5 VSSD.t643 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1469 VSSD.t1072 a_7948_7637.t13 clkload0.X.t13 VSSD.t1071 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1470 a_5055_3285.t1 a_5342_3563.t5 VDDD.t199 VDDD.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1471 VSSD.t1051 a_10851_5461.t6 CF[7].t2 VSSD.t1050 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1472 a_2509_11169.t0 a_2291_10927.t4 VDDD.t204 VDDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1473 VSSD.t419 a_4619_4636.t5 a_4550_4765.t1 VSSD.t418 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1474 SWP[8].t0 a_1651_4917.t7 VDDD.t1270 VDDD.t1269 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1475 VDDD.t1323 a_10667_9599.t8 DOUT[0].t0 VDDD.t1322 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1476 a_10746_6031.t0 a_9669_6037.t5 a_10584_6409.t0 VDDD.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1477 a_2659_10761.t0 a_2143_10389.t7 a_2564_10749.t0 VSSD.t810 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1478 a_2196_10927.t1 x2/net8.t5 VSSD.t437 VSSD.t436 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1479 VSSD.t498 EN.t58 a_9821_7485.t1 VSSD.t497 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1480 a_9112_10761.t1 a_8031_10389.t4 a_8765_10357.t0 VDDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1481 a_4181_6575.t1 a_4146_6827.t5 a_3859_6549.t1 VSSD.t1635 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1482 a_7708_9117.t2 a_7494_9117.t5 VDDD.t124 VDDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1483 VDDD.t1640 a_7331_9269.t16 x3/COMP_BUF_N.t1 VDDD.t1639 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1484 a_4463_8893.t0 CF[0].t10 VDDD.t1578 VDDD.t1577 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1485 a_7723_11775.t0 EN.t59 VDDD.t1487 VDDD.t1486 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1486 VSSD.t367 x3/COMP_BUF_P.t32 a_2974_4943.t1 VSSD.t366 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1487 a_7348_5487.t0 x3/COMP_BUF_P.t33 VDDD.t450 VDDD.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1488 VDDD.t996 VSSD.t1947 VDDD.t995 VDDD.t994 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1489 a_10286_7119.t1 a_9209_7125.t5 a_10124_7497.t1 VDDD.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1490 VDDD.t1489 EN.t60 a_5040_10383.t2 VDDD.t1488 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1491 VDDD.t1447 a_4993_3829.t5 a_4883_3855.t2 VDDD.t1446 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1492 a_1941_10927.t1 a_1775_10927.t6 VSSD.t529 VSSD.t528 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1493 VSSD.t1613 x2/net6.t7 x2/net12.t3 VSSD.t1612 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1494 a_6942_6941.t2 a_6855_6717.t6 a_6538_6827.t1 VDDD.t1485 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1495 a_10035_4943.t1 CLKS.t107 VDDD.t308 VDDD.t307 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1496 a_7201_11445.t1 a_6983_11849.t5 VSSD.t320 VSSD.t319 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1497 VDDD.t716 a_7171_7637.t8 DOUT[6].t0 VDDD.t715 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1498 VDDD.t377 a_10759_6335.t7 CF[8].t2 VDDD.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1499 a_10207_8725.t0 EN.t61 VDDD.t1491 VDDD.t1490 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1500 a_8183_5461.t2 a_8008_5487.t5 a_8362_5487.t0 VSSD.t1024 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1501 a_8262_6031.t1 a_7185_6037.t5 a_8100_6409.t2 VDDD.t597 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1502 VSSD.t330 a_2779_6005.t5 a_2710_6031.t1 VSSD.t329 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1503 a_5366_8029.t0 a_4647_7805.t7 a_4803_7900.t1 VSSD.t1745 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1504 a_10478_7485.t1 EN.t62 VSSD.t1138 VSSD.t1137 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1505 a_6081_7663.t0 a_5915_7663.t6 VDDD.t113 VDDD.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1506 CLKSB.t1 CLKS.t108 VSSD.t247 VSSD.t246 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1507 a_1754_8339.t1 a_2032_8323.t4 a_1988_8207.t0 VDDD.t726 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1508 VDDD.t722 x2/net13.t18 CLKS.t3 VDDD.t721 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1509 a_2585_11477.t0 a_2419_11477.t6 VDDD.t1284 VDDD.t1283 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1510 a_7367_4765.t1 CLKS.t109 VDDD.t310 VDDD.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1511 a_4550_4765.t3 a_4424_4667.t4 a_4146_4651.t2 VSSD.t707 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1512 VDDD.t464 a_10492_5321.t5 a_10667_5247.t2 VDDD.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1513 a_3399_10687.t2 EN.t63 VDDD.t1493 VDDD.t1492 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1514 a_7185_6037.t0 a_7019_6037.t6 VDDD.t6 VDDD.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1515 a_4057_12015.t0 a_3891_12015.t4 VDDD.t99 VDDD.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1516 a_10846_9661.t1 EN.t64 VSSD.t1140 VSSD.t1139 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1517 VDDD.t999 VSSD.t1948 VDDD.t998 VDDD.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1518 VDDD.t1395 a_10851_5461.t7 a_10838_5853.t0 VDDD.t1394 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1519 a_8008_5487.t3 a_6927_5487.t6 a_7661_5729.t3 VDDD.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1520 a_1789_8573.t0 a_1754_8339.t5 a_1467_8181.t0 VSSD.t1587 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1521 a_1941_10927.t0 a_1775_10927.t7 VDDD.t690 VDDD.t689 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1522 a_2833_9839.t0 EN.t65 VSSD.t1142 VSSD.t1141 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1523 a_10785_3311.t0 a_9595_3311.t7 a_10676_3311.t2 VSSD.t1121 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1524 VSSD.t1088 x3/COMP_BUF_N.t30 a_5366_8029.t3 VSSD.t1087 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1525 VSSD.t337 x3/COMP_BUF_N.t31 a_7574_6941.t1 VSSD.t336 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1526 VSSD.t1291 VDDD.t2078 VSSD.t1290 VSSD.t1289 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1527 VDDD.t415 x3/COMP_BUF_N.t32 a_7574_6941.t0 VDDD.t414 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1528 VSSD.t1082 a_10299_7423.t8 DOUT[3].t2 VSSD.t1081 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1529 VDDD.t775 a_3859_8725.t7 SWN[0].t0 VDDD.t774 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1530 a_7723_11775.t1 a_7548_11849.t4 a_7902_11837.t1 VSSD.t1704 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1531 VDDD.t1002 VSSD.t1949 VDDD.t1001 VDDD.t1000 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1532 a_9112_10761.t2 a_8197_10389.t5 a_8765_10357.t1 VSSD.t132 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1533 a_7948_7637.t3 clknet_1_0__leaf_CLK.t48 VSSD.t429 VSSD.t428 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1534 VSSD.t1288 VDDD.t2079 VSSD.t1287 VSSD.t1286 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1535 x3/COMP_BUF_P.t1 a_8435_8181.t18 VDDD.t926 VDDD.t925 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1536 VSSD.t610 a_7654_4943.t28 clknet_1_0__leaf_CLK.t22 VSSD.t609 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1537 VSSD.t1285 VDDD.t2080 VSSD.t1284 VSSD.t1283 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1538 a_9467_10927.t1 a_8951_10927.t5 a_9372_10927.t3 VSSD.t1150 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1539 a_5113_7663.t0 a_4734_8029.t5 a_5041_7663.t0 VSSD.t103 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1540 x3/COMP_BUF_N.t11 a_7331_9269.t17 VSSD.t1630 VSSD.t1629 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1541 a_10145_4917.t1 a_9927_5321.t4 VDDD.t1356 VDDD.t1355 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1542 a_2790_8207.t1 a_2071_8449.t5 a_2227_8181.t2 VSSD.t524 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1543 a_7324_9117.t0 a_6803_8725.t6 VDDD.t1566 VDDD.t1565 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1544 clknet_1_0__leaf_CLK.t11 a_7654_4943.t29 VDDD.t647 VDDD.t646 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1545 VDDD.t600 a_7753_6005.t4 a_7643_6031.t1 VDDD.t599 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1546 a_5171_11445.t2 a_5015_11713.t6 a_5316_11471.t2 VDDD.t1372 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1547 VSSD.t680 a_4895_10357.t5 a_4826_10383.t3 VSSD.t679 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1548 VSSD.t27 clknet_0_CLK.t43 a_7654_4943.t4 VSSD.t26 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1549 VSSD.t1282 VDDD.t2081 VSSD.t1281 VSSD.t1280 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1550 a_6796_8573.t3 SWP[5].t5 VSSD.t651 VSSD.t650 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1551 a_6378_3677.t2 a_5659_3453.t5 a_5815_3548.t1 VSSD.t634 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1552 VSSD.t1279 VDDD.t2082 VSSD.t1278 VSSD.t1257 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1553 VDDD.t1005 VSSD.t1950 VDDD.t1004 VDDD.t1003 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1554 VSSD.t305 a_1835_9813.t7 x2/net8.t2 VSSD.t304 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1555 a_7093_3311.t0 a_6927_3311.t7 VDDD.t1895 VDDD.t1894 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1556 VSSD.t454 a_8459_4159.t6 a_8393_4233.t0 VSSD.t453 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1557 VSSD.t713 CF[3].t9 a_8126_2767.t1 VSSD.t712 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1558 a_4625_12257.t3 a_4407_12015.t5 VSSD.t1611 VSSD.t1610 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1559 a_10846_9839.t1 EN.t66 VSSD.t1588 VSSD.t1139 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1560 a_3399_10687.t1 a_3224_10761.t5 a_3578_10749.t0 VSSD.t69 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1561 VDDD.t838 a_9287_10687.t7 x2/net5.t1 VDDD.t837 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1562 VDDD.t1008 VSSD.t1951 VDDD.t1007 VDDD.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1563 a_5659_3453.t0 clknet_1_0__leaf_CLK.t49 VDDD.t580 VDDD.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1564 a_4457_10749.t1 a_4422_10515.t5 a_4135_10357.t1 VSSD.t868 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1565 VSSD.t1844 a_2019_6005.t8 SWN[8].t2 VSSD.t1843 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1566 VDDD.t1011 VSSD.t1952 VDDD.t1010 VDDD.t1009 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1567 VDDD.t872 a_10207_8725.t7 a_10194_9117.t1 VDDD.t871 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1568 x2/net6.t0 a_3399_10687.t8 VDDD.t176 VDDD.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1569 VSSD.t17 a_10759_4159.t7 CF[5].t3 VSSD.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1570 VSSD.t955 CF[2].t8 a_6378_3677.t1 VSSD.t954 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1571 VDDD.t1014 VSSD.t1953 VDDD.t1013 VDDD.t1012 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1572 a_10492_5321.t0 a_9411_4949.t7 a_10145_4917.t0 VDDD.t1459 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1573 VDDD.t1017 VSSD.t1954 VDDD.t1016 VDDD.t1015 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1574 VSSD.t785 clknet_1_1__leaf_CLK.t43 a_6927_10927.t1 VSSD.t784 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1575 VSSD.t1277 VDDD.t2083 VSSD.t1276 VSSD.t1275 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1576 VSSD.t1074 a_7948_7637.t14 clkload0.X.t12 VSSD.t1073 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1577 SWN[1].t0 a_6251_6549.t8 VDDD.t739 VDDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1578 clkload0.X.t0 a_7948_7637.t15 VDDD.t1410 VDDD.t1409 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1579 CF[1].t0 a_5055_3285.t8 VDDD.t1 VDDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1580 VDDD.t1020 VSSD.t1955 VDDD.t1019 VDDD.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1581 a_9927_9673.t1 a_9411_9301.t5 a_9832_9661.t1 VSSD.t1023 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1582 a_1988_9117.t1 a_1467_8725.t7 VDDD.t420 VDDD.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1583 a_10035_9295.t0 a_9411_9301.t6 a_9927_9673.t0 VDDD.t1361 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1584 a_6125_3311.t0 a_5746_3677.t5 a_6053_3311.t1 VSSD.t770 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1585 VDDD.t1337 a_4411_11445.t7 x2/net1.t1 VDDD.t1336 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1586 a_8435_8181.t0 COMP_P.t4 VDDD.t422 VDDD.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1587 a_4407_12015.t1 a_4057_12015.t4 a_4312_12015.t1 VDDD.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1588 VSSD.t787 clknet_1_1__leaf_CLK.t44 a_8031_10389.t1 VSSD.t786 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1589 SWP[7].t0 a_1835_4373.t8 VDDD.t390 VDDD.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1590 a_10127_6031.t1 a_9503_6037.t4 a_10019_6409.t2 VDDD.t915 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1591 VSSD.t1274 VDDD.t2084 VSSD.t1273 VSSD.t1272 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1592 VSSD.t1271 VDDD.t2085 VSSD.t1270 VSSD.t1269 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1593 a_4057_12015.t1 a_3891_12015.t5 VSSD.t73 VSSD.t72 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1594 VDDD.t1023 VSSD.t1956 VDDD.t1022 VDDD.t1021 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1595 VSSD.t1268 VDDD.t2086 VSSD.t1267 VSSD.t1266 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1596 VDDD.t649 a_7654_4943.t30 clknet_1_0__leaf_CLK.t12 VDDD.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1597 a_9924_4221.t2 CF[6].t8 VSSD.t1624 VSSD.t1623 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1598 VSSD.t1265 VDDD.t2087 VSSD.t1264 VSSD.t1263 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1599 a_5607_10927.t1 a_5161_10927.t3 a_5511_10927.t1 VSSD.t66 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1600 VSSD.t900 a_4135_10357.t8 x2/net7.t2 VSSD.t899 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1601 VDDD.t1026 VSSD.t1957 VDDD.t1025 VDDD.t1024 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1602 VDDD.t1029 VSSD.t1958 VDDD.t1028 VDDD.t1027 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1603 x2/net13.t2 x2/net12.t10 VSSD.t647 VSSD.t646 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1604 VSSD.t757 a_8435_8181.t19 x3/COMP_BUF_P.t9 VSSD.t756 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1605 VSSD.t249 CLKS.t110 a_10281_3133.t0 VSSD.t248 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1606 VSSD.t389 CF[0].t11 a_7019_6037.t1 VSSD.t388 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1607 VDDD.t760 clknet_1_1__leaf_CLK.t45 a_6927_10927.t0 VDDD.t759 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1608 a_9669_3861.t1 a_9503_3861.t6 VSSD.t1579 VSSD.t1578 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1609 VDDD.t1032 VSSD.t1959 VDDD.t1031 VDDD.t1030 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1610 VDDD.t1035 VSSD.t1960 VDDD.t1034 VDDD.t1033 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1611 a_4929_6575.t1 a_4550_6941.t5 a_4857_6575.t1 VSSD.t1699 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1612 VDDD.t1964 CKO.t16 a_8951_8751.t0 VDDD.t1963 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1613 clknet_0_CLK.t4 a_6813_7093.t31 VDDD.t1503 VDDD.t1502 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1614 VSSD.t1837 CKO.t17 a_8951_7663.t1 VSSD.t1836 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1615 VSSD.t1590 EN.t67 a_9729_8751.t0 VSSD.t1589 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1616 VDDD.t626 a_7999_4373.t6 a_7986_4765.t0 VDDD.t625 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1617 VSSD.t599 clknet_1_1__leaf_CLK.t46 a_1775_10927.t1 VSSD.t598 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1618 VDDD.t82 a_5815_3548.t4 a_5746_3677.t1 VDDD.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1619 VDDD.t1281 a_6803_2741.t7 CF[2].t2 VDDD.t1280 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1620 a_10141_8751.t1 a_8951_8751.t7 a_10032_8751.t2 VSSD.t1021 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1621 clknet_0_CLK.t19 a_6813_7093.t32 VSSD.t1148 VSSD.t1147 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1622 a_7158_8029.t0 a_6081_7663.t5 a_6996_7663.t2 VDDD.t411 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1623 VDDD.t254 CLKS.t111 a_6803_8725.t2 VDDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1624 a_10032_7663.t0 a_9117_7663.t4 a_9685_7905.t0 VSSD.t432 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1625 a_10219_5853.t1 CLKS.t112 VDDD.t256 VDDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1626 VDDD.t566 a_10207_10901.t6 x2/net11.t0 VDDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1627 VSSD.t1262 VDDD.t2088 VSSD.t1261 VSSD.t1260 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1628 VSSD.t210 CLKS.t113 a_2157_5487.t0 VSSD.t209 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1629 a_5040_10383.t0 a_4826_10383.t5 VDDD.t849 VDDD.t848 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1630 clknet_0_CLK.t3 a_6813_7093.t33 VDDD.t1505 VDDD.t1504 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1631 a_9467_7663.t0 a_9117_7663.t5 a_9372_7663.t0 VDDD.t583 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1632 a_5015_11713.t1 clknet_1_1__leaf_CLK.t47 VSSD.t601 VSSD.t600 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1633 a_10237_6005.t3 a_10019_6409.t4 VSSD.t1809 VSSD.t1808 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1634 a_10386_8751.t0 EN.t68 VSSD.t1592 VSSD.t1591 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1635 VSSD.t926 a_8183_5461.t7 SWP[1].t2 VSSD.t925 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1636 CLKS.t4 x2/net13.t19 VDDD.t724 VDDD.t723 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1637 a_5481_3133.t0 a_5102_2767.t4 a_5409_3133.t0 VSSD.t34 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1638 a_5182_4765.t2 a_4463_4541.t6 a_4619_4636.t3 VSSD.t834 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1639 VSSD.t1259 VDDD.t2089 VSSD.t1258 VSSD.t1257 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1640 VSSD.t212 CLKS.t114 a_5101_5487.t1 VSSD.t211 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1641 a_7535_6409.t0 a_7019_6037.t7 a_7440_6397.t2 VSSD.t3 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1642 VDDD.t762 clknet_1_1__leaf_CLK.t48 a_1775_10927.t0 VDDD.t761 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1643 VDDD.t1111 VSSD.t1961 VDDD.t1110 VDDD.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1644 a_6999_8207.t0 a_6375_8213.t7 a_6891_8585.t1 VDDD.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1645 VDDD.t614 a_8459_4159.t7 a_8446_3855.t0 VDDD.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1646 VSSD.t539 a_4411_2741.t8 SWP[4].t2 VSSD.t538 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1647 VDDD.t193 a_5307_7093.t16 FINAL.t2 VDDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1648 a_6813_7093.t4 CLK.t5 VSSD.t361 VSSD.t360 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1649 VDDD.t1114 VSSD.t1962 VDDD.t1113 VDDD.t1112 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1650 clkload0.X.t11 a_7948_7637.t16 VSSD.t1076 VSSD.t1075 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1651 a_10145_9269.t2 a_9927_9673.t4 VSSD.t854 VSSD.t853 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1652 a_2439_9981.t1 clknet_1_1__leaf_CLK.t49 VSSD.t603 VSSD.t602 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1653 VDDD.t1117 VSSD.t1963 VDDD.t1116 VDDD.t1115 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1654 x2/net12.t2 x2/net6.t8 VSSD.t865 VSSD.t864 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1655 a_9575_8029.t1 a_8951_7663.t6 a_9467_7663.t3 VDDD.t1230 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1656 VDDD.t1582 EN.t69 a_4411_11445.t2 VDDD.t1581 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1657 a_5849_5487.t0 a_5470_5853.t4 a_5777_5487.t0 VSSD.t1692 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1658 a_10851_5461.t0 CLKS.t115 VDDD.t258 VDDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1659 a_6693_7663.t0 a_6649_7905.t4 a_6527_7663.t0 VSSD.t760 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1660 a_10386_10927.t1 EN.t70 VSSD.t1594 VSSD.t1593 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1661 VSSD.t1256 VDDD.t2090 VSSD.t1255 VSSD.t1254 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1662 VSSD.t1595 EN.t71 a_1789_8573.t1 VSSD.t478 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1663 VSSD.t1253 VDDD.t2091 VSSD.t1252 VSSD.t1251 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1664 VDDD.t1966 CKO.t18 a_5915_7663.t0 VDDD.t1965 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1665 VDDD.t930 a_6649_7905.t5 a_6539_8029.t1 VDDD.t929 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1666 a_1988_8207.t1 a_1467_8181.t7 VDDD.t446 VDDD.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1667 VSSD.t1250 VDDD.t2092 VSSD.t1249 VSSD.t1248 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1668 a_10693_6409.t0 a_9503_6037.t5 a_10584_6409.t2 VSSD.t747 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1669 a_2071_8449.t1 CKO.t19 VSSD.t1838 VSSD.t1160 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1670 VSSD.t640 a_10207_10901.t7 a_10141_10927.t1 VSSD.t639 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1671 SWP[9].t0 a_4779_5461.t6 VDDD.t538 VDDD.t537 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1672 a_4564_8029.t0 a_4043_7637.t7 VDDD.t1887 VDDD.t1886 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1673 VSSD.t1152 a_2595_5724.t5 a_2526_5853.t1 VSSD.t1151 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1674 VSSD.t152 a_5307_7093.t17 FINAL.t10 VSSD.t151 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1675 VDDD.t1628 a_2439_4541.t6 a_2400_4667.t0 VDDD.t1627 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1676 a_10654_10205.t0 a_9577_9839.t5 a_10492_9839.t3 VDDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1677 VDDD.t1220 a_1835_9813.t8 x2/net8.t0 VDDD.t1219 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1678 a_8183_10901.t2 EN.t72 VDDD.t1584 VDDD.t1583 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1679 VDDD.t1120 VSSD.t1964 VDDD.t1119 VDDD.t1118 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1680 a_4647_7805.t1 CF[4].t8 VSSD.t630 VSSD.t629 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1681 a_8425_6603.t1 FINAL.t19 a_8339_6603.t1 VSSD.t458 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1682 VSSD.t1247 VDDD.t2093 VSSD.t1246 VSSD.t1245 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1683 VDDD.t883 a_10676_3311.t5 a_10851_3285.t2 VDDD.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1684 a_2595_5724.t0 a_2439_5629.t7 a_2740_5853.t1 VDDD.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1685 a_9924_6397.t0 CF[9].t9 VDDD.t958 VDDD.t957 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1686 VDDD.t1252 EN.t73 a_2372_9117.t2 VDDD.t1251 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1687 VSSD.t339 x3/COMP_BUF_N.t33 a_5090_8207.t3 VSSD.t338 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1688 a_10194_11293.t1 a_9117_10927.t4 a_10032_10927.t3 VDDD.t1368 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1689 VSSD.t1244 VDDD.t2094 VSSD.t1243 VSSD.t1242 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1690 a_2595_4636.t0 a_2400_4667.t5 a_2905_4399.t1 VSSD.t226 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1691 a_4857_4399.t0 CLKS.t116 VSSD.t214 VSSD.t213 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1692 a_9464_7485.t2 SWP[3].t5 VDDD.t155 VDDD.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1693 a_7705_3311.t0 a_7661_3553.t5 a_7539_3311.t0 VSSD.t953 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1694 a_7661_5729.t2 a_7443_5487.t5 VSSD.t1739 VSSD.t1738 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1695 a_8170_5853.t0 a_7093_5487.t4 a_8008_5487.t1 VDDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1696 a_2595_10076.t3 a_2439_9981.t6 a_2740_10205.t0 VDDD.t1622 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1697 a_2157_9839.t0 a_2122_10091.t5 a_1835_9813.t0 VSSD.t1018 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1698 a_10746_2767.t1 a_9669_2773.t5 a_10584_3145.t1 VDDD.t779 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1699 VDDD.t1390 a_4463_6717.t6 a_4424_6843.t0 VDDD.t1389 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1700 a_4739_10625.t0 clknet_1_1__leaf_CLK.t50 VDDD.t530 VDDD.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1701 a_10584_4233.t2 a_9669_3861.t3 a_10237_3829.t3 VSSD.t1806 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1702 a_2526_5853.t3 a_2400_5755.t4 a_2122_5739.t3 VSSD.t744 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1703 a_8765_10357.t3 a_8547_10761.t5 VSSD.t989 VSSD.t988 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1704 a_4054_8339.t3 a_4332_8323.t5 a_4288_8207.t1 VDDD.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1705 VDDD.t1348 clknet_1_0__leaf_CLK.t50 a_6927_3311.t0 VDDD.t1347 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1706 VDDD.t651 a_7654_4943.t31 clknet_1_0__leaf_CLK.t13 VDDD.t650 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1707 a_2122_4651.t3 a_2439_4541.t7 a_2397_4399.t1 VSSD.t1614 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1708 VSSD.t1098 a_5171_11445.t5 a_5102_11471.t3 VSSD.t1097 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1709 x2/net11.t2 a_10207_10901.t8 VSSD.t642 VSSD.t641 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1710 x3/COMP_BUF_N.t10 a_7331_9269.t18 VSSD.t1632 VSSD.t1631 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1711 a_3158_5853.t1 a_2400_5755.t5 a_2595_5724.t3 VDDD.t909 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1712 VSSD.t1001 clknet_1_0__leaf_CLK.t51 a_7948_7637.t2 VSSD.t1000 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1713 SWP[2].t2 a_7999_4373.t7 VSSD.t460 VSSD.t459 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1714 a_2755_10761.t1 a_2309_10389.t3 a_2659_10761.t2 VSSD.t1752 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1715 a_7331_9269.t0 COMP_N.t5 VDDD.t212 VDDD.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1716 a_7407_3009.t1 clknet_1_0__leaf_CLK.t52 VSSD.t1003 VSSD.t1002 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1717 clknet_1_0__leaf_CLK.t14 a_7654_4943.t32 VSSD.t485 VSSD.t484 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1718 VSSD.t1241 VDDD.t2095 VSSD.t1240 VSSD.t1239 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1719 VDDD.t1380 a_10759_3071.t7 CF[3].t1 VDDD.t1379 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1720 VDDD.t1123 VSSD.t1965 VDDD.t1122 VDDD.t1121 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1721 VSSD.t1238 VDDD.t2096 VSSD.t1237 VSSD.t1222 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1722 VDDD.t1126 VSSD.t1966 VDDD.t1125 VDDD.t1124 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1723 VSSD.t440 a_10943_6549.t8 a_10877_6575.t1 VSSD.t439 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1724 VSSD.t391 CF[0].t12 a_5307_7093.t4 VSSD.t390 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1725 a_7661_11169.t1 a_7443_10927.t5 VSSD.t196 VSSD.t195 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1726 a_7539_10927.t1 a_7093_10927.t4 a_7443_10927.t3 VSSD.t730 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1727 a_10465_6575.t1 a_10421_6817.t5 a_10299_6575.t1 VSSD.t474 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1728 VSSD.t1236 VDDD.t2097 VSSD.t1235 VSSD.t1234 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1729 a_4895_10357.t2 a_4700_10499.t5 a_5205_10749.t1 VSSD.t1030 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1730 a_10329_3553.t1 a_10111_3311.t4 VDDD.t750 VDDD.t749 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1731 VDDD.t1311 a_10207_7637.t7 DOUT[4].t0 VDDD.t1310 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1732 VDDD.t970 a_7723_11775.t7 x2/net3.t0 VDDD.t969 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1733 VDDD.t1129 VSSD.t1967 VDDD.t1128 VDDD.t1127 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1734 a_6102_5853.t3 a_5344_5755.t5 a_5539_5724.t2 VDDD.t746 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1735 DOUT[2].t0 a_10207_8725.t8 VDDD.t874 VDDD.t873 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1736 VDDD.t260 CLKS.t117 a_4043_7637.t0 VDDD.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1737 VSSD.t29 clknet_0_CLK.t44 a_6077_9813.t3 VSSD.t28 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1738 a_2071_8893.t0 CKO.t20 VDDD.t1968 VDDD.t1967 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1739 VDDD.t1132 VSSD.t1968 VDDD.t1131 VDDD.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1740 a_8197_10389.t0 a_8031_10389.t5 VDDD.t141 VDDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1741 VDDD.t1889 a_4043_7637.t8 SWN[4].t0 VDDD.t1888 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1742 a_7797_6397.t1 a_7753_6005.t5 a_7631_6409.t0 VSSD.t442 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1743 VSSD.t216 CLKS.t118 a_7125_8751.t1 VSSD.t215 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1744 VDDD.t683 a_2071_8449.t6 a_2032_8323.t1 VDDD.t682 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1745 VDDD.t787 a_7661_5729.t5 a_7551_5853.t2 VDDD.t786 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1746 a_10108_6575.t3 EN.t74 VSSD.t916 VSSD.t915 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1747 VDDD.t532 clknet_1_1__leaf_CLK.t51 a_2143_10389.t0 VDDD.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1748 a_10654_4943.t1 a_9577_4949.t5 a_10492_5321.t2 VDDD.t612 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1749 VSSD.t174 x2/TRIG1.t5 a_5734_11471.t3 VSSD.t173 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1750 VDDD.t1135 VSSD.t1969 VDDD.t1134 VDDD.t1133 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1751 VSSD.t1233 VDDD.t2098 VSSD.t1232 VSSD.t1231 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1752 x3/COMP_BUF_P.t0 a_8435_8181.t20 VDDD.t928 VDDD.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1753 a_5081_12015.t0 a_3891_12015.t6 a_4972_12015.t0 VSSD.t74 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1754 a_3153_11445.t3 a_2935_11849.t5 VSSD.t946 VSSD.t945 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1755 CF[2].t3 a_6803_2741.t8 VSSD.t1748 VSSD.t1747 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1756 VDDD.t1137 VSSD.t1970 VDDD.t1136 VDDD.t1030 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1757 clkload0.X.t10 a_7948_7637.t17 VSSD.t593 VSSD.t592 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1758 VSSD.t1230 VDDD.t2099 VSSD.t1229 VSSD.t1228 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1759 a_2509_11169.t1 a_2291_10927.t5 VSSD.t158 VSSD.t157 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1760 a_9761_5487.t0 a_9595_5487.t6 VDDD.t1914 VDDD.t1913 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1761 VDDD.t1254 EN.t75 a_2372_8207.t2 VDDD.t1253 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1762 a_7986_4765.t1 a_6909_4399.t5 a_7824_4399.t1 VDDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1763 VDDD.t1140 VSSD.t1971 VDDD.t1139 VDDD.t1138 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1764 VDDD.t208 a_5383_5629.t7 a_5344_5755.t0 VDDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1765 VDDD.t1675 CLKS.t119 a_4948_8029.t1 VDDD.t1674 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1766 VDDD.t1248 clknet_0_CLK.t45 a_6077_9813.t5 VDDD.t1247 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1767 VSSD.t1733 a_5515_4159.t8 SWP[5].t2 VSSD.t1732 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1768 VSSD.t176 a_5171_2741.t5 a_5102_2767.t2 VSSD.t175 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1769 clknet_1_0__leaf_CLK.t15 a_7654_4943.t33 VDDD.t653 VDDD.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1770 a_5316_6031.t1 a_5102_6031.t5 VDDD.t934 VDDD.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1771 a_2122_7915.t2 a_2400_7931.t5 a_2356_8029.t1 VDDD.t1534 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1772 VSSD.t759 a_8435_8181.t21 x3/COMP_BUF_P.t8 VSSD.t758 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1773 VDDD.t951 a_8765_10357.t5 a_8655_10383.t0 VDDD.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1774 VSSD.t701 a_4619_8988.t5 a_4550_9117.t2 VSSD.t700 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1775 a_9563_10927.t0 a_9117_10927.t5 a_9467_10927.t3 VSSD.t1029 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1776 a_10035_9295.t2 EN.t76 VDDD.t1256 VDDD.t1255 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1777 VDDD.t1507 a_6813_7093.t34 clknet_0_CLK.t2 VDDD.t1506 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1778 a_7440_6397.t1 x3/COMP_BUF_P.t34 VSSD.t858 VSSD.t857 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1779 VSSD.t1049 a_4463_6717.t7 a_4424_6843.t1 VSSD.t1048 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1780 VDDD.t1143 VSSD.t1972 VDDD.t1142 VDDD.t1141 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1781 VDDD.t1315 a_6813_7093.t35 clknet_0_CLK.t1 VDDD.t1314 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1782 a_2556_4943.t0 a_2342_4943.t5 VDDD.t429 VDDD.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1783 VDDD.t1146 VSSD.t1973 VDDD.t1145 VDDD.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1784 VSSD.t974 a_6813_7093.t36 clknet_0_CLK.t18 VSSD.t973 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1785 a_8008_5487.t0 a_7093_5487.t5 a_7661_5729.t0 VSSD.t68 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1786 a_3031_10901.t1 a_2856_10927.t5 a_3210_10927.t0 VSSD.t762 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1787 VSSD.t564 a_5015_3009.t7 a_4976_2883.t1 VSSD.t563 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1788 VDDD.t586 a_10492_9673.t5 a_10667_9599.t1 VDDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1789 a_2767_10383.t2 EN.t77 VDDD.t1258 VDDD.t1257 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1790 a_7719_4233.t2 a_7203_3861.t6 a_7624_4221.t3 VSSD.t300 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1791 a_10016_5487.t2 CF[8].t8 VSSD.t1641 VSSD.t1640 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1792 VDDD.t1350 a_10584_6409.t5 a_10759_6335.t2 VDDD.t1349 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1793 a_2905_7663.t0 a_2526_8029.t5 a_2833_7663.t0 VSSD.t121 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1794 a_2585_11477.t1 a_2419_11477.t7 VSSD.t944 VSSD.t943 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1795 VSSD.t1227 VDDD.t2100 VSSD.t1226 VSSD.t1225 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1796 a_2397_7663.t0 a_1835_7637.t7 VSSD.t591 VSSD.t590 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1797 VSSD.t1224 VDDD.t2101 VSSD.t1223 VSSD.t1222 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1798 a_4550_9117.t0 a_4424_9019.t4 a_4146_9003.t0 VSSD.t548 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1799 VDDD.t370 a_2227_8988.t4 a_2158_9117.t2 VDDD.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1800 a_9117_10927.t1 a_8951_10927.t6 VSSD.t1113 VSSD.t1112 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1801 a_5729_11169.t2 a_5511_10927.t5 VDDD.t527 VDDD.t526 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1802 a_10127_2767.t2 a_9503_2773.t6 a_10019_3145.t0 VDDD.t1890 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1803 a_3870_5075.t2 a_4148_5059.t5 a_4104_4943.t1 VDDD.t1211 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1804 VSSD.t1221 VDDD.t2102 VSSD.t1220 VSSD.t1219 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1805 a_2255_5185.t0 CF[8].t9 VDDD.t1647 VDDD.t1646 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1806 VDDD.t195 a_5307_7093.t18 FINAL.t1 VDDD.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1807 a_4619_8988.t2 a_4463_8893.t6 a_4764_9117.t2 VDDD.t1553 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1808 a_4463_4541.t1 CF[6].t9 VSSD.t1626 VSSD.t1625 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1809 a_1938_5075.t1 a_2255_5185.t7 a_2213_5309.t0 VSSD.t1751 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1810 VDDD.t1275 a_4739_10625.t6 a_4700_10499.t0 VDDD.t1274 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1811 VDDD.t616 a_8459_4159.t8 SWP[3].t0 VDDD.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1812 a_4698_6163.t0 a_4976_6147.t3 a_4932_6031.t0 VDDD.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1813 a_9685_8993.t3 a_9467_8751.t5 VSSD.t1849 VSSD.t1848 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1814 VDDD.t1149 VSSD.t1974 VDDD.t1148 VDDD.t1147 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1815 VSSD.t918 EN.t78 a_10189_9661.t1 VSSD.t917 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1816 a_10943_6549.t0 CLKS.t120 VDDD.t1677 VDDD.t1676 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1817 a_10145_9269.t3 a_9927_9673.t5 VDDD.t1202 VDDD.t1201 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1818 a_5161_10927.t1 a_4995_10927.t6 VSSD.t1847 VSSD.t1846 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1819 a_6238_11293.t1 a_5161_10927.t4 a_6076_10927.t0 VDDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1820 clknet_0_CLK.t17 a_6813_7093.t37 VSSD.t976 VSSD.t975 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1821 a_2740_4765.t0 a_2526_4765.t5 VDDD.t568 VDDD.t567 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1822 a_9575_8029.t2 EN.t79 VDDD.t1260 VDDD.t1259 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1823 a_10115_4233.t1 a_9669_3861.t4 a_10019_4233.t3 VSSD.t1807 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1824 a_9117_10927.t0 a_8951_10927.t7 VDDD.t1455 VDDD.t1454 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1825 VDDD.t781 CKO.t21 a_9043_7125.t0 VDDD.t780 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1826 a_5182_9117.t0 a_4424_9019.t5 a_4619_8988.t1 VDDD.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1827 VDDD.t1892 a_8008_3311.t5 a_8183_3285.t2 VDDD.t895 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1828 VDDD.t1325 a_4619_6812.t5 a_4550_6941.t2 VDDD.t1324 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1829 VDDD.t1679 CLKS.t121 a_8615_7457.t0 VDDD.t1678 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1830 VSSD.t1005 clknet_1_0__leaf_CLK.t53 a_9411_4949.t1 VSSD.t1004 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1831 VSSD.t375 a_6077_9813.t32 clknet_1_1__leaf_CLK.t17 VSSD.t374 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1832 a_2172_4943.t0 a_1651_4917.t8 VDDD.t74 VDDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1833 a_10237_6005.t2 a_10019_6409.t5 VDDD.t1420 VDDD.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1834 VSSD.t1218 VDDD.t2103 VSSD.t1217 VSSD.t1216 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1835 VDDD.t628 a_7999_4373.t8 SWP[2].t0 VDDD.t627 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1836 CF[8].t3 a_10759_6335.t8 VDDD.t379 VDDD.t378 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1837 CLKS.t12 x2/net13.t20 VDDD.t1404 VDDD.t1403 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1838 a_5815_3548.t0 a_5659_3453.t6 a_5960_3677.t1 VDDD.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1839 VDDD.t1692 a_7407_8893.t6 a_7368_9019.t1 VDDD.t1691 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1840 VDDD.t783 CKO.t22 a_9411_9301.t0 VDDD.t782 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1841 a_10492_9673.t0 a_9411_9301.t7 a_10145_9269.t0 VDDD.t1362 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1842 a_9777_7093.t0 a_9559_7497.t4 VDDD.t1246 VDDD.t1245 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1843 VDDD.t1236 a_8275_6335.t8 SWP[0].t0 VDDD.t1235 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1844 a_7902_11837.t0 EN.t80 VSSD.t1779 VSSD.t1778 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1845 VDDD.t1152 VSSD.t1975 VDDD.t1151 VDDD.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1846 a_5161_10927.t0 a_4995_10927.t7 VDDD.t1974 VDDD.t1973 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1847 VSSD.t487 a_7654_4943.t34 clknet_1_0__leaf_CLK.t16 VSSD.t486 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1848 a_7631_8511.t2 EN.t81 VDDD.t1900 VDDD.t1899 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1849 a_4871_4233.t1 a_4425_3861.t5 a_4775_4233.t3 VSSD.t872 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1850 a_4371_8449.t0 CF[5].t9 VSSD.t21 VSSD.t20 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1851 VSSD.t1683 CLKS.t122 a_4365_7663.t0 VSSD.t1682 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1852 VSSD.t1215 VDDD.t2104 VSSD.t1214 VSSD.t1213 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1853 VSSD.t1780 EN.t82 a_10189_9839.t1 VSSD.t917 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1854 a_6649_7905.t2 a_6431_7663.t5 VDDD.t80 VDDD.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1855 a_6983_11849.t1 a_6633_11477.t5 a_6888_11837.t0 VDDD.t1367 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1856 a_10838_5853.t1 a_9761_5487.t5 a_10676_5487.t0 VDDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1857 VSSD.t867 x2/net6.t9 a_5458_10383.t1 VSSD.t866 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1858 a_3583_4917.t2 a_3870_5075.t5 VDDD.t1514 VDDD.t1513 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1859 VSSD.t806 a_7723_11775.t8 a_7657_11849.t0 VSSD.t805 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1860 a_2227_8988.t2 a_2071_8893.t7 a_2372_9117.t0 VDDD.t847 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1861 VDDD.t1681 CLKS.t123 a_2740_5853.t0 VDDD.t1680 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1862 a_10584_6409.t3 a_9503_6037.t6 a_10237_6005.t1 VDDD.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1863 a_5307_7093.t3 CF[0].t13 VSSD.t393 VSSD.t392 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1864 a_6378_3677.t3 a_5620_3579.t4 a_5815_3548.t3 VDDD.t1512 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1865 VSSD.t1212 VDDD.t2105 VSSD.t1211 VSSD.t1210 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1866 x3/COMP_BUF_N.t9 a_7331_9269.t19 VSSD.t1634 VSSD.t1633 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1867 VDDD.t458 a_6077_9813.t33 clknet_1_1__leaf_CLK.t5 VDDD.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1868 a_7719_4233.t1 a_7369_3861.t4 a_7624_4221.t2 VDDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1869 VDDD.t460 a_6077_9813.t34 clknet_1_1__leaf_CLK.t4 VDDD.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1870 x2/TRIG1.t0 a_5147_11989.t8 VDDD.t712 VDDD.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1871 clknet_1_0__leaf_CLK.t0 a_7654_4943.t35 VDDD.t347 VDDD.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1872 a_2833_5487.t0 CLKS.t124 VSSD.t1685 VSSD.t1684 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1873 a_10124_7497.t3 a_9043_7125.t7 a_9777_7093.t2 VDDD.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1874 a_3578_10749.t1 EN.t83 VSSD.t1782 VSSD.t1781 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1875 a_10203_6575.t3 a_9687_6575.t4 a_10108_6575.t1 VSSD.t684 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1876 a_10768_6575.t1 a_9687_6575.t5 a_10421_6817.t0 VDDD.t853 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1877 VDDD.t1155 VSSD.t1976 VDDD.t1154 VDDD.t1153 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1878 a_5102_11471.t0 a_4976_11587.t4 a_4698_11603.t0 VSSD.t64 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1879 VDDD.t855 CLK.t6 a_6813_7093.t1 VDDD.t854 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1880 a_4581_5309.t0 CLKS.t125 VSSD.t1687 VSSD.t1686 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1881 a_2659_10761.t3 a_2309_10389.t4 a_2564_10749.t1 VDDD.t960 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1882 VSSD.t1209 VDDD.t2106 VSSD.t1208 VSSD.t1207 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1883 SWN[3].t0 a_6803_8725.t7 VDDD.t1568 VDDD.t1567 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1884 VSSD.t1206 VDDD.t2107 VSSD.t1205 VSSD.t1204 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1885 x2/net1.t0 a_4411_11445.t8 VDDD.t936 VDDD.t935 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1886 a_7548_11849.t1 a_6467_11477.t6 a_7201_11445.t3 VDDD.t676 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1887 a_2877_10357.t0 a_2659_10761.t5 VSSD.t97 VSSD.t96 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1888 a_2790_9117.t0 a_2032_9019.t4 a_2227_8988.t1 VDDD.t877 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1889 clknet_1_1__leaf_CLK.t3 a_6077_9813.t35 VDDD.t462 VDDD.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1890 a_9924_3133.t0 CF[4].t9 VDDD.t802 VDDD.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1891 a_8117_5487.t0 a_6927_5487.t7 a_8008_5487.t2 VSSD.t113 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1892 a_9467_7663.t2 a_8951_7663.t7 a_9372_7663.t1 VSSD.t882 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1893 a_7090_9003.t3 a_7407_8893.t7 a_7365_8751.t1 VSSD.t1696 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1894 a_9669_6037.t0 a_9503_6037.t7 VDDD.t918 VDDD.t917 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1895 a_4826_10383.t0 a_4739_10625.t7 a_4422_10515.t0 VDDD.t1273 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1896 a_7827_3855.t0 a_7203_3861.t7 a_7719_4233.t3 VDDD.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1897 VSSD.t1203 VDDD.t2108 VSSD.t1202 VSSD.t1201 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1898 VDDD.t109 a_5659_3453.t7 a_5620_3579.t0 VDDD.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1899 a_9853_6575.t0 a_9687_6575.t6 VDDD.t743 VDDD.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1900 a_8655_10383.t1 a_8031_10389.t6 a_8547_10761.t0 VDDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1901 VSSD.t1689 CLKS.t126 a_5377_3311.t0 VSSD.t1688 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1902 a_6077_9813.t6 clknet_0_CLK.t46 VSSD.t906 VSSD.t905 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1903 a_10281_4221.t0 a_10237_3829.t5 a_10115_4233.t0 VSSD.t51 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1904 VSSD.t46 a_1835_5461.t7 SWN[7].t2 VSSD.t45 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1905 VDDD.t444 a_10851_3285.t8 CF[4].t1 VDDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1906 VDDD.t1659 CLKS.t127 a_1651_4917.t0 VDDD.t1658 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1907 VSSD.t1065 x2/net13.t21 CLKS.t13 VSSD.t1064 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1908 VDDD.t417 x3/COMP_BUF_N.t34 a_5090_8207.t2 VDDD.t416 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1909 x2/net5.t2 a_9287_10687.t8 VSSD.t674 VSSD.t673 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1910 VDDD.t785 CKO.t23 a_9411_9839.t0 VDDD.t784 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1911 VDDD.t1158 VSSD.t1977 VDDD.t1157 VDDD.t1156 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1912 a_8117_10927.t0 a_6927_10927.t6 a_8008_10927.t2 VSSD.t1096 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1913 CF[5].t2 a_10759_4159.t8 VSSD.t19 VSSD.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1914 a_5171_6005.t1 a_4976_6147.t4 a_5481_6397.t1 VSSD.t301 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1915 a_8284_4233.t0 a_7369_3861.t5 a_7937_3829.t0 VSSD.t102 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1916 VDDD.t1703 a_7548_11849.t5 a_7723_11775.t2 VDDD.t1702 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1917 a_10938_4221.t0 CLKS.t128 VSSD.t1649 VSSD.t1648 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1918 a_5684_5853.t0 a_5470_5853.t5 VDDD.t1685 VDDD.t1684 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1919 VDDD.t544 a_7631_8511.t8 a_7618_8207.t1 VDDD.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1920 a_2526_8029.t0 a_2439_7805.t6 a_2122_7915.t0 VDDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1921 VDDD.t1161 VSSD.t1978 VDDD.t1160 VDDD.t1159 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1922 VDDD.t1164 VSSD.t1979 VDDD.t1163 VDDD.t1162 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1923 VSSD.t595 a_7948_7637.t18 clkload0.X.t9 VSSD.t594 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1924 VDDD.t1167 VSSD.t1980 VDDD.t1166 VDDD.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1925 a_5511_10927.t0 a_5161_10927.t5 a_5416_10927.t3 VDDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1926 VSSD.t387 a_4779_5461.t7 SWP[9].t2 VSSD.t386 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1927 a_5182_9117.t3 a_4463_8893.t7 a_4619_8988.t3 VSSD.t1571 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1928 VSSD.t1784 EN.t84 a_2553_10927.t1 VSSD.t1783 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1929 VSSD.t1200 VDDD.t2109 VSSD.t1199 VSSD.t1198 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1930 SWP[1].t0 a_8183_5461.t8 VDDD.t202 VDDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1931 a_6813_7093.t0 CLK.t7 VDDD.t1555 VDDD.t1554 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1932 a_3767_8181.t2 a_4054_8339.t5 VDDD.t1401 VDDD.t1400 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1933 VDDD.t1170 VSSD.t1981 VDDD.t1169 VDDD.t1168 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1934 VDDD.t1898 a_4371_8449.t7 a_4332_8323.t0 VDDD.t1897 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1935 a_8362_5487.t1 CLKS.t129 VSSD.t1651 VSSD.t1650 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1936 a_4733_6397.t1 a_4698_6163.t4 a_4411_6005.t1 VSSD.t1716 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1937 a_10421_6817.t2 a_10203_6575.t5 VDDD.t1698 VDDD.t1697 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1938 VSSD.t383 clknet_1_1__leaf_CLK.t52 a_4995_10927.t1 VSSD.t382 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1939 VSSD.t1197 VDDD.t2110 VSSD.t1196 VSSD.t1195 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1940 a_2227_8181.t3 a_2071_8449.t7 a_2372_8207.t1 VDDD.t684 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1941 VSSD.t1194 VDDD.t2111 VSSD.t1193 VSSD.t1192 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1942 a_4734_8029.t3 a_4608_7931.t4 a_4330_7915.t1 VSSD.t588 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1943 clknet_0_CLK.t0 a_6813_7093.t38 VDDD.t1317 VDDD.t1316 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1944 VDDD.t1910 a_9777_7093.t5 a_9667_7119.t2 VDDD.t1909 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1945 VSSD.t79 a_2439_7805.t7 a_2400_7931.t1 VSSD.t78 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1946 a_9832_5309.t1 CF[7].t7 VDDD.t907 VDDD.t906 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1947 VSSD.t1191 VDDD.t2112 VSSD.t1190 VSSD.t1189 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1948 a_6942_6941.t3 a_6816_6843.t5 a_6538_6827.t3 VSSD.t1795 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1949 a_2595_10076.t2 a_2400_10107.t5 a_2905_9839.t0 VSSD.t1168 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1950 a_4680_4221.t1 x3/COMP_BUF_P.t35 VSSD.t860 VSSD.t859 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1951 a_10237_2741.t2 a_10019_3145.t4 VSSD.t1719 VSSD.t1718 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1952 VDDD.t1661 CLKS.t130 a_4672_8207.t0 VDDD.t1660 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1953 a_4411_11445.t1 a_4698_11603.t5 VDDD.t97 VDDD.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1954 VSSD.t377 a_6077_9813.t36 clknet_1_1__leaf_CLK.t16 VSSD.t376 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1955 a_9777_7093.t1 a_9559_7497.t5 VSSD.t904 VSSD.t903 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1956 VSSD.t63 a_5815_3548.t5 a_5746_3677.t2 VSSD.t62 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1957 VDDD.t1465 a_4187_5185.t5 a_4148_5059.t0 VDDD.t1464 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1958 VSSD.t1786 EN.t85 a_6693_7663.t1 VSSD.t1785 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1959 x2/net10.t2 a_3675_11775.t8 VSSD.t585 VSSD.t584 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1960 a_4698_11603.t3 a_5015_11713.t7 a_4973_11837.t1 VSSD.t1035 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1961 a_2356_5853.t0 a_1835_5461.t8 VDDD.t1313 VDDD.t1312 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1962 a_2122_10091.t3 a_2439_9981.t7 a_2397_9839.t1 VSSD.t1617 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1963 clknet_1_1__leaf_CLK.t2 a_6077_9813.t37 VDDD.t1598 VDDD.t1597 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1964 VDDD.t534 clknet_1_1__leaf_CLK.t53 a_4995_10927.t0 VDDD.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1965 a_8435_8181.t1 COMP_P.t5 VDDD.t424 VDDD.t423 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1966 a_2790_8207.t0 a_2032_8323.t5 a_2227_8181.t0 VDDD.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1967 clkload0.X.t8 a_7948_7637.t19 VSSD.t597 VSSD.t596 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1968 a_7090_2899.t0 a_7368_2883.t5 a_7324_2767.t0 VDDD.t1327 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1969 a_3224_10761.t2 a_2309_10389.t5 a_2877_10357.t2 VSSD.t796 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1970 CF[0].t2 a_8183_3285.t7 VSSD.t503 VSSD.t502 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1971 a_10219_5853.t2 a_9595_5487.t7 a_10111_5487.t2 VDDD.t1915 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1972 VDDD.t1707 SWP[9].t5 a_3158_8029.t3 VDDD.t1706 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1973 x2/net13.t3 x2/net12.t11 VSSD.t649 VSSD.t648 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1974 a_7933_4399.t1 a_6743_4399.t7 a_7824_4399.t3 VSSD.t445 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1975 VDDD.t851 a_6076_10927.t5 a_6251_10901.t1 VDDD.t850 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1976 a_4274_4943.t3 a_4187_5185.t6 a_3870_5075.t1 VDDD.t1466 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1977 a_4857_8751.t0 CLKS.t131 VSSD.t1653 VSSD.t1652 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1978 a_5300_5853.t1 a_4779_5461.t8 VDDD.t540 VDDD.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1979 VDDD.t1172 VSSD.t1982 VDDD.t1171 VDDD.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1980 a_10019_4233.t0 a_9503_3861.t7 a_9924_4221.t0 VSSD.t1580 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1981 a_5316_2767.t0 a_5102_2767.t5 VDDD.t44 VDDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1982 a_9853_6575.t1 a_9687_6575.t7 VSSD.t576 VSSD.t575 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1983 a_4803_7900.t3 a_4608_7931.t5 a_5113_7663.t1 VSSD.t589 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1984 a_4739_10625.t1 clknet_1_1__leaf_CLK.t54 VSSD.t385 VSSD.t384 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1985 CKO.t3 a_8339_6603.t4 VSSD.t1800 VSSD.t1799 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1986 VDDD.t1600 a_6077_9813.t38 clknet_1_1__leaf_CLK.t1 VDDD.t1599 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1987 VSSD.t1007 clknet_1_0__leaf_CLK.t54 a_9503_6037.t1 VSSD.t1006 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1988 VDDD.t756 a_1835_7637.t8 DOUT[9].t0 VDDD.t755 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1989 VDDD.t1602 a_6077_9813.t39 clknet_1_1__leaf_CLK.t0 VDDD.t1601 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1990 a_5746_3677.t3 a_5620_3579.t5 a_5342_3563.t3 VSSD.t1153 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1991 VDDD.t1175 VSSD.t1983 VDDD.t1174 VDDD.t1173 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1992 VSSD.t1655 CLKS.t132 a_4181_4399.t1 VSSD.t1654 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1993 a_7521_4399.t0 a_7477_4641.t5 a_7355_4399.t0 VSSD.t1089 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1994 a_4906_4943.t0 a_4187_5185.t7 a_4343_4917.t2 VSSD.t999 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1995 VDDD.t49 VSSD.t1984 VDDD.t48 VDDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1996 a_10145_4917.t2 a_9927_5321.t5 VSSD.t1017 VSSD.t1016 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1997 a_2439_5629.t0 CF[7].t8 VSSD.t324 VSSD.t323 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1998 clknet_1_0__leaf_CLK.t1 a_7654_4943.t36 VDDD.t349 VDDD.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1999 VSSD.t978 a_6813_7093.t39 clknet_0_CLK.t16 VSSD.t977 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2000 a_7801_8751.t0 CLKS.t133 VSSD.t1657 VSSD.t1656 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2001 a_1835_7637.t1 a_2122_7915.t5 VDDD.t18 VDDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2002 VDDD.t1651 a_7331_9269.t20 x3/COMP_BUF_N.t0 VDDD.t1650 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2003 a_6996_7663.t1 a_5915_7663.t7 a_6649_7905.t0 VDDD.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2004 a_5734_11471.t0 a_4976_11587.t5 a_5171_11445.t0 VDDD.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2005 VSSD.t1659 CLKS.t134 a_7705_3311.t1 VSSD.t1658 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2006 VDDD.t90 a_10584_3145.t5 a_10759_3071.t1 VDDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2007 VDDD.t164 a_4343_4917.t5 a_4274_4943.t0 VDDD.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2008 FINAL.t9 a_5307_7093.t19 VSSD.t154 VSSD.t153 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2009 CLKS.t14 x2/net13.t22 VDDD.t1406 VDDD.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2010 a_9832_5309.t2 CF[7].t9 VSSD.t326 VSSD.t325 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2011 VSSD.t1788 EN.t86 a_4733_11837.t1 VSSD.t1787 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2012 a_6999_8207.t1 EN.t87 VDDD.t673 VDDD.t672 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2013 a_3662_11471.t1 a_2585_11477.t5 a_3500_11849.t3 VDDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2014 VDDD.t52 VSSD.t1985 VDDD.t51 VDDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2015 SWP[6].t0 a_3859_4373.t8 VDDD.t470 VDDD.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2016 VDDD.t197 a_5307_7093.t20 FINAL.t0 VDDD.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2017 a_10654_9295.t1 a_9577_9301.t5 a_10492_9673.t3 VDDD.t763 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2018 a_8197_10389.t1 a_8031_10389.t7 VSSD.t141 VSSD.t140 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2019 VSSD.t294 a_2227_8988.t5 a_2158_9117.t3 VSSD.t293 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2020 VDDD.t60 x3/COMP_BUF_N.t35 a_5734_6031.t0 VDDD.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2021 clknet_1_0__leaf_CLK.t2 a_7654_4943.t37 VSSD.t277 VSSD.t276 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2022 a_4764_9117.t1 a_4550_9117.t5 VDDD.t1657 VDDD.t1656 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2023 a_10759_4159.t1 a_10584_4233.t5 a_10938_4221.t1 VSSD.t349 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2024 VDDD.t262 CLKS.t135 a_1835_5461.t0 VDDD.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2025 VSSD.t852 clknet_1_1__leaf_CLK.t55 a_2143_10389.t1 VSSD.t851 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2026 VSSD.t1582 a_6803_8725.t8 SWN[3].t2 VSSD.t1581 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X2027 a_9685_11169.t1 a_9467_10927.t5 VDDD.t1904 VDDD.t1903 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2028 a_4698_2899.t3 a_4976_2883.t5 a_4932_2767.t1 VDDD.t1880 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2029 VDDD.t55 VSSD.t1986 VDDD.t54 VDDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2030 DOUT[7].t0 a_1467_8181.t8 VDDD.t448 VDDD.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2031 VSSD.t218 CLKS.t136 a_10465_6575.t0 VSSD.t217 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2032 a_9563_8751.t0 a_9117_8751.t5 a_9467_8751.t0 VSSD.t724 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2033 VDDD.t1449 clknet_1_0__leaf_CLK.t55 a_9503_2773.t0 VDDD.t1448 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2034 a_4515_12381.t0 a_3891_12015.t7 a_4407_12015.t0 VDDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2035 VDDD.t264 CLKS.t137 a_4779_5461.t0 VDDD.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2036 a_5102_6031.t0 a_4976_6147.t5 a_4698_6163.t1 VSSD.t302 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2037 VSSD.t220 CLKS.t138 a_7797_6397.t0 VSSD.t219 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2038 VSSD.t222 CLKS.t139 a_4733_6397.t0 VSSD.t221 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2039 a_2157_5487.t1 a_2122_5739.t5 a_1835_5461.t2 VSSD.t438 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2040 VDDD.t351 a_7654_4943.t38 clknet_1_0__leaf_CLK.t3 VDDD.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2041 a_7443_10927.t2 a_7093_10927.t5 a_7348_10927.t2 VDDD.t886 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2042 a_2158_9117.t0 a_2032_9019.t5 a_1754_9003.t3 VSSD.t549 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2043 a_4619_4636.t2 a_4463_4541.t7 a_4764_4765.t1 VDDD.t788 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2044 a_10930_6941.t1 a_9853_6575.t5 a_10768_6575.t3 VDDD.t1883 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2045 FINAL.t8 a_5307_7093.t21 VSSD.t1093 VSSD.t1092 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2046 a_5416_10927.t1 x2/net1.t5 VSSD.t1805 VSSD.t1804 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2047 VSSD.t1188 VDDD.t2113 VSSD.t1187 VSSD.t1186 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2048 a_10329_3553.t2 a_10111_3311.t5 VSSD.t583 VSSD.t582 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2049 a_10237_2741.t3 a_10019_3145.t5 VDDD.t1721 VDDD.t1720 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2050 CF[3].t2 a_10759_3071.t8 VDDD.t1382 VDDD.t1381 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X2051 a_5015_6273.t1 CF[2].t9 VSSD.t957 VSSD.t956 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2052 x3/COMP_BUF_N.t8 a_7331_9269.t21 VSSD.t1643 VSSD.t1642 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2053 a_7091_11471.t2 EN.t88 VDDD.t675 VDDD.t674 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2054 a_10127_3855.t2 CLKS.t140 VDDD.t266 VDDD.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2055 a_7456_8585.t3 a_6541_8213.t5 a_7109_8181.t3 VSSD.t99 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2056 VSSD.t972 a_10207_7637.t8 a_10141_7663.t0 VSSD.t971 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2057 a_4411_6005.t2 a_4698_6163.t5 VDDD.t1716 VDDD.t1715 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2058 VDDD.t804 a_8183_3285.t8 CF[0].t3 VDDD.t803 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2059 VDDD.t58 VSSD.t1987 VDDD.t57 VDDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2060 a_10019_4233.t2 a_9669_3861.t5 a_9924_4221.t3 VDDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2061 VSSD.t1067 x2/net13.t23 CLKS.t15 VSSD.t1066 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2062 a_5101_5487.t0 a_5066_5739.t5 a_4779_5461.t2 VSSD.t753 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2063 a_4972_12015.t1 a_4057_12015.t5 a_4625_12257.t0 VSSD.t476 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2064 VDDD.t794 a_3031_10901.t8 x2/net9.t0 VDDD.t793 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2065 VSSD.t279 a_7654_4943.t39 clknet_1_0__leaf_CLK.t4 VSSD.t278 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2066 a_7091_11471.t1 a_6467_11477.t7 a_6983_11849.t3 VDDD.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2067 a_7574_6941.t3 a_6855_6717.t7 a_7011_6812.t2 VSSD.t1725 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2068 VSSD.t908 clknet_0_CLK.t47 a_6077_9813.t7 VSSD.t907 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2069 a_5182_4765.t3 a_4424_4667.t5 a_4619_4636.t1 VDDD.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2070 a_1973_5309.t1 a_1938_5075.t5 a_1651_4917.t2 VSSD.t1736 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2071 a_7245_11837.t0 a_7201_11445.t5 a_7079_11849.t1 VSSD.t1127 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2072 VSSD.t411 a_8183_10901.t8 a_8117_10927.t1 VSSD.t410 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2073 a_10601_9839.t0 a_9411_9839.t7 a_10492_9839.t0 VSSD.t139 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2074 a_2649_5309.t1 CLKS.t141 VSSD.t224 VSSD.t223 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2075 a_8008_10927.t3 a_6927_10927.t7 a_7661_11169.t2 VDDD.t1439 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2076 VSSD.t1185 VDDD.t2114 VSSD.t1184 VSSD.t1183 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2077 DOUT[8].t2 a_1467_8725.t8 VSSD.t343 VSSD.t342 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2078 a_10584_3145.t3 a_9503_2773.t7 a_10237_2741.t1 VDDD.t1891 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2079 a_2465_8573.t1 EN.t89 VSSD.t515 VSSD.t514 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2080 a_4380_9117.t0 a_3859_8725.t8 VDDD.t777 VDDD.t776 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2081 VSSD.t296 a_10851_5461.t8 a_10785_5487.t1 VSSD.t295 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
R0 a_2122_10091.n3 a_2122_10091.n2 636.953
R1 a_2122_10091.n1 a_2122_10091.t5 366.856
R2 a_2122_10091.n2 a_2122_10091.n0 300.2
R3 a_2122_10091.n2 a_2122_10091.n1 225.036
R4 a_2122_10091.n1 a_2122_10091.t4 174.056
R5 a_2122_10091.n0 a_2122_10091.t1 70.0005
R6 a_2122_10091.n3 a_2122_10091.t2 68.0124
R7 a_2122_10091.t0 a_2122_10091.n3 63.3219
R8 a_2122_10091.n0 a_2122_10091.t3 61.6672
R9 VDDD VDDD.t478 1725.39
R10 VDDD VDDD.t981 1719.47
R11 VDDD VDDD.t1027 1719.47
R12 VDDD.t1833 VDDD 1719.47
R13 VDDD.t1115 VDDD 1719.47
R14 VDDD VDDD.t1781 1719.47
R15 VDDD.t981 VDDD 1547.82
R16 VDDD.t1027 VDDD 1547.82
R17 VDDD VDDD.t1833 1547.82
R18 VDDD VDDD.t1115 1547.82
R19 VDDD.t478 VDDD 1547.82
R20 VDDD.t1781 VDDD 1547.82
R21 VDDD VDDD.t1041 975.178
R22 VDDD VDDD.t1071 975.178
R23 VDDD VDDD.t1033 975.178
R24 VDDD VDDD.t1147 975.178
R25 VDDD VDDD.t1750 975.178
R26 VDDD VDDD.t1787 975.178
R27 VDDD.t1041 VDDD 877.827
R28 VDDD.t1071 VDDD 877.827
R29 VDDD.t1033 VDDD 877.827
R30 VDDD.t1147 VDDD 877.827
R31 VDDD.t1750 VDDD 877.827
R32 VDDD.t1787 VDDD 877.827
R33 VDDD.n3426 VDDD.t816 877.144
R34 VDDD.n1568 VDDD.t516 812.014
R35 VDDD.n1134 VDDD.t1325 806.787
R36 VDDD.n313 VDDD.t204 806.511
R37 VDDD.n3596 VDDD.t1441 806.511
R38 VDDD.n3581 VDDD.t527 806.511
R39 VDDD.n3543 VDDD.t404 806.511
R40 VDDD.n3536 VDDD.t240 806.511
R41 VDDD.n3338 VDDD.t745 806.511
R42 VDDD.n3385 VDDD.t842 806.511
R43 VDDD.n697 VDDD.t1202 806.511
R44 VDDD.n741 VDDD.t466 806.511
R45 VDDD.n596 VDDD.t859 806.511
R46 VDDD.n1069 VDDD.t932 806.511
R47 VDDD.n1062 VDDD.t80 806.511
R48 VDDD.n886 VDDD.t558 806.511
R49 VDDD.n1013 VDDD.t1941 806.511
R50 VDDD.n971 VDDD.t1268 806.511
R51 VDDD.n1330 VDDD.t1246 806.511
R52 VDDD.n1397 VDDD.t1378 806.511
R53 VDDD.n2838 VDDD.t865 806.511
R54 VDDD.n1274 VDDD.t1876 806.511
R55 VDDD.n2764 VDDD.t1436 806.511
R56 VDDD.n2721 VDDD.t1210 806.511
R57 VDDD.n2720 VDDD.t1420 806.511
R58 VDDD.n2919 VDDD.t382 806.511
R59 VDDD.n1621 VDDD.t1649 806.511
R60 VDDD.n1578 VDDD.t164 806.511
R61 VDDD.n2657 VDDD.t667 806.511
R62 VDDD.n1906 VDDD.t603 806.511
R63 VDDD.n2342 VDDD.t750 806.511
R64 VDDD.n1668 VDDD.t162 806.511
R65 VDDD.n2389 VDDD.t1736 806.511
R66 VDDD.n3750 VDDD.t1612 806.511
R67 VDDD.n3173 VDDD.t1823 806.484
R68 VDDD.n8 VDDD.t480 804.731
R69 VDDD.n14 VDDD.t479 804.731
R70 VDDD.n3822 VDDD.t1783 804.731
R71 VDDD.n7 VDDD.t1782 804.731
R72 VDDD.n258 VDDD.t1857 804.731
R73 VDDD.n3510 VDDD.t1140 804.731
R74 VDDD.n224 VDDD.t1139 804.731
R75 VDDD.n334 VDDD.t495 804.731
R76 VDDD.n3605 VDDD.t494 804.731
R77 VDDD.n285 VDDD.t504 804.731
R78 VDDD.n3662 VDDD.t1760 804.731
R79 VDDD.n241 VDDD.t1759 804.731
R80 VDDD.t1080 VDDD.n234 804.731
R81 VDDD.t1858 VDDD.n254 804.731
R82 VDDD.n261 VDDD.t1040 804.731
R83 VDDD.n265 VDDD.t1005 804.731
R84 VDDD.n292 VDDD.t498 804.731
R85 VDDD.n287 VDDD.t1794 804.731
R86 VDDD.n295 VDDD.t1172 804.731
R87 VDDD.n298 VDDD.t1065 804.731
R88 VDDD.t1037 VDDD.n496 804.731
R89 VDDD.n505 VDDD.t977 804.731
R90 VDDD.n396 VDDD.t500 804.731
R91 VDDD.t1097 VDDD.n509 804.731
R92 VDDD.n3451 VDDD.t1785 804.731
R93 VDDD.t1786 VDDD.n3447 804.731
R94 VDDD.t1001 VDDD.n3301 804.731
R95 VDDD.n378 VDDD.t1143 804.731
R96 VDDD.n421 VDDD.t1142 804.731
R97 VDDD.n482 VDDD.t519 804.731
R98 VDDD.n400 VDDD.t492 804.731
R99 VDDD.n403 VDDD.t1738 804.731
R100 VDDD.n3352 VDDD.t1023 804.731
R101 VDDD.t1045 VDDD.n3344 804.731
R102 VDDD.n3355 VDDD.t985 804.731
R103 VDDD.n3358 VDDD.t513 804.731
R104 VDDD.n635 VDDD.t1829 804.731
R105 VDDD.n3187 VDDD.t1861 804.731
R106 VDDD.n3179 VDDD.t1860 804.731
R107 VDDD.n3222 VDDD.t1824 804.731
R108 VDDD.n3244 VDDD.t972 804.731
R109 VDDD.t1813 VDDD.n577 804.731
R110 VDDD.n658 VDDD.t1152 804.731
R111 VDDD.n720 VDDD.t1151 804.731
R112 VDDD.n639 VDDD.t1837 804.731
R113 VDDD.n672 VDDD.t1816 804.731
R114 VDDD.n675 VDDD.t1792 804.731
R115 VDDD.n3190 VDDD.t980 804.731
R116 VDDD.n3193 VDDD.t507 804.731
R117 VDDD.n776 VDDD.t1798 804.731
R118 VDDD.n779 VDDD.t1842 804.731
R119 VDDD.n765 VDDD.t1845 804.731
R120 VDDD.n790 VDDD.t1844 804.731
R121 VDDD.t995 VDDD.n784 804.731
R122 VDDD.n807 VDDD.t1113 804.731
R123 VDDD.n940 VDDD.t1803 804.731
R124 VDDD.n943 VDDD.t1017 804.731
R125 VDDD.n1441 VDDD.t1052 804.731
R126 VDDD.n1444 VDDD.t1847 804.731
R127 VDDD.n1170 VDDD.t1743 804.731
R128 VDDD.n1164 VDDD.t1742 804.731
R129 VDDD.n1170 VDDD.t1073 804.731
R130 VDDD.n1164 VDDD.t1072 804.731
R131 VDDD.n1163 VDDD.t1059 804.731
R132 VDDD.n1157 VDDD.t1058 804.731
R133 VDDD.n1163 VDDD.t1043 804.731
R134 VDDD.n1157 VDDD.t1042 804.731
R135 VDDD.n1156 VDDD.t489 804.731
R136 VDDD.n2974 VDDD.t488 804.731
R137 VDDD.t990 VDDD.n1335 804.731
R138 VDDD.n1173 VDDD.t1137 804.731
R139 VDDD.n1176 VDDD.t1032 804.731
R140 VDDD.n1263 VDDD.t55 804.731
R141 VDDD.n1299 VDDD.t1054 804.731
R142 VDDD.n1302 VDDD.t58 804.731
R143 VDDD.n2888 VDDD.t1146 804.731
R144 VDDD.n2891 VDDD.t1754 804.731
R145 VDDD.t1776 VDDD.n1570 804.731
R146 VDDD.t1062 VDDD.n2696 804.731
R147 VDDD.n1821 VDDD.t515 804.731
R148 VDDD.n1829 VDDD.t1049 804.731
R149 VDDD.n1761 VDDD.t1780 804.731
R150 VDDD.n1704 VDDD.t1779 804.731
R151 VDDD.n1728 VDDD.t521 804.731
R152 VDDD.n1737 VDDD.t522 804.731
R153 VDDD.n1693 VDDD.t486 804.731
R154 VDDD.n1696 VDDD.t993 804.731
R155 VDDD.n2629 VDDD.t1757 804.731
R156 VDDD.n2632 VDDD.t1826 804.731
R157 VDDD.n2507 VDDD.t1149 804.731
R158 VDDD.n2501 VDDD.t1148 804.731
R159 VDDD.n2507 VDDD.t1774 804.731
R160 VDDD.n2501 VDDD.t1773 804.731
R161 VDDD.n2500 VDDD.t1035 804.731
R162 VDDD.n2494 VDDD.t1034 804.731
R163 VDDD.n2500 VDDD.t1095 804.731
R164 VDDD.n2494 VDDD.t1094 804.731
R165 VDDD.n1892 VDDD.t999 804.731
R166 VDDD.n1895 VDDD.t1078 804.731
R167 VDDD.n1657 VDDD.t1122 804.731
R168 VDDD.n2447 VDDD.t1089 804.731
R169 VDDD.n1644 VDDD.t1090 804.731
R170 VDDD.n1934 VDDD.t1746 804.731
R171 VDDD.t1128 VDDD.n1936 804.731
R172 VDDD.n2510 VDDD.t1840 804.731
R173 VDDD.n2513 VDDD.t1167 804.731
R174 VDDD.n2062 VDDD.t1806 804.731
R175 VDDD.n2086 VDDD.t1805 804.731
R176 VDDD.n2061 VDDD.t1831 804.731
R177 VDDD.n2148 VDDD.t1832 804.731
R178 VDDD.n1989 VDDD.t1093 804.731
R179 VDDD.n1992 VDDD.t1811 804.731
R180 VDDD.n2242 VDDD.t1789 804.731
R181 VDDD.n2236 VDDD.t1788 804.731
R182 VDDD.n2242 VDDD.t1852 804.731
R183 VDDD.n2236 VDDD.t1851 804.731
R184 VDDD.n2235 VDDD.t1752 804.731
R185 VDDD.n2229 VDDD.t1751 804.731
R186 VDDD.n2235 VDDD.t1821 804.731
R187 VDDD.n2229 VDDD.t1820 804.731
R188 VDDD.n2225 VDDD.t1819 804.731
R189 VDDD.n2190 VDDD.t1818 804.731
R190 VDDD.n2034 VDDD.t1120 804.731
R191 VDDD.n2164 VDDD.t1119 804.731
R192 VDDD.n2162 VDDD.t1111 804.731
R193 VDDD.n1978 VDDD.t1772 804.731
R194 VDDD.n1970 VDDD.t1771 804.731
R195 VDDD.n1969 VDDD.t477 804.731
R196 VDDD.n2015 VDDD.t476 804.731
R197 VDDD.n1985 VDDD.t1155 804.731
R198 VDDD.t1025 VDDD.n2077 804.731
R199 VDDD.n2245 VDDD.t49 804.731
R200 VDDD.n2248 VDDD.t975 804.731
R201 VDDD.n71 VDDD.t1835 804.731
R202 VDDD.n52 VDDD.t1834 804.731
R203 VDDD.n46 VDDD.t1117 804.731
R204 VDDD.n72 VDDD.t1116 804.731
R205 VDDD.n199 VDDD.t983 804.731
R206 VDDD.n125 VDDD.t982 804.731
R207 VDDD.n178 VDDD.t1029 804.731
R208 VDDD.n172 VDDD.t1028 804.731
R209 VDDD.n327 VDDD.t1286 803.572
R210 VDDD.n3669 VDDD.t1904 803.572
R211 VDDD.n3429 VDDD.t846 803.572
R212 VDDD.n430 VDDD.t1936 803.572
R213 VDDD.n474 VDDD.t1329 803.572
R214 VDDD.n3214 VDDD.t370 803.572
R215 VDDD.n3139 VDDD.t1331 803.572
R216 VDDD.n3056 VDDD.t1902 803.572
R217 VDDD.n965 VDDD.t618 803.572
R218 VDDD.n1463 VDDD.t1698 803.572
R219 VDDD.n2832 VDDD.t1429 803.572
R220 VDDD.n2924 VDDD.t407 803.572
R221 VDDD.n1854 VDDD.t771 803.572
R222 VDDD.n1719 VDDD.t1356 803.572
R223 VDDD.n2662 VDDD.t946 803.572
R224 VDDD.n2435 VDDD.t20 803.572
R225 VDDD.n2430 VDDD.t82 803.572
R226 VDDD.n2120 VDDD.t754 803.572
R227 VDDD.n2036 VDDD.t224 803.572
R228 VDDD.n2002 VDDD.t1721 803.572
R229 VDDD.t1877 VDDD.t98 790.188
R230 VDDD.n1382 VDDD.t1505 783.403
R231 VDDD.n3446 VDDD.t456 780.471
R232 VDDD.n1735 VDDD.t355 779.372
R233 VDDD.n842 VDDD.t1410 777.706
R234 VDDD.n510 VDDD.t1097 751.957
R235 VDDD.t1857 VDDD.n257 751.692
R236 VDDD.n236 VDDD.t1080 751.692
R237 VDDD.n255 VDDD.t1858 751.692
R238 VDDD.t498 VDDD.n291 751.692
R239 VDDD.t1794 VDDD.n286 751.692
R240 VDDD.n497 VDDD.t1037 751.692
R241 VDDD.n3302 VDDD.t1001 751.692
R242 VDDD.t1023 VDDD.n3351 751.692
R243 VDDD.n3347 VDDD.t1045 751.692
R244 VDDD.t972 VDDD.n3243 751.692
R245 VDDD.n578 VDDD.t1813 751.692
R246 VDDD.t1837 VDDD.n638 751.692
R247 VDDD.n786 VDDD.t995 751.692
R248 VDDD.t1113 VDDD.n806 751.692
R249 VDDD.n1337 VDDD.t990 751.692
R250 VDDD.n1597 VDDD.t1776 751.692
R251 VDDD.n2697 VDDD.t1062 751.692
R252 VDDD.t1122 VDDD.n1656 751.692
R253 VDDD.t1746 VDDD.n1933 751.692
R254 VDDD.n1937 VDDD.t1128 751.692
R255 VDDD.t504 VDDD.n284 725.173
R256 VDDD.t1040 VDDD.n260 725.173
R257 VDDD.t1005 VDDD.n264 725.173
R258 VDDD.t1172 VDDD.n294 725.173
R259 VDDD.t1065 VDDD.n297 725.173
R260 VDDD.t977 VDDD.n504 725.173
R261 VDDD.t500 VDDD.n395 725.173
R262 VDDD.t1785 VDDD.n3450 725.173
R263 VDDD.n3448 VDDD.t1786 725.173
R264 VDDD.t519 VDDD.n481 725.173
R265 VDDD.t492 VDDD.n399 725.173
R266 VDDD.t1738 VDDD.n402 725.173
R267 VDDD.t985 VDDD.n3354 725.173
R268 VDDD.t513 VDDD.n3357 725.173
R269 VDDD.t1829 VDDD.n634 725.173
R270 VDDD.t1816 VDDD.n671 725.173
R271 VDDD.t1792 VDDD.n674 725.173
R272 VDDD.t980 VDDD.n3189 725.173
R273 VDDD.t507 VDDD.n3192 725.173
R274 VDDD.t1798 VDDD.n775 725.173
R275 VDDD.t1842 VDDD.n778 725.173
R276 VDDD.t1803 VDDD.n939 725.173
R277 VDDD.t1017 VDDD.n942 725.173
R278 VDDD.t1052 VDDD.n1440 725.173
R279 VDDD.t1847 VDDD.n1443 725.173
R280 VDDD.t1137 VDDD.n1172 725.173
R281 VDDD.t1032 VDDD.n1175 725.173
R282 VDDD.t55 VDDD.n1262 725.173
R283 VDDD.t1054 VDDD.n1298 725.173
R284 VDDD.t58 VDDD.n1301 725.173
R285 VDDD.t1146 VDDD.n2887 725.173
R286 VDDD.t1754 VDDD.n2890 725.173
R287 VDDD.t1049 VDDD.n1828 725.173
R288 VDDD.t486 VDDD.n1692 725.173
R289 VDDD.t993 VDDD.n1695 725.173
R290 VDDD.t1757 VDDD.n2628 725.173
R291 VDDD.t1826 VDDD.n2631 725.173
R292 VDDD.t999 VDDD.n1891 725.173
R293 VDDD.t1078 VDDD.n1894 725.173
R294 VDDD.t1840 VDDD.n2509 725.173
R295 VDDD.t1167 VDDD.n2512 725.173
R296 VDDD.t1093 VDDD.n1988 725.173
R297 VDDD.t1811 VDDD.n1991 725.173
R298 VDDD.t1111 VDDD.n2161 725.173
R299 VDDD.t1155 VDDD.n1984 725.173
R300 VDDD.n2078 VDDD.t1025 725.173
R301 VDDD.t49 VDDD.n2244 725.173
R302 VDDD.t975 VDDD.n2247 725.173
R303 VDDD.n1344 VDDD.t624 675.293
R304 VDDD.n1355 VDDD.t622 671.408
R305 VDDD.t1799 VDDD 669.701
R306 VDDD.n792 VDDD.t357 669.332
R307 VDDD.n3346 VDDD.t1358 668.764
R308 VDDD.n641 VDDD.t439 668.764
R309 VDDD.n955 VDDD.t1580 668.747
R310 VDDD.n350 VDDD.t1923 667.778
R311 VDDD.n3583 VDDD.t1694 667.778
R312 VDDD.n3372 VDDD.t1462 667.778
R313 VDDD.n3333 VDDD.t687 667.778
R314 VDDD.n456 VDDD.t1244 667.778
R315 VDDD.n3124 VDDD.t1952 667.778
R316 VDDD.n3045 VDDD.t1193 667.778
R317 VDDD.n883 VDDD.t417 667.778
R318 VDDD.n917 VDDD.t1707 667.778
R319 VDDD.n920 VDDD.t1214 667.778
R320 VDDD.n1368 VDDD.t415 667.778
R321 VDDD.n2801 VDDD.t60 667.778
R322 VDDD.n1251 VDDD.t1453 667.778
R323 VDDD.n2778 VDDD.t450 667.778
R324 VDDD.n2777 VDDD.t914 667.778
R325 VDDD.n1554 VDDD.t1643 667.778
R326 VDDD.n1553 VDDD.t958 667.778
R327 VDDD.n2934 VDDD.t831 667.778
R328 VDDD.n2932 VDDD.t1422 667.778
R329 VDDD.n1615 VDDD.t942 667.778
R330 VDDD.n2672 VDDD.t1451 667.778
R331 VDDD.n2670 VDDD.t1734 667.778
R332 VDDD.n1928 VDDD.t1630 667.778
R333 VDDD.n1952 VDDD.t34 667.778
R334 VDDD.n1665 VDDD.t1732 667.778
R335 VDDD.n3774 VDDD.t1878 667.778
R336 VDDD.n272 VDDD.t938 667.751
R337 VDDD.n3535 VDDD.t1703 667.751
R338 VDDD.n3419 VDDD.t620 667.751
R339 VDDD.n689 VDDD.t1208 667.751
R340 VDDD.n847 VDDD.t244 667.751
R341 VDDD.n893 VDDD.t452 667.751
R342 VDDD.n931 VDDD.t18 667.751
R343 VDDD.n1461 VDDD.t1431 667.751
R344 VDDD.n2816 VDDD.t1716 667.751
R345 VDDD.n2812 VDDD.t922 667.751
R346 VDDD.n2750 VDDD.t560 667.751
R347 VDDD.n2728 VDDD.t1350 667.751
R348 VDDD.n1809 VDDD.t1687 667.751
R349 VDDD.n1576 VDDD.t1212 667.751
R350 VDDD.n2350 VDDD.t1663 667.751
R351 VDDD.n1673 VDDD.t1892 667.751
R352 VDDD.n3742 VDDD.t1516 667.751
R353 VDDD.n305 VDDD.t588 666.404
R354 VDDD.n313 VDDD.t1177 666.366
R355 VDDD.n1330 VDDD.t214 666.366
R356 VDDD.n3606 VDDD.t97 664.455
R357 VDDD.n3637 VDDD.t472 664.455
R358 VDDD.n3565 VDDD.t851 664.455
R359 VDDD.n240 VDDD.t1366 664.455
R360 VDDD.n3511 VDDD.t634 664.455
R361 VDDD.n3396 VDDD.t85 664.455
R362 VDDD.n422 VDDD.t120 664.455
R363 VDDD.n461 VDDD.t1912 664.455
R364 VDDD.n3186 VDDD.t427 664.455
R365 VDDD.n683 VDDD.t586 664.455
R366 VDDD.n3256 VDDD.t605 664.455
R367 VDDD.n841 VDDD.t386 664.455
R368 VDDD.n998 VDDD.t1401 664.455
R369 VDDD.n1475 VDDD.t1541 664.455
R370 VDDD.n1230 VDDD.t1642 664.455
R371 VDDD.n1387 VDDD.t655 664.455
R372 VDDD.n1290 VDDD.t1932 664.455
R373 VDDD.n1307 VDDD.t342 664.455
R374 VDDD.n2875 VDDD.t879 664.455
R375 VDDD.n2910 VDDD.t590 664.455
R376 VDDD.n1780 VDDD.t464 664.455
R377 VDDD.n2599 VDDD.t1514 664.455
R378 VDDD.n2618 VDDD.t1863 664.455
R379 VDDD.n2648 VDDD.t1873 664.455
R380 VDDD.n2352 VDDD.t883 664.455
R381 VDDD.n2461 VDDD.t199 664.455
R382 VDDD.n2470 VDDD.t876 664.455
R383 VDDD.n1886 VDDD.t1305 664.455
R384 VDDD.n2058 VDDD.t1303 664.455
R385 VDDD.n2191 VDDD.t230 664.455
R386 VDDD.n2014 VDDD.t90 664.455
R387 VDDD.n479 VDDD.t692 664.069
R388 VDDD.n1493 VDDD.t155 664.069
R389 VDDD.n3298 VDDD.t1618 663.471
R390 VDDD.n3558 VDDD.t93 663.426
R391 VDDD.n3548 VDDD.t174 663.426
R392 VDDD.n3656 VDDD.t1196 663.426
R393 VDDD.n714 VDDD.t1483 663.426
R394 VDDD.n721 VDDD.t1376 663.426
R395 VDDD.n610 VDDD.t940 663.426
R396 VDDD.n3229 VDDD.t920 663.426
R397 VDDD.n857 VDDD.t818 663.426
R398 VDDD.n872 VDDD.t796 663.426
R399 VDDD.n879 VDDD.t1954 663.426
R400 VDDD.n1127 VDDD.t1950 663.426
R401 VDDD.n1822 VDDD.t1730 663.426
R402 VDDD.n1754 VDDD.t907 663.426
R403 VDDD.n1608 VDDD.t911 663.426
R404 VDDD.n2440 VDDD.t913 663.426
R405 VDDD.n2419 VDDD.t1299 663.426
R406 VDDD.n2407 VDDD.t572 663.426
R407 VDDD.n2107 VDDD.t62 663.426
R408 VDDD.n2041 VDDD.t1728 663.426
R409 VDDD.n2314 VDDD.t802 663.426
R410 VDDD VDDD.t1130 636.293
R411 VDDD.t711 VDDD.t1515 636.293
R412 VDDD.t1817 VDDD.t1807 617.668
R413 VDDD.n1403 VDDD.n1372 611.122
R414 VDDD.n1397 VDDD.n1379 611.122
R415 VDDD.n1687 VDDD.n1686 611.122
R416 VDDD.n530 VDDD.n520 610.861
R417 VDDD.n1396 VDDD.n1380 610.098
R418 VDDD.n1371 VDDD.n1370 609.615
R419 VDDD.n1410 VDDD.n1409 609.615
R420 VDDD.n518 VDDD.n517 609.37
R421 VDDD.n1809 VDDD.n1808 608.676
R422 VDDD.n3464 VDDD.n368 606.42
R423 VDDD.n525 VDDD.n523 606.42
R424 VDDD.n1377 VDDD.n1376 606.42
R425 VDDD.n1689 VDDD.n1688 606.42
R426 VDDD.n1801 VDDD.n1685 606.42
R427 VDDD.n1741 VDDD.n1736 605.581
R428 VDDD.n820 VDDD.n819 605.432
R429 VDDD.n838 VDDD.n827 605.432
R430 VDDD.n1084 VDDD.n839 605.432
R431 VDDD.n515 VDDD.n514 605.186
R432 VDDD.n540 VDDD.n512 605.186
R433 VDDD.n1364 VDDD.n1363 605.186
R434 VDDD.n1806 VDDD.n1683 605.186
R435 VDDD.n1862 VDDD.n1812 605.186
R436 VDDD.n320 VDDD.n319 604.457
R437 VDDD.n3568 VDDD.n3480 604.457
R438 VDDD.n3537 VDDD.n3493 604.457
R439 VDDD.n3421 VDDD.n3311 604.457
R440 VDDD.n465 VDDD.n464 604.457
R441 VDDD.n3146 VDDD.n644 604.457
R442 VDDD.n706 VDDD.n705 604.457
R443 VDDD.n1068 VDDD.n849 604.457
R444 VDDD.n1012 VDDD.n892 604.457
R445 VDDD.n957 VDDD.n932 604.457
R446 VDDD.n1456 VDDD.n1455 604.457
R447 VDDD.n2824 VDDD.n2814 604.457
R448 VDDD.n1277 VDDD.n1276 604.457
R449 VDDD.n2751 VDDD.n1289 604.457
R450 VDDD.n2727 VDDD.n1309 604.457
R451 VDDD.n2726 VDDD.n1310 604.457
R452 VDDD.n2917 VDDD.n2873 604.457
R453 VDDD.n2590 VDDD.n2589 604.457
R454 VDDD.n2655 VDDD.n2617 604.457
R455 VDDD.n1904 VDDD.n1903 604.457
R456 VDDD.n2349 VDDD.n2348 604.457
R457 VDDD.n2464 VDDD.n2463 604.457
R458 VDDD.n2468 VDDD.n2433 604.457
R459 VDDD.n2388 VDDD.n1672 604.457
R460 VDDD.n3744 VDDD.n33 604.457
R461 VDDD.n3597 VDDD.n349 604.394
R462 VDDD.n3580 VDDD.n357 604.394
R463 VDDD.n3485 VDDD.n3484 604.394
R464 VDDD.n734 VDDD.n716 604.394
R465 VDDD.n1055 VDDD.n859 604.394
R466 VDDD.n979 VDDD.n919 604.394
R467 VDDD.n2847 VDDD.n2846 604.394
R468 VDDD.n1265 VDDD.n1264 604.394
R469 VDDD.n2780 VDDD.n1267 604.394
R470 VDDD.n1531 VDDD.n1530 604.394
R471 VDDD.n1548 VDDD.n1532 604.394
R472 VDDD.n2939 VDDD.n1249 604.394
R473 VDDD.n2863 VDDD.n2862 604.394
R474 VDDD.n2677 VDDD.n2604 604.394
R475 VDDD.n2606 VDDD.n2605 604.394
R476 VDDD.n1945 VDDD.n1931 604.394
R477 VDDD.n1947 VDDD.n1946 604.394
R478 VDDD.n17 VDDD.n16 604.394
R479 VDDD.n3220 VDDD.n3219 604.011
R480 VDDD.n2163 VDDD.n2042 601.996
R481 VDDD.n3298 VDDD.n3297 601.926
R482 VDDD.n282 VDDD.n281 601.741
R483 VDDD.n322 VDDD.n321 601.679
R484 VDDD.n3590 VDDD.n3589 601.679
R485 VDDD.n355 VDDD.n354 601.679
R486 VDDD.n3491 VDDD.n3490 601.679
R487 VDDD.n3379 VDDD.n3378 601.679
R488 VDDD.n3336 VDDD.n3335 601.679
R489 VDDD.n709 VDDD.n708 601.679
R490 VDDD.n851 VDDD.n850 601.679
R491 VDDD.n1021 VDDD.n885 601.679
R492 VDDD.n889 VDDD.n888 601.679
R493 VDDD.n923 VDDD.n922 601.679
R494 VDDD.n926 VDDD.n925 601.679
R495 VDDD.n1458 VDDD.n1457 601.679
R496 VDDD.n2808 VDDD.n2807 601.679
R497 VDDD.n2804 VDDD.n2803 601.679
R498 VDDD.n2771 VDDD.n1272 601.679
R499 VDDD.n2769 VDDD.n1273 601.679
R500 VDDD.n1315 VDDD.n1314 601.679
R501 VDDD.n1526 VDDD.n1525 601.679
R502 VDDD.n2869 VDDD.n2868 601.679
R503 VDDD.n1591 VDDD.n1590 601.679
R504 VDDD.n1588 VDDD.n1587 601.679
R505 VDDD.n2612 VDDD.n2611 601.679
R506 VDDD.n1926 VDDD.n1914 601.679
R507 VDDD.n1917 VDDD.n1915 601.679
R508 VDDD.n2399 VDDD.n1667 601.679
R509 VDDD.n2392 VDDD.n2391 601.679
R510 VDDD.n3755 VDDD.n28 601.679
R511 VDDD.n1662 VDDD.n1660 601.359
R512 VDDD.n3603 VDDD.n3602 601.338
R513 VDDD.n2188 VDDD.n2187 601.338
R514 VDDD.n3269 VDDD.n3268 601.311
R515 VDDD.n1385 VDDD.n1384 601.311
R516 VDDD.n3643 VDDD.n3642 601.189
R517 VDDD.n1662 VDDD.n1661 601.112
R518 VDDD.n307 VDDD.n280 601.097
R519 VDDD.n3564 VDDD.n3481 601.097
R520 VDDD.n3650 VDDD.n227 601.097
R521 VDDD.n554 VDDD.n499 601.097
R522 VDDD.n3366 VDDD.n3343 601.097
R523 VDDD.n3330 VDDD.n3329 601.097
R524 VDDD.n463 VDDD.n375 601.097
R525 VDDD.n665 VDDD.n664 601.097
R526 VDDD.n724 VDDD.n722 601.097
R527 VDDD.n616 VDDD.n580 601.097
R528 VDDD.n3235 VDDD.n3174 601.097
R529 VDDD.n3038 VDDD.n772 601.097
R530 VDDD.n877 VDDD.n876 601.097
R531 VDDD.n1039 VDDD.n875 601.097
R532 VDDD.n882 VDDD.n881 601.097
R533 VDDD.n916 VDDD.n913 601.097
R534 VDDD.n1334 VDDD.n1333 601.097
R535 VDDD.n1367 VDDD.n1366 601.097
R536 VDDD.n1488 VDDD.n1339 601.097
R537 VDDD.n1125 VDDD.n1122 601.097
R538 VDDD.n2792 VDDD.n1258 601.097
R539 VDDD.n1826 VDDD.n1825 601.097
R540 VDDD.n1748 VDDD.n1732 601.097
R541 VDDD.n1601 VDDD.n1596 601.097
R542 VDDD.n1609 VDDD.n1594 601.097
R543 VDDD.n2575 VDDD.n1640 601.097
R544 VDDD.n2408 VDDD.n2406 601.097
R545 VDDD.n2308 VDDD.n1974 601.097
R546 VDDD.n3529 VDDD.n3497 600.105
R547 VDDD.n216 VDDD.n215 600.105
R548 VDDD.n3341 VDDD.n3340 600.105
R549 VDDD.n3391 VDDD.n3332 600.105
R550 VDDD.n389 VDDD.n388 600.105
R551 VDDD.n3207 VDDD.n3183 600.105
R552 VDDD.n688 VDDD.n687 600.105
R553 VDDD.n758 VDDD.n757 600.105
R554 VDDD.n846 VDDD.n845 600.105
R555 VDDD.n907 VDDD.n905 600.105
R556 VDDD.n964 VDDD.n928 600.105
R557 VDDD.n1450 VDDD.n1449 600.105
R558 VDDD.n1151 VDDD.n1149 600.105
R559 VDDD.n2831 VDDD.n2809 600.105
R560 VDDD.n2878 VDDD.n2877 600.105
R561 VDDD.n1863 VDDD.n1811 600.105
R562 VDDD.n1707 VDDD.n1706 600.105
R563 VDDD.n2595 VDDD.n1575 600.105
R564 VDDD.n2621 VDDD.n2620 600.105
R565 VDDD.n2370 VDDD.n1885 600.105
R566 VDDD.n2129 VDDD.n2060 600.105
R567 VDDD.n1998 VDDD.n1997 600.105
R568 VDDD.n279 VDDD.n278 598.383
R569 VDDD.n3549 VDDD.n3487 598.383
R570 VDDD.n220 VDDD.n219 598.383
R571 VDDD.n449 VDDD.n380 598.383
R572 VDDD.n3132 VDDD.n3131 598.383
R573 VDDD.n715 VDDD.n713 598.383
R574 VDDD.n591 VDDD.n588 598.383
R575 VDDD.n764 VDDD.n763 598.383
R576 VDDD.n858 VDDD.n856 598.383
R577 VDDD.n1498 VDDD.n1332 598.383
R578 VDDD.n1378 VDDD.n1375 598.383
R579 VDDD.n2981 VDDD.n1133 598.383
R580 VDDD.n2925 VDDD.n2870 598.383
R581 VDDD.n1849 VDDD.n1818 598.383
R582 VDDD.n1727 VDDD.n1718 598.383
R583 VDDD.n2663 VDDD.n2613 598.383
R584 VDDD.n2454 VDDD.n2437 598.383
R585 VDDD.n2477 VDDD.n2429 598.383
R586 VDDD.n2065 VDDD.n2064 598.383
R587 VDDD.n2176 VDDD.n2038 598.383
R588 VDDD.n1968 VDDD.n1967 598.383
R589 VDDD.n3290 VDDD.n3289 598.361
R590 VDDD.n3435 VDDD.n3434 598.237
R591 VDDD.n370 VDDD.n369 592.856
R592 VDDD.n2088 VDDD.n2087 592.159
R593 VDDD VDDD.t1853 588.942
R594 VDDD.t1611 VDDD.t638 583.023
R595 VDDD VDDD.t1848 568.994
R596 VDDD VDDD.t1112 568.994
R597 VDDD.n129 VDDD.t508 544.548
R598 VDDD.t1159 VDDD.n3707 544.548
R599 VDDD.t1074 VDDD 515.284
R600 VDDD.t1018 VDDD 511.926
R601 VDDD VDDD.t1156 494.238
R602 VDDD.t1276 VDDD.t1767 480.036
R603 VDDD.t1079 VDDD.t1856 463.252
R604 VDDD.t1060 VDDD.t1775 463.252
R605 VDDD.t1130 VDDD 458.724
R606 VDDD.t1454 VDDD.t1195 448.146
R607 VDDD.t1617 VDDD.t1274 448.146
R608 VDDD.t1359 VDDD.t1375 448.146
R609 VDDD.t1456 VDDD.t906 448.146
R610 VDDD.t825 VDDD.t912 448.146
R611 VDDD.t1688 VDDD.t801 448.146
R612 VDDD.t555 VDDD.t61 448.146
R613 VDDD.t1036 VDDD.t691 438.075
R614 VDDD.t1729 VDDD.t514 438.075
R615 VDDD.t1121 VDDD.t1298 438.075
R616 VDDD VDDD.t1018 414.577
R617 VDDD.t1623 VDDD.t100 414.33
R618 VDDD.n2945 VDDD.t1170 396.406
R619 VDDD.n2885 VDDD.t525 396.406
R620 VDDD.n1247 VDDD.t1169 391.005
R621 VDDD.n2884 VDDD.t524 391.005
R622 VDDD.n3172 VDDD.t1126 390.875
R623 VDDD.n3155 VDDD.t1838 390.875
R624 VDDD.n1248 VDDD.t483 390.062
R625 VDDD.n2557 VDDD.t1076 389.361
R626 VDDD.n1939 VDDD.t1129 389.361
R627 VDDD.n2023 VDDD.t1809 389.361
R628 VDDD.n289 VDDD.t1795 389.046
R629 VDDD.n3349 VDDD.t1046 389.046
R630 VDDD.n621 VDDD.t1850 389.046
R631 VDDD.n804 VDDD.t1114 389.046
R632 VDDD.n3241 VDDD.t973 388.721
R633 VDDD.n247 VDDD.t1081 388.656
R634 VDDD.n516 VDDD.t1098 388.656
R635 VDDD.n521 VDDD.t1762 388.656
R636 VDDD.n367 VDDD.t1763 388.656
R637 VDDD.n410 VDDD.t1765 388.656
R638 VDDD.n415 VDDD.t1766 388.656
R639 VDDD.n582 VDDD.t1814 388.656
R640 VDDD.n571 VDDD.t1125 388.656
R641 VDDD.n788 VDDD.t996 388.656
R642 VDDD.n873 VDDD.t1013 388.656
R643 VDDD.n1033 VDDD.t1014 388.656
R644 VDDD.n914 VDDD.t987 388.656
R645 VDDD.n984 VDDD.t988 388.656
R646 VDDD.n1476 VDDD.t1010 388.656
R647 VDDD.n1451 VDDD.t1011 388.656
R648 VDDD.n1390 VDDD.t1083 388.656
R649 VDDD.n1100 VDDD.t1084 388.656
R650 VDDD.n1131 VDDD.t1163 388.656
R651 VDDD.n2979 VDDD.t1164 388.656
R652 VDDD.n2786 VDDD.t1086 388.656
R653 VDDD.n1253 VDDD.t1087 388.656
R654 VDDD.n1535 VDDD.t1019 388.656
R655 VDDD.n1536 VDDD.t1020 388.656
R656 VDDD.n2880 VDDD.t1748 388.656
R657 VDDD.n2895 VDDD.t1749 388.656
R658 VDDD.n1602 VDDD.t1777 388.656
R659 VDDD.n2563 VDDD.t1075 388.656
R660 VDDD.n1649 VDDD.t1123 388.656
R661 VDDD.n2142 VDDD.t1768 388.656
R662 VDDD.n2148 VDDD.t1769 388.656
R663 VDDD.n2217 VDDD.t1808 388.656
R664 VDDD.n1977 VDDD.t1800 388.656
R665 VDDD.n2075 VDDD.t1801 388.656
R666 VDDD.n501 VDDD.t1038 388.656
R667 VDDD.n3304 VDDD.t1002 388.656
R668 VDDD.n3325 VDDD.t1007 388.656
R669 VDDD.n3401 VDDD.t1008 388.656
R670 VDDD.n470 VDDD.t51 388.656
R671 VDDD.n473 VDDD.t52 388.656
R672 VDDD.n669 VDDD.t1056 388.656
R673 VDDD.n681 VDDD.t1057 388.656
R674 VDDD.n935 VDDD.t1067 388.656
R675 VDDD.n948 VDDD.t1068 388.656
R676 VDDD.n1340 VDDD.t991 388.656
R677 VDDD.n1116 VDDD.t1174 388.656
R678 VDDD.n2999 VDDD.t1175 388.656
R679 VDDD.n2817 VDDD.t482 388.656
R680 VDDD.n1535 VDDD.t1069 388.656
R681 VDDD.n1536 VDDD.t1070 388.656
R682 VDDD.n1792 VDDD.t1740 388.656
R683 VDDD.n1703 VDDD.t1741 388.656
R684 VDDD.n2623 VDDD.t1134 388.656
R685 VDDD.n2626 VDDD.t1135 388.656
R686 VDDD.n3729 VDDD.t1131 388.656
R687 VDDD.n36 VDDD.t1132 388.656
R688 VDDD VDDD.t169 387.695
R689 VDDD.n290 VDDD.t497 387.682
R690 VDDD.n3350 VDDD.t1022 387.682
R691 VDDD.n1932 VDDD.t1745 387.682
R692 VDDD.n3157 VDDD.t1849 385.026
R693 VDDD.n2700 VDDD.t1061 385.026
R694 VDDD.n3828 VDDD.t1157 381.443
R695 VDDD.n50 VDDD.t1160 381.443
R696 VDDD.n3701 VDDD.t1161 381.443
R697 VDDD.n141 VDDD.t509 381.443
R698 VDDD.n126 VDDD.t510 381.443
R699 VDDD.n131 VDDD.t1854 381.443
R700 VDDD.n132 VDDD.t1855 381.443
R701 VDDD.n3831 VDDD.t1158 381.443
R702 VDDD.n507 VDDD.t978 381.44
R703 VDDD.n2080 VDDD.t1026 381.44
R704 VDDD.n393 VDDD.t501 381.44
R705 VDDD.n283 VDDD.t503 380.193
R706 VDDD.n259 VDDD.t1039 380.193
R707 VDDD.n263 VDDD.t1004 380.193
R708 VDDD.n293 VDDD.t1171 380.193
R709 VDDD.n296 VDDD.t1064 380.193
R710 VDDD.n480 VDDD.t518 380.193
R711 VDDD.n398 VDDD.t491 380.193
R712 VDDD.n401 VDDD.t1737 380.193
R713 VDDD.n3353 VDDD.t984 380.193
R714 VDDD.n3356 VDDD.t512 380.193
R715 VDDD.n633 VDDD.t1828 380.193
R716 VDDD.n670 VDDD.t1815 380.193
R717 VDDD.n673 VDDD.t1791 380.193
R718 VDDD.n3188 VDDD.t979 380.193
R719 VDDD.n3191 VDDD.t506 380.193
R720 VDDD.n774 VDDD.t1797 380.193
R721 VDDD.n777 VDDD.t1841 380.193
R722 VDDD.n938 VDDD.t1802 380.193
R723 VDDD.n941 VDDD.t1016 380.193
R724 VDDD.n1439 VDDD.t1051 380.193
R725 VDDD.n1442 VDDD.t1846 380.193
R726 VDDD.n1171 VDDD.t1136 380.193
R727 VDDD.n1174 VDDD.t1031 380.193
R728 VDDD.n1261 VDDD.t54 380.193
R729 VDDD.n1297 VDDD.t1053 380.193
R730 VDDD.n1300 VDDD.t57 380.193
R731 VDDD.n2886 VDDD.t1145 380.193
R732 VDDD.n2889 VDDD.t1753 380.193
R733 VDDD.n1827 VDDD.t1048 380.193
R734 VDDD.n1691 VDDD.t485 380.193
R735 VDDD.n1694 VDDD.t992 380.193
R736 VDDD.n2627 VDDD.t1756 380.193
R737 VDDD.n2630 VDDD.t1825 380.193
R738 VDDD.n1890 VDDD.t998 380.193
R739 VDDD.n1893 VDDD.t1077 380.193
R740 VDDD.n2508 VDDD.t1839 380.193
R741 VDDD.n2511 VDDD.t1166 380.193
R742 VDDD.n1987 VDDD.t1092 380.193
R743 VDDD.n1990 VDDD.t1810 380.193
R744 VDDD.n2160 VDDD.t1110 380.193
R745 VDDD.n1983 VDDD.t1154 380.193
R746 VDDD.n2243 VDDD.t48 380.193
R747 VDDD.n2246 VDDD.t974 380.193
R748 VDDD VDDD.t689 367.579
R749 VDDD.t961 VDDD.t633 360.866
R750 VDDD.t96 VDDD.t1336 360.866
R751 VDDD.t896 VDDD.t471 360.866
R752 VDDD.t774 VDDD.t604 360.866
R753 VDDD.t426 VDDD.t372 360.866
R754 VDDD.t1579 VDDD.t943 360.866
R755 VDDD.t463 VDDD.t1342 360.866
R756 VDDD.t1302 VDDD.t1280 360.866
R757 VDDD.t229 VDDD.t751 360.866
R758 VDDD VDDD.t1563 357.51
R759 VDDD.t1744 VDDD 357.51
R760 VDDD VDDD.t1219 354.152
R761 VDDD.n815 VDDD.t366 347.019
R762 VDDD.n3482 VDDD.t610 343.579
R763 VDDD.n3081 VDDD.t874 343.579
R764 VDDD.n1073 VDDD.t1557 343.579
R765 VDDD.n958 VDDD.t756 343.579
R766 VDDD.n1437 VDDD.t596 343.579
R767 VDDD.n2825 VDDD.t536 343.579
R768 VDDD.n2734 VDDD.t1293 343.579
R769 VDDD.n1900 VDDD.t1412 343.579
R770 VDDD.n34 VDDD.t712 343.579
R771 VDDD.n3495 VDDD.t1921 343.577
R772 VDDD.n376 VDDD.t836 343.577
R773 VDDD.n3090 VDDD.t1948 343.577
R774 VDDD.n908 VDDD.t12 343.577
R775 VDDD.n2819 VDDD.t68 343.577
R776 VDDD.n2744 VDDD.t1234 343.577
R777 VDDD.n3010 VDDD.t1384 340.344
R778 VDDD.n1785 VDDD.t1343 340.303
R779 VDDD.n329 VDDD.t790 340.012
R780 VDDD.n246 VDDD.t564 340.012
R781 VDDD.n3508 VDDD.t962 340.012
R782 VDDD.n414 VDDD.t1655 340.012
R783 VDDD.n3345 VDDD.t1220 340.012
R784 VDDD.n3200 VDDD.t373 340.012
R785 VDDD.n640 VDDD.t1564 340.012
R786 VDDD.n574 VDDD.t775 340.012
R787 VDDD.n797 VDDD.t1290 340.012
R788 VDDD.n1000 VDDD.t1889 340.012
R789 VDDD.n1153 VDDD.t1104 340.012
R790 VDDD.n2745 VDDD.t202 340.012
R791 VDDD.n2905 VDDD.t72 340.012
R792 VDDD.n1807 VDDD.t741 340.012
R793 VDDD.n2597 VDDD.t1185 340.012
R794 VDDD.n2649 VDDD.t409 340.012
R795 VDDD.n2456 VDDD.t857 340.012
R796 VDDD.n2368 VDDD.t665 340.012
R797 VDDD.n3612 VDDD.t1337 340.01
R798 VDDD.n336 VDDD.t897 340.01
R799 VDDD.n3324 VDDD.t118 340.01
R800 VDDD.n3400 VDDD.t176 340.01
R801 VDDD.n1083 VDDD.t1309 340.01
R802 VDDD.n950 VDDD.t944 340.01
R803 VDDD.n1454 VDDD.t1418 340.01
R804 VDDD.n2733 VDDD.t379 340.01
R805 VDDD.n2911 VDDD.t102 340.01
R806 VDDD.n1573 VDDD.t552 340.01
R807 VDDD.n2643 VDDD.t1705 340.01
R808 VDDD.n1902 VDDD.t833 340.01
R809 VDDD.n2475 VDDD.t707 340.01
R810 VDDD.n1887 VDDD.t246 340.01
R811 VDDD.n2137 VDDD.t1281 340.01
R812 VDDD.n2197 VDDD.t752 340.01
R813 VDDD.n1982 VDDD.t1382 340.01
R814 VDDD VDDD.n3170 339.046
R815 VDDD VDDD.n810 339.046
R816 VDDD.n548 VDDD.t38 339.002
R817 VDDD.n595 VDDD.t724 338.892
R818 VDDD.n583 VDDD.t722 338.108
R819 VDDD.n1346 VDDD.t855 336.522
R820 VDDD.n1817 VDDD.t26 336.522
R821 VDDD VDDD.t1003 334.012
R822 VDDD VDDD.t490 334.012
R823 VDDD VDDD.t1790 334.012
R824 VDDD VDDD.t1796 334.012
R825 VDDD VDDD.t1050 334.012
R826 VDDD VDDD.t56 334.012
R827 VDDD VDDD.t484 334.012
R828 VDDD VDDD.t997 334.012
R829 VDDD VDDD.t1091 334.012
R830 VDDD VDDD.t1727 332.332
R831 VDDD.t1591 VDDD.t1903 330.654
R832 VDDD.t526 VDDD.t1480 330.654
R833 VDDD.t658 VDDD.t1440 330.654
R834 VDDD.t203 VDDD.t1589 330.654
R835 VDDD.t1935 VDDD.t1868 330.654
R836 VDDD.t1251 VDDD.t369 330.654
R837 VDDD.t1478 VDDD.t1245 330.654
R838 VDDD.t307 VDDD.t1355 330.654
R839 VDDD.t303 VDDD.t1720 330.654
R840 VDDD.t331 VDDD.t753 330.654
R841 VDDD.t1241 VDDD.t223 330.654
R842 VDDD.t69 VDDD.t1747 325.618
R843 VDDD.n3030 VDDD.n817 323.053
R844 VDDD.t508 VDDD 322.587
R845 VDDD VDDD.t1159 322.587
R846 VDDD.t1156 VDDD 322.587
R847 VDDD.n1430 VDDD.n1345 322.329
R848 VDDD.n1436 VDDD.n1342 322.329
R849 VDDD.t11 VDDD.t1884 322.262
R850 VDDD.n3309 VDDD.n3308 320.976
R851 VDDD.n657 VDDD.n656 320.976
R852 VDDD.n3129 VDDD.n653 320.976
R853 VDDD.n604 VDDD.n585 320.976
R854 VDDD.n590 VDDD.n589 320.976
R855 VDDD.n598 VDDD.n592 320.976
R856 VDDD.n3044 VDDD.n767 320.976
R857 VDDD.n771 VDDD.n770 320.976
R858 VDDD.n3007 VDDD.n1112 320.976
R859 VDDD.n1118 VDDD.n1115 320.976
R860 VDDD.t1396 VDDD.t171 319.627
R861 VDDD VDDD.t1715 317.226
R862 VDDD.n3709 VDDD 316.668
R863 VDDD.n3708 VDDD 316.668
R864 VDDD.t835 VDDD.t1924 315.548
R865 VDDD.n1417 VDDD.n1416 315.334
R866 VDDD.n1814 VDDD.n1813 315.334
R867 VDDD.n544 VDDD.n543 313.897
R868 VDDD.n503 VDDD.n502 311.983
R869 VDDD.n1353 VDDD.n1352 311.149
R870 VDDD.n1855 VDDD.n1816 311.149
R871 VDDD.n647 VDDD.n646 310.5
R872 VDDD.n2993 VDDD.n1126 310.5
R873 VDDD.t1793 VDDD.t496 308.834
R874 VDDD.t1044 VDDD.t1021 308.834
R875 VDDD.n2294 VDDD.t1024 308.834
R876 VDDD.n3138 VDDD.n649 307.204
R877 VDDD.n651 VDDD.n650 307.204
R878 VDDD.n3036 VDDD.n773 307.204
R879 VDDD.n816 VDDD.n814 307.204
R880 VDDD.n3028 VDDD.n818 307.204
R881 VDDD.n3000 VDDD.n1119 307.204
R882 VDDD.n1124 VDDD.n1123 307.204
R883 VDDD.t1285 VDDD.t937 307.156
R884 VDDD.t1430 VDDD.t1697 307.156
R885 VDDD.n5 VDDD.t1998 306.735
R886 VDDD.n12 VDDD.t2059 306.735
R887 VDDD.n3613 VDDD.t2091 306.735
R888 VDDD.n3675 VDDD.t2013 306.735
R889 VDDD.n225 VDDD.t2060 306.735
R890 VDDD.n428 VDDD.t2062 306.735
R891 VDDD.n3181 VDDD.t1982 306.735
R892 VDDD.n723 VDDD.t2065 306.735
R893 VDDD.n3236 VDDD.t2111 306.735
R894 VDDD.n759 VDDD.t2009 306.735
R895 VDDD.n1150 VDDD.t1980 306.735
R896 VDDD.n1159 VDDD.t1994 306.735
R897 VDDD.n1159 VDDD.t2030 306.735
R898 VDDD.n1166 VDDD.t2006 306.735
R899 VDDD.n1166 VDDD.t2045 306.735
R900 VDDD.n1824 VDDD.t1997 306.735
R901 VDDD.n1730 VDDD.t2109 306.735
R902 VDDD.n1709 VDDD.t2032 306.735
R903 VDDD.n2441 VDDD.t2020 306.735
R904 VDDD.n2496 VDDD.t2022 306.735
R905 VDDD.n2496 VDDD.t2093 306.735
R906 VDDD.n2503 VDDD.t2041 306.735
R907 VDDD.n2503 VDDD.t2107 306.735
R908 VDDD.n2131 VDDD.t1992 306.735
R909 VDDD.n2108 VDDD.t2114 306.735
R910 VDDD.n2170 VDDD.t2073 306.735
R911 VDDD.n2198 VDDD.t1983 306.735
R912 VDDD.n2008 VDDD.t2102 306.735
R913 VDDD.n1972 VDDD.t2039 306.735
R914 VDDD.n2231 VDDD.t1985 306.735
R915 VDDD.n2231 VDDD.t2015 306.735
R916 VDDD.n2238 VDDD.t1996 306.735
R917 VDDD.n2238 VDDD.t2033 306.735
R918 VDDD.n74 VDDD.t2029 306.735
R919 VDDD.n107 VDDD.t2092 306.735
R920 VDDD.n174 VDDD.t2027 306.735
R921 VDDD.n123 VDDD.t2007 306.735
R922 VDDD.t1103 VDDD.t487 305.478
R923 VDDD.t1913 VDDD.t957 293.728
R924 VDDD.t449 VDDD.t5 293.728
R925 VDDD.t1391 VDDD.t1629 293.728
R926 VDDD.t1346 VDDD.t1611 292.991
R927 VDDD.t100 VDDD.t637 292.991
R928 VDDD.t638 VDDD.t1623 287.072
R929 VDDD.t1822 VDDD.t919 283.658
R930 VDDD.t989 VDDD.t154 283.658
R931 VDDD VDDD.t1063 280.3
R932 VDDD.t976 VDDD 280.3
R933 VDDD VDDD.t511 280.3
R934 VDDD VDDD.t505 280.3
R935 VDDD VDDD.t1015 280.3
R936 VDDD VDDD.t1030 280.3
R937 VDDD VDDD.t53 280.3
R938 VDDD VDDD.t1144 280.3
R939 VDDD VDDD.t1047 280.3
R940 VDDD VDDD.t1165 280.3
R941 VDDD VDDD.t47 280.3
R942 VDDD VDDD.t1755 278.623
R943 VDDD VDDD.t696 273.587
R944 VDDD.t637 VDDD.t1877 272.274
R945 VDDD.t1691 VDDD 270.231
R946 VDDD VDDD.t1906 270.231
R947 VDDD.t1150 VDDD 261.837
R948 VDDD.t1540 VDDD 261.837
R949 VDDD.t496 VDDD 260.159
R950 VDDD.t1021 VDDD 260.159
R951 VDDD.t971 VDDD 260.159
R952 VDDD.t986 VDDD 260.159
R953 VDDD.t1082 VDDD 260.159
R954 VDDD VDDD.t1168 260.159
R955 VDDD.t523 VDDD 260.159
R956 VDDD.t1133 VDDD 260.159
R957 VDDD.t1767 VDDD 260.159
R958 VDDD.t1807 VDDD 260.159
R959 VDDD.t1365 VDDD 258.481
R960 VDDD VDDD.t119 258.481
R961 VDDD.t89 VDDD 258.481
R962 VDDD VDDD.t1289 256.803
R963 VDDD.n518 VDDD.t76 255.154
R964 VDDD.t1525 VDDD.t1346 254.518
R965 VDDD.n3428 VDDD.t1616 250.724
R966 VDDD.n684 VDDD.t324 250.724
R967 VDDD.n270 VDDD.t794 250.464
R968 VDDD.n956 VDDD.t1536 250.464
R969 VDDD.n1438 VDDD.t956 250.464
R970 VDDD.n3008 VDDD.t739 250.464
R971 VDDD.n2813 VDDD.t538 250.464
R972 VDDD.n2743 VDDD.t1264 250.464
R973 VDDD.n3736 VDDD.t170 250.464
R974 VDDD.n455 VDDD.t838 250.463
R975 VDDD.n1468 VDDD.t1414 250.463
R976 VDDD.n2735 VDDD.t377 250.463
R977 VDDD.n2357 VDDD.t375 250.463
R978 VDDD.n2677 VDDD.t548 249.407
R979 VDDD.n3420 VDDD.t814 248.843
R980 VDDD.t169 VDDD.t711 248.599
R981 VDDD.t1515 VDDD.t1396 248.599
R982 VDDD.t171 VDDD.t1525 248.599
R983 VDDD.t98 VDDD.t893 248.599
R984 VDDD.n3647 VDDD.t45 248.411
R985 VDDD.n3171 VDDD.t947 248.411
R986 VDDD.n1155 VDDD.t1105 248.411
R987 VDDD.t469 VDDD.n2682 248.411
R988 VDDD.n2361 VDDD.t803 248.411
R989 VDDD.t81 VDDD.t706 248.411
R990 VDDD.t856 VDDD.t19 248.411
R991 VDDD.t1379 VDDD.n2021 248.411
R992 VDDD.n3305 VDDD.t1614 248.219
R993 VDDD.n504 VDDD.t2034 247.744
R994 VDDD.n2078 VDDD.t2066 247.744
R995 VDDD.n1940 VDDD.t616 247.293
R996 VDDD.n395 VDDD.t2078 246.734
R997 VDDD.n3557 VDDD.t608 246.112
R998 VDDD.n249 VDDD.t566 246.112
R999 VDDD.n3504 VDDD.t46 246.112
R1000 VDDD.n413 VDDD.t1653 246.112
R1001 VDDD.n3345 VDDD.t1216 246.112
R1002 VDDD.n3187 VDDD.t840 246.112
R1003 VDDD.n640 VDDD.t1568 246.112
R1004 VDDD.n685 VDDD.t1620 246.112
R1005 VDDD.n3250 VDDD.t948 246.112
R1006 VDDD.n799 VDDD.t1311 246.112
R1007 VDDD.n843 VDDD.t716 246.112
R1008 VDDD.n997 VDDD.t1885 246.112
R1009 VDDD.n1224 VDDD.t1106 246.112
R1010 VDDD.n1296 VDDD.t1930 246.112
R1011 VDDD.n2881 VDDD.t70 246.112
R1012 VDDD.n1684 VDDD.t628 246.112
R1013 VDDD.n2598 VDDD.t470 246.112
R1014 VDDD.n2622 VDDD.t390 246.112
R1015 VDDD.n2358 VDDD.t444 246.112
R1016 VDDD.n2453 VDDD.t1 246.112
R1017 VDDD.n2363 VDDD.t804 246.112
R1018 VDDD.n3614 VDDD.t936 246.111
R1019 VDDD.n3631 VDDD.t899 246.111
R1020 VDDD.n3528 VDDD.t970 246.111
R1021 VDDD.n3407 VDDD.t116 246.111
R1022 VDDD.n3326 VDDD.t251 246.111
R1023 VDDD.n680 VDDD.t1323 246.111
R1024 VDDD.n948 VDDD.t448 246.111
R1025 VDDD.n1086 VDDD.t1307 246.111
R1026 VDDD.n991 VDDD.t8 246.111
R1027 VDDD.n1243 VDDD.t697 246.111
R1028 VDDD.n2742 VDDD.t1236 246.111
R1029 VDDD.n2879 VDDD.t1970 246.111
R1030 VDDD.n1702 VDDD.t1606 246.111
R1031 VDDD.n2625 VDDD.t1270 246.111
R1032 VDDD.n2478 VDDD.t1341 246.111
R1033 VDDD.n2056 VDDD.t1277 246.111
R1034 VDDD.n2199 VDDD.t705 246.111
R1035 VDDD.n1982 VDDD.t1380 246.111
R1036 VDDD.n284 VDDD.t2097 245.667
R1037 VDDD.n260 VDDD.t1987 245.667
R1038 VDDD.n264 VDDD.t2052 245.667
R1039 VDDD.n294 VDDD.t2074 245.667
R1040 VDDD.n297 VDDD.t2001 245.667
R1041 VDDD.n481 VDDD.t2010 245.667
R1042 VDDD.n399 VDDD.t2084 245.667
R1043 VDDD.n402 VDDD.t2064 245.667
R1044 VDDD.n3354 VDDD.t2037 245.667
R1045 VDDD.n3357 VDDD.t1995 245.667
R1046 VDDD.n634 VDDD.t2014 245.667
R1047 VDDD.n671 VDDD.t2104 245.667
R1048 VDDD.n674 VDDD.t2067 245.667
R1049 VDDD.n3189 VDDD.t2035 245.667
R1050 VDDD.n3192 VDDD.t2000 245.667
R1051 VDDD.n775 VDDD.t2063 245.667
R1052 VDDD.n778 VDDD.t2031 245.667
R1053 VDDD.n939 VDDD.t1993 245.667
R1054 VDDD.n942 VDDD.t2101 245.667
R1055 VDDD.n1440 VDDD.t2023 245.667
R1056 VDDD.n1443 VDDD.t1991 245.667
R1057 VDDD.n1172 VDDD.t2096 245.667
R1058 VDDD.n1175 VDDD.t2058 245.667
R1059 VDDD.n1262 VDDD.t2088 245.667
R1060 VDDD.n1298 VDDD.t2026 245.667
R1061 VDDD.n1301 VDDD.t2090 245.667
R1062 VDDD.n2887 VDDD.t2098 245.667
R1063 VDDD.n2890 VDDD.t2019 245.667
R1064 VDDD.n1828 VDDD.t1999 245.667
R1065 VDDD.n1692 VDDD.t1989 245.667
R1066 VDDD.n1695 VDDD.t2053 245.667
R1067 VDDD.n2628 VDDD.t2056 245.667
R1068 VDDD.n2631 VDDD.t1981 245.667
R1069 VDDD.n1891 VDDD.t2087 245.667
R1070 VDDD.n1894 VDDD.t2017 245.667
R1071 VDDD.n2509 VDDD.t2011 245.667
R1072 VDDD.n2512 VDDD.t2089 245.667
R1073 VDDD.n1988 VDDD.t2008 245.667
R1074 VDDD.n1991 VDDD.t1979 245.667
R1075 VDDD.n2161 VDDD.t2070 245.667
R1076 VDDD.n1984 VDDD.t2086 245.667
R1077 VDDD.n2244 VDDD.t2082 245.667
R1078 VDDD.n2247 VDDD.t2051 245.667
R1079 VDDD.n3145 VDDD.t1638 243.512
R1080 VDDD.n3829 VDDD.t2047 242.282
R1081 VDDD.n51 VDDD.t2048 242.282
R1082 VDDD.n142 VDDD.t2072 242.282
R1083 VDDD.n133 VDDD.t2099 242.282
R1084 VDDD.n828 VDDD.t926 240.214
R1085 VDDD.n2988 VDDD.t147 240.214
R1086 VDDD.n3449 VDDD.t2021 238.976
R1087 VDDD.t354 VDDD 236.661
R1088 VDDD.n3243 VDDD.t2075 235.319
R1089 VDDD.t1508 VDDD.t678 234.982
R1090 VDDD.t94 VDDD.t1262 234.982
R1091 VDDD.t848 VDDD.t1229 234.982
R1092 VDDD.t847 VDDD.t269 234.982
R1093 VDDD.t1230 VDDD.t811 234.982
R1094 VDDD.t713 VDDD.t1939 234.982
R1095 VDDD.t1402 VDDD.t121 234.982
R1096 VDDD.t1695 VDDD.t1683 234.982
R1097 VDDD.t1684 VDDD.t206 234.982
R1098 VDDD.t1463 VDDD.t772 234.982
R1099 VDDD.t1363 VDDD.t380 234.982
R1100 VDDD.t1890 VDDD.t383 234.982
R1101 VDDD.t734 VDDD.t43 234.982
R1102 VDDD.t323 VDDD.t1947 233.304
R1103 VDDD.t1259 VDDD.t1843 233.304
R1104 VDDD.t1510 VDDD.t1437 231.625
R1105 VDDD.t185 VDDD.t1205 231.625
R1106 VDDD.t1836 VDDD.t1827 231.625
R1107 VDDD.t220 VDDD.t929 231.625
R1108 VDDD.n129 VDDD 227.882
R1109 VDDD VDDD.n3708 227.882
R1110 VDDD.t1853 VDDD 221.964
R1111 VDDD.n3707 VDDD 221.964
R1112 VDDD.n3709 VDDD 221.964
R1113 VDDD.t1804 VDDD.t808 221.555
R1114 VDDD.t565 VDDD 219.876
R1115 VDDD VDDD.t601 219.876
R1116 VDDD.t615 VDDD 219.876
R1117 VDDD.t112 VDDD 216.519
R1118 VDDD.n291 VDDD.t2094 213.148
R1119 VDDD.n3351 VDDD.t2085 213.148
R1120 VDDD.n1933 VDDD.t2054 213.148
R1121 VDDD.n3646 VDDD.n269 213.119
R1122 VDDD.n3462 VDDD.n3293 213.119
R1123 VDDD.n1482 VDDD.n1481 213.119
R1124 VDDD.n3009 VDDD.n1101 213.119
R1125 VDDD.n2860 VDDD.n2859 213.119
R1126 VDDD.n2492 VDDD.n2491 213.119
R1127 VDDD.n3645 VDDD.n3644 213.119
R1128 VDDD.n1796 VDDD.n1795 213.119
R1129 VDDD.n3708 VDDD.n15 213.119
R1130 VDDD.n3715 VDDD.n3709 213.119
R1131 VDDD.n3707 VDDD.n3706 213.119
R1132 VDDD.n139 VDDD.n129 213.119
R1133 VDDD.n2939 VDDD.n2861 212.665
R1134 VDDD.n522 VDDD.t2016 210.964
R1135 VDDD.n411 VDDD.t2018 210.964
R1136 VDDD.n471 VDDD.t1986 210.964
R1137 VDDD.n679 VDDD.t2038 210.964
R1138 VDDD.n915 VDDD.t2069 210.964
R1139 VDDD.n937 VDDD.t2050 210.964
R1140 VDDD.n1474 VDDD.t2079 210.964
R1141 VDDD.n1389 VDDD.t2040 210.964
R1142 VDDD.n1117 VDDD.t2083 210.964
R1143 VDDD.n1132 VDDD.t2106 210.964
R1144 VDDD.n1247 VDDD.t2108 210.964
R1145 VDDD.n2884 VDDD.t2112 210.964
R1146 VDDD.n1791 VDDD.t2012 210.964
R1147 VDDD.n2624 VDDD.t2068 210.964
R1148 VDDD.n2055 VDDD.t2025 210.964
R1149 VDDD.n3730 VDDD.t2036 210.964
R1150 VDDD.n397 VDDD.t499 210.55
R1151 VDDD.n2556 VDDD.n2493 210.55
R1152 VDDD.n2292 VDDD.n2291 210.55
R1153 VDDD.n2692 VDDD.n2683 210.365
R1154 VDDD.n268 VDDD.n267 210.155
R1155 VDDD.n3170 VDDD.n3169 210.144
R1156 VDDD.n810 VDDD.n809 210.012
R1157 VDDD.n3648 VDDD.n3647 209.368
R1158 VDDD.n3398 VDDD.n3397 209.368
R1159 VDDD.n3292 VDDD.n3291 209.368
R1160 VDDD.n3248 VDDD.n3171 209.368
R1161 VDDD.n3101 VDDD.n3100 209.368
R1162 VDDD.n3099 VDDD.n3098 209.368
R1163 VDDD.n990 VDDD.n910 209.368
R1164 VDDD.n3035 VDDD.n811 209.368
R1165 VDDD.n909 VDDD.n861 209.368
R1166 VDDD.n1222 VDDD.n1155 209.368
R1167 VDDD.n1483 VDDD.t241 209.368
R1168 VDDD.n2741 VDDD.n2740 209.368
R1169 VDDD.n2739 VDDD.n2738 209.368
R1170 VDDD.n2682 VDDD.n2681 209.368
R1171 VDDD.n1794 VDDD.n1793 209.368
R1172 VDDD.n2362 VDDD.n2361 209.368
R1173 VDDD.n2360 VDDD.n2359 209.368
R1174 VDDD.n2295 VDDD.n2294 209.368
R1175 VDDD.t1856 VDDD 206.45
R1176 VDDD.t341 VDDD.t378 206.45
R1177 VDDD.t201 VDDD.t1931 206.45
R1178 VDDD.t481 VDDD 206.45
R1179 VDDD VDDD.t1060 206.45
R1180 VDDD.t882 VDDD.t832 206.45
R1181 VDDD VDDD.t1764 203.093
R1182 VDDD.t1328 VDDD 203.093
R1183 VDDD.t117 VDDD 203.093
R1184 VDDD VDDD.t971 203.093
R1185 VDDD.t893 VDDD 192.369
R1186 VDDD VDDD.t397 184.63
R1187 VDDD.t1063 VDDD 182.952
R1188 VDDD.t499 VDDD 182.952
R1189 VDDD.t511 VDDD 182.952
R1190 VDDD.t1827 VDDD 182.952
R1191 VDDD.n3171 VDDD 182.952
R1192 VDDD.t505 VDDD 182.952
R1193 VDDD.n910 VDDD 182.952
R1194 VDDD.t1015 VDDD 182.952
R1195 VDDD.t1030 VDDD 182.952
R1196 VDDD.t53 VDDD 182.952
R1197 VDDD VDDD.n2860 182.952
R1198 VDDD.t1144 VDDD 182.952
R1199 VDDD.t1047 VDDD 182.952
R1200 VDDD.t1755 VDDD 182.952
R1201 VDDD.t1165 VDDD 182.952
R1202 VDDD.n2293 VDDD 182.952
R1203 VDDD.t47 VDDD 182.952
R1204 VDDD.t561 VDDD.t1866 181.273
R1205 VDDD.t1486 VDDD.t1918 181.273
R1206 VDDD.t1864 VDDD.t13 181.273
R1207 VDDD.t871 VDDD.t1490 181.273
R1208 VDDD.t1565 VDDD.t253 181.273
R1209 VDDD.t1287 VDDD.t1476 181.273
R1210 VDDD.t1558 VDDD.t670 181.273
R1211 VDDD.t1666 VDDD.t9 181.273
R1212 VDDD.t593 VDDD.t1676 181.273
R1213 VDDD.t1385 VDDD.t337 181.273
R1214 VDDD.t305 VDDD.t1107 181.273
R1215 VDDD.t1344 VDDD.t399 181.273
R1216 VDDD.t549 VDDD.t319 181.273
R1217 VDDD.t1664 VDDD.t613 181.273
R1218 VDDD.t1387 VDDD.t395 181.273
R1219 VDDD.t1278 VDDD.t293 181.273
R1220 VDDD VDDD.n268 179.595
R1221 VDDD VDDD.n3099 179.595
R1222 VDDD VDDD.n909 179.595
R1223 VDDD.t241 VDDD 179.595
R1224 VDDD.n1155 VDDD 179.595
R1225 VDDD VDDD.n1794 179.595
R1226 VDDD.n2683 VDDD 179.595
R1227 VDDD.n2493 VDDD 179.595
R1228 VDDD.n2292 VDDD 179.595
R1229 VDDD.t255 VDDD.t1419 176.238
R1230 VDDD.t1875 VDDD.t325 176.238
R1231 VDDD.t1672 VDDD.t602 176.238
R1232 VDDD VDDD.t231 172.881
R1233 VDDD.t935 VDDD.t493 171.202
R1234 VDDD.t493 VDDD.t898 171.202
R1235 VDDD.t1006 VDDD.t115 171.202
R1236 VDDD.t250 VDDD.t1006 171.202
R1237 VDDD.t1215 VDDD.t1044 171.202
R1238 VDDD.t1322 VDDD.t1055 171.202
R1239 VDDD.t1567 VDDD.t1836 171.202
R1240 VDDD.t1310 VDDD.t994 171.202
R1241 VDDD.t1605 VDDD.t1739 171.202
R1242 VDDD.t1269 VDDD.t1133 171.202
R1243 VDDD.t704 VDDD.t1817 171.202
R1244 VDDD VDDD.t1446 169.524
R1245 VDDD.n617 VDDD.n579 169.398
R1246 VDDD.n800 VDDD.n787 169.398
R1247 VDDD.t878 VDDD.t261 167.845
R1248 VDDD.t1969 VDDD.t71 167.845
R1249 VDDD.t1862 VDDD.t1658 167.845
R1250 VDDD.t389 VDDD.t1704 167.845
R1251 VDDD.t88 VDDD.t1372 166.167
R1252 VDDD.t824 VDDD.t87 166.167
R1253 VDDD.t581 VDDD.t1942 166.167
R1254 VDDD.t1229 VDDD.t418 166.167
R1255 VDDD.t1273 VDDD.t845 166.167
R1256 VDDD.t1532 VDDD.t1622 166.167
R1257 VDDD.t1099 VDDD.t960 166.167
R1258 VDDD.t877 VDDD.t847 166.167
R1259 VDDD.t369 VDDD.t700 166.167
R1260 VDDD.t1901 VDDD.t1701 166.167
R1261 VDDD.t583 VDDD.t1230 166.167
R1262 VDDD.t1879 VDDD.t1604 166.167
R1263 VDDD.t1896 VDDD.t1940 166.167
R1264 VDDD.t685 VDDD.t684 166.167
R1265 VDDD.t1933 VDDD.t617 166.167
R1266 VDDD.t1712 VDDD.t1724 166.167
R1267 VDDD.t1682 VDDD.t1324 166.167
R1268 VDDD.t1425 VDDD.t110 166.167
R1269 VDDD.t1428 VDDD.t539 166.167
R1270 VDDD.t406 VDDD.t862 166.167
R1271 VDDD.t1355 VDDD.t1459 166.167
R1272 VDDD.t345 VDDD.t1458 166.167
R1273 VDDD.t601 VDDD.t1332 166.167
R1274 VDDD.t867 VDDD.t788 166.167
R1275 VDDD.t163 VDDD.t1466 166.167
R1276 VDDD.t945 VDDD.t1625 166.167
R1277 VDDD.t1432 VDDD.t1735 166.167
R1278 VDDD.t1893 VDDD.t168 166.167
R1279 VDDD.t1943 VDDD.t541 166.167
R1280 VDDD.t1326 VDDD.t554 166.167
R1281 VDDD.t1484 VDDD.t734 166.167
R1282 VDDD.t223 VDDD.t735 166.167
R1283 VDDD.t1439 VDDD.t1702 164.488
R1284 VDDD VDDD.t1581 164.488
R1285 VDDD.t1207 VDDD.t1362 164.488
R1286 VDDD.t698 VDDD.t1822 164.488
R1287 VDDD.t243 VDDD.t219 164.488
R1288 VDDD.t1722 VDDD.t989 164.488
R1289 VDDD.t678 VDDD.t1591 162.81
R1290 VDDD.t674 VDDD.t1510 162.81
R1291 VDDD.t1868 VDDD.t94 162.81
R1292 VDDD.t950 VDDD.t656 162.81
R1293 VDDD.t1205 VDDD.t644 162.81
R1294 VDDD.t811 VDDD.t1259 162.81
R1295 VDDD.t929 VDDD.t668 162.81
R1296 VDDD.t1426 VDDD.t1680 162.81
R1297 VDDD.t231 VDDD.t307 162.81
R1298 VDDD.t428 VDDD.t335 162.81
R1299 VDDD.t383 VDDD.t303 162.81
R1300 VDDD.t808 VDDD.t331 162.81
R1301 VDDD.t753 VDDD 162.81
R1302 VDDD.t609 VDDD.t1300 161.131
R1303 VDDD VDDD.t297 161.131
R1304 VDDD.t287 VDDD 159.452
R1305 VDDD.t1195 VDDD.t83 154.417
R1306 VDDD.t886 VDDD.t173 154.417
R1307 VDDD.t691 VDDD.t178 154.417
R1308 VDDD.t1482 VDDD.t1189 154.417
R1309 VDDD.t919 VDDD.t877 154.417
R1310 VDDD.t817 VDDD.t1101 154.417
R1311 VDDD.t154 VDDD.t1712 154.417
R1312 VDDD.t844 VDDD.t1949 154.417
R1313 VDDD.t1419 VDDD.t1209 154.417
R1314 VDDD.t277 VDDD.t255 154.417
R1315 VDDD.t1517 VDDD.t591 154.417
R1316 VDDD.t915 VDDD.t1915 154.417
R1317 VDDD.t412 VDDD.t701 154.417
R1318 VDDD.t957 VDDD.t412 154.417
R1319 VDDD.t1435 VDDD.t1875 154.417
R1320 VDDD.t325 VDDD.t391 154.417
R1321 VDDD.t599 VDDD.t786 154.417
R1322 VDDD.t1194 VDDD.t727 154.417
R1323 VDDD.t868 VDDD.t252 154.417
R1324 VDDD.t252 VDDD.t449 154.417
R1325 VDDD.t1168 VDDD.t481 154.417
R1326 VDDD.t830 VDDD.t954 154.417
R1327 VDDD.t954 VDDD.t1421 154.417
R1328 VDDD.t1747 VDDD.t523 154.417
R1329 VDDD.t906 VDDD.t345 154.417
R1330 VDDD.t1332 VDDD.t1729 154.417
R1331 VDDD.t1450 VDDD.t268 154.417
R1332 VDDD.t268 VDDD.t1733 154.417
R1333 VDDD.t602 VDDD.t749 154.417
R1334 VDDD.t265 VDDD.t1672 154.417
R1335 VDDD.t77 VDDD.t1318 154.417
R1336 VDDD.t453 VDDD.t1393 154.417
R1337 VDDD.t33 VDDD.t1204 154.417
R1338 VDDD.t1629 VDDD.t33 154.417
R1339 VDDD.t1127 VDDD.t1744 154.417
R1340 VDDD.t912 VDDD.t1943 154.417
R1341 VDDD.t801 VDDD.t778 154.417
R1342 VDDD.t61 VDDD.t1326 154.417
R1343 VDDD.t1727 VDDD.t1484 154.417
R1344 VDDD.t682 VDDD.t1402 151.06
R1345 VDDD.t206 VDDD.t225 151.06
R1346 VDDD.t92 VDDD.t607 146.025
R1347 VDDD.t693 VDDD.t837 146.025
R1348 VDDD.t1324 VDDD 146.025
R1349 VDDD.t339 VDDD.t1426 146.025
R1350 VDDD.t281 VDDD.t428 146.025
R1351 VDDD.t1509 VDDD.t1368 144.346
R1352 VDDD.t885 VDDD.t1439 144.346
R1353 VDDD.t200 VDDD.t1261 144.346
R1354 VDDD.t177 VDDD.t139 144.346
R1355 VDDD.t517 VDDD.t950 144.346
R1356 VDDD.t21 VDDD.t37 144.346
R1357 VDDD.t1247 VDDD.t21 144.346
R1358 VDDD.t23 VDDD.t1247 144.346
R1359 VDDD.t459 VDDD.t23 144.346
R1360 VDDD.t1601 VDDD.t125 144.346
R1361 VDDD.t1597 VDDD.t1601 144.346
R1362 VDDD.t127 VDDD.t1597 144.346
R1363 VDDD.t461 VDDD.t131 144.346
R1364 VDDD.t821 VDDD.t457 144.346
R1365 VDDD.t1178 VDDD.t133 144.346
R1366 VDDD.t606 VDDD.t1100 144.346
R1367 VDDD.t1621 VDDD.t1533 144.346
R1368 VDDD.t1362 VDDD.t763 144.346
R1369 VDDD.t1552 VDDD.t723 144.346
R1370 VDDD.t1560 VDDD.t1552 144.346
R1371 VDDD.t700 VDDD.t807 144.346
R1372 VDDD.t1701 VDDD.t371 144.346
R1373 VDDD.t436 VDDD.t1530 144.346
R1374 VDDD.t1526 VDDD.t436 144.346
R1375 VDDD.t1409 VDDD.t1528 144.346
R1376 VDDD.t219 VDDD.t1102 144.346
R1377 VDDD.t1603 VDDD.t442 144.346
R1378 VDDD.t425 VDDD.t726 144.346
R1379 VDDD.t1496 VDDD.t1554 144.346
R1380 VDDD.t965 VDDD.t237 144.346
R1381 VDDD.t237 VDDD.t1500 144.346
R1382 VDDD.t181 VDDD.t179 144.346
R1383 VDDD.t183 VDDD.t235 144.346
R1384 VDDD.t843 VDDD.t1682 144.346
R1385 VDDD.t916 VDDD.t413 144.346
R1386 VDDD.t91 VDDD.t160 144.346
R1387 VDDD.t111 VDDD.t227 144.346
R1388 VDDD.t710 VDDD.t908 144.346
R1389 VDDD.t766 VDDD.t354 144.346
R1390 VDDD.t764 VDDD.t766 144.346
R1391 VDDD.t1607 VDDD.t764 144.346
R1392 VDDD.t348 VDDD.t1609 144.346
R1393 VDDD.t650 VDDD.t646 144.346
R1394 VDDD.t652 VDDD.t648 144.346
R1395 VDDD.t27 VDDD.t25 144.346
R1396 VDDD.t1188 VDDD.t866 144.346
R1397 VDDD.t1719 VDDD.t1373 144.346
R1398 VDDD.t454 VDDD.t1928 144.346
R1399 VDDD.t167 VDDD.t405 144.346
R1400 VDDD.t1891 VDDD.t779 144.346
R1401 VDDD.t553 VDDD.t1327 144.346
R1402 VDDD.t735 VDDD.t1880 144.346
R1403 VDDD.t131 VDDD.t819 142.668
R1404 VDDD.t1257 VDDD.t747 142.668
R1405 VDDD.t1271 VDDD.t1398 142.668
R1406 VDDD.t416 VDDD.t1879 142.668
R1407 VDDD.t863 VDDD.t909 142.668
R1408 VDDD.t862 VDDD.t381 142.668
R1409 VDDD.t1977 VDDD.t350 142.668
R1410 VDDD.t788 VDDD.t941 142.668
R1411 VDDD.t1626 VDDD.t1374 142.668
R1412 VDDD.t1625 VDDD.t666 142.668
R1413 VDDD.t1731 VDDD.t1893 142.668
R1414 VDDD.n3463 VDDD.n370 141.531
R1415 VDDD.t563 VDDD.t565 140.989
R1416 VDDD.t1866 VDDD.t1365 140.989
R1417 VDDD.t1368 VDDD.t561 140.989
R1418 VDDD.t135 VDDD.t1454 140.989
R1419 VDDD.t45 VDDD.t961 140.989
R1420 VDDD.t607 VDDD.t609 140.989
R1421 VDDD.t1300 VDDD.t887 140.989
R1422 VDDD.t1581 VDDD.t96 140.989
R1423 VDDD.t1336 VDDD.t935 140.989
R1424 VDDD.t898 VDDD.t896 140.989
R1425 VDDD.t471 VDDD.t1470 140.989
R1426 VDDD.t689 VDDD.t761 140.989
R1427 VDDD.t1652 VDDD.t1654 140.989
R1428 VDDD.t119 VDDD.t1864 140.989
R1429 VDDD.t13 VDDD.t200 140.989
R1430 VDDD.t891 VDDD.t140 140.989
R1431 VDDD.t1274 VDDD.t529 140.989
R1432 VDDD.t1615 VDDD.t1613 140.989
R1433 VDDD.t115 VDDD.t117 140.989
R1434 VDDD.t175 VDDD.t250 140.989
R1435 VDDD.t248 VDDD.t606 140.989
R1436 VDDD.t1533 VDDD.t1217 140.989
R1437 VDDD.t1219 VDDD.t1215 140.989
R1438 VDDD.t1963 VDDD.t1359 140.989
R1439 VDDD.t65 VDDD.t1691 140.989
R1440 VDDD.t473 VDDD.t209 140.989
R1441 VDDD.t1544 VDDD.t1550 140.989
R1442 VDDD.t1550 VDDD.t1546 140.989
R1443 VDDD.t253 VDDD.t438 140.989
R1444 VDDD.t1563 VDDD.t1567 140.989
R1445 VDDD.t1906 VDDD.t1577 140.989
R1446 VDDD.t1403 VDDD.t717 140.989
R1447 VDDD.t719 VDDD.t1405 140.989
R1448 VDDD.t776 VDDD.t1560 140.989
R1449 VDDD.t604 VDDD.t287 140.989
R1450 VDDD.t1967 VDDD.t698 140.989
R1451 VDDD.t807 VDDD.t419 140.989
R1452 VDDD.t1227 VDDD.t426 140.989
R1453 VDDD.t372 VDDD.t839 140.989
R1454 VDDD.t1289 VDDD.t1310 140.989
R1455 VDDD.t1476 VDDD.t356 140.989
R1456 VDDD.t371 VDDD.t1287 140.989
R1457 VDDD.t1442 VDDD.t423 140.989
R1458 VDDD.t421 VDDD.t1442 140.989
R1459 VDDD.t927 VDDD.t1199 140.989
R1460 VDDD.t385 VDDD.t1409 140.989
R1461 VDDD.t1899 VDDD.t385 140.989
R1462 VDDD.t1965 VDDD.t112 140.989
R1463 VDDD.t440 VDDD.t799 140.989
R1464 VDDD.t1886 VDDD.t1603 140.989
R1465 VDDD.t451 VDDD.t259 140.989
R1466 VDDD.t9 VDDD.t451 140.989
R1467 VDDD.t1523 VDDD.t103 140.989
R1468 VDDD.t1534 VDDD.t1933 140.989
R1469 VDDD.t1870 VDDD.t17 140.989
R1470 VDDD.t726 VDDD.t445 140.989
R1471 VDDD.t780 VDDD.t1722 140.989
R1472 VDDD.t1678 VDDD.t623 140.989
R1473 VDDD.t623 VDDD.t828 140.989
R1474 VDDD.t1314 VDDD 140.989
R1475 VDDD.t337 VDDD.t654 140.989
R1476 VDDD.t1571 VDDD.t1569 140.989
R1477 VDDD.t196 VDDD.t1571 140.989
R1478 VDDD.t192 VDDD.t148 140.989
R1479 VDDD.t1249 VDDD.t152 140.989
R1480 VDDD.t146 VDDD.t1249 140.989
R1481 VDDD.t1107 VDDD.t843 140.989
R1482 VDDD.t1641 VDDD.t305 140.989
R1483 VDDD.t1105 VDDD.t1103 140.989
R1484 VDDD.t1292 VDDD.t1929 140.989
R1485 VDDD.t378 VDDD.t376 140.989
R1486 VDDD.t257 VDDD.t341 140.989
R1487 VDDD.t285 VDDD.t1349 140.989
R1488 VDDD.t205 VDDD.t1394 140.989
R1489 VDDD.t361 VDDD.t1913 140.989
R1490 VDDD.t1235 VDDD.t1233 140.989
R1491 VDDD.t1263 VDDD.t201 140.989
R1492 VDDD.t1931 VDDD.t289 140.989
R1493 VDDD.t559 VDDD.t393 140.989
R1494 VDDD.t1231 VDDD.t597 140.989
R1495 VDDD.t5 VDDD.t1573 140.989
R1496 VDDD.t1221 VDDD.t207 140.989
R1497 VDDD.t539 VDDD.t1291 140.989
R1498 VDDD.t921 VDDD.t263 140.989
R1499 VDDD.t694 VDDD.t111 140.989
R1500 VDDD.t696 VDDD.t67 140.989
R1501 VDDD.t904 VDDD.t708 140.989
R1502 VDDD.t949 VDDD.t1971 140.989
R1503 VDDD.t261 VDDD.t589 140.989
R1504 VDDD.t101 VDDD.t1969 140.989
R1505 VDDD.t71 VDDD.t69 140.989
R1506 VDDD.t399 VDDD.t463 140.989
R1507 VDDD.t612 VDDD.t1344 140.989
R1508 VDDD.t577 VDDD.t1456 140.989
R1509 VDDD.t1538 VDDD.t1468 140.989
R1510 VDDD.t1633 VDDD.t1186 140.989
R1511 VDDD.t866 VDDD.t1182 140.989
R1512 VDDD.t401 VDDD.t1211 140.989
R1513 VDDD.t1211 VDDD.t549 140.989
R1514 VDDD.t902 VDDD.t1627 140.989
R1515 VDDD.t1646 VDDD.t1717 140.989
R1516 VDDD.t267 VDDD.t387 140.989
R1517 VDDD.t1658 VDDD.t1872 140.989
R1518 VDDD.t408 VDDD.t389 140.989
R1519 VDDD.t1704 VDDD.t1269 140.989
R1520 VDDD.t1411 VDDD.t443 140.989
R1521 VDDD.t832 VDDD.t374 140.989
R1522 VDDD.t317 VDDD.t882 140.989
R1523 VDDD.t1239 VDDD.t1662 140.989
R1524 VDDD.t1203 VDDD.t757 140.989
R1525 VDDD.t575 VDDD.t1391 140.989
R1526 VDDD.t613 VDDD.t895 140.989
R1527 VDDD.t895 VDDD.t1670 140.989
R1528 VDDD.t662 VDDD.t167 140.989
R1529 VDDD.t1894 VDDD.t1347 140.989
R1530 VDDD.t579 VDDD.t108 140.989
R1531 VDDD.t39 VDDD.t825 140.989
R1532 VDDD.t395 VDDD.t89 140.989
R1533 VDDD.t779 VDDD.t1387 140.989
R1534 VDDD.t1448 VDDD.t1688 140.989
R1535 VDDD.t631 VDDD.t555 140.989
R1536 VDDD.t1327 VDDD.t1278 140.989
R1537 VDDD.t293 VDDD.t1302 140.989
R1538 VDDD.t1880 VDDD.t702 140.989
R1539 VDDD.t297 VDDD.t229 140.989
R1540 VDDD.t751 VDDD.t704 140.989
R1541 VDDD.t239 VDDD.t1486 139.311
R1542 VDDD VDDD.t455 139.311
R1543 VDDD.t1490 VDDD.t1201 139.311
R1544 VDDD.t670 VDDD.t931 139.311
R1545 VDDD.t1604 VDDD.t1897 139.311
R1546 VDDD.t708 VDDD.t830 139.311
R1547 VDDD.t1464 VDDD.t867 139.311
R1548 VDDD.t1717 VDDD.t1450 139.311
R1549 VDDD.t168 VDDD.t1433 139.311
R1550 VDDD.t677 VDDD.t759 137.633
R1551 VDDD.t782 VDDD.t1961 137.633
R1552 VDDD.t947 VDDD.t1124 137.633
R1553 VDDD.t1521 VDDD.t884 137.633
R1554 VDDD.t1066 VDDD.t447 137.633
R1555 VDDD.t1830 VDDD.t1276 137.633
R1556 VDDD.t467 VDDD.t791 135.954
R1557 VDDD.t1415 VDDD.t635 135.954
R1558 VDDD VDDD.t1423 135.954
R1559 VDDD VDDD.t1334 134.276
R1560 VDDD.t688 VDDD.t1176 134.276
R1561 VDDD.t213 VDDD.t810 134.276
R1562 VDDD.t1609 VDDD 134.276
R1563 VDDD.t646 VDDD.t1686 134.276
R1564 VDDD.n3646 VDDD.t86 132.597
R1565 VDDD.n3645 VDDD.t3 132.597
R1566 VDDD.t1243 VDDD.t835 132.597
R1567 VDDD.n3397 VDDD.t84 132.597
R1568 VDDD.t1660 VDDD.t557 132.597
R1569 VDDD.t1554 VDDD 132.597
R1570 VDDD.t1648 VDDD.t321 132.597
R1571 VDDD.t313 VDDD.t161 132.597
R1572 VDDD.n1937 VDDD.t2076 131.529
R1573 VDDD.t1585 VDDD.t1874 130.919
R1574 VDDD.t819 VDDD.t75 130.919
R1575 VDDD.t881 VDDD.t1255 130.919
R1576 VDDD.t1690 VDDD.t1639 130.919
R1577 VDDD.t411 VDDD.t672 130.919
R1578 VDDD.t1467 VDDD.t106 130.919
R1579 VDDD.t1926 VDDD.t4 130.919
R1580 VDDD.t768 VDDD.t732 130.919
R1581 VDDD.t1460 VDDD.t31 130.919
R1582 VDDD.t1298 VDDD 130.919
R1583 VDDD.n2562 VDDD.t2044 129.344
R1584 VDDD.n3408 VDDD.t2071 129.344
R1585 VDDD.n1040 VDDD.t2080 129.344
R1586 VDDD.n2901 VDDD.t2046 129.344
R1587 VDDD.n2787 VDDD.t2043 129.344
R1588 VDDD.n1543 VDDD.t2081 129.344
R1589 VDDD.n1543 VDDD.t2004 129.344
R1590 VDDD.n268 VDDD 129.24
R1591 VDDD.t1583 VDDD.t969 129.24
R1592 VDDD.t499 VDDD 129.24
R1593 VDDD.t418 VDDD.t1000 129.24
R1594 VDDD.n3099 VDDD 129.24
R1595 VDDD.t1619 VDDD.t1595 129.24
R1596 VDDD.n810 VDDD 129.24
R1597 VDDD.t715 VDDD.t1899 129.24
R1598 VDDD.n2739 VDDD 129.24
R1599 VDDD.n1794 VDDD 129.24
R1600 VDDD.n2360 VDDD 129.24
R1601 VDDD.n2021 VDDD 129.24
R1602 VDDD.t1761 VDDD.t461 127.562
R1603 VDDD.t585 VDDD.t323 127.562
R1604 VDDD VDDD.t844 127.562
R1605 VDDD.t299 VDDD.t1312 127.562
R1606 VDDD.t301 VDDD.t73 127.562
R1607 VDDD.t1003 VDDD 125.883
R1608 VDDD.t490 VDDD 125.883
R1609 VDDD.n3292 VDDD 125.883
R1610 VDDD.n3397 VDDD 125.883
R1611 VDDD.t1790 VDDD 125.883
R1612 VDDD.n3100 VDDD 125.883
R1613 VDDD.t211 VDDD.t328 125.883
R1614 VDDD.t1548 VDDD.t730 125.883
R1615 VDDD.n3170 VDDD 125.883
R1616 VDDD.t1796 VDDD 125.883
R1617 VDDD.n811 VDDD 125.883
R1618 VDDD.t1953 VDDD.t41 125.883
R1619 VDDD.t188 VDDD.t598 125.883
R1620 VDDD.t1050 VDDD 125.883
R1621 VDDD.t241 VDDD 125.883
R1622 VDDD.t150 VDDD 125.883
R1623 VDDD.t56 VDDD 125.883
R1624 VDDD.n2740 VDDD 125.883
R1625 VDDD.n2860 VDDD 125.883
R1626 VDDD.t746 VDDD.t1296 125.883
R1627 VDDD.t484 VDDD 125.883
R1628 VDDD.n2683 VDDD 125.883
R1629 VDDD.t1223 VDDD.t910 125.883
R1630 VDDD.t997 VDDD 125.883
R1631 VDDD.t571 VDDD.t63 125.883
R1632 VDDD.n2493 VDDD 125.883
R1633 VDDD.t1091 VDDD 125.883
R1634 VDDD.n2294 VDDD 125.883
R1635 VDDD VDDD.n2293 125.883
R1636 VDDD VDDD.n2292 125.883
R1637 VDDD.t827 VDDD.t2 124.206
R1638 VDDD.t1488 VDDD 124.206
R1639 VDDD VDDD.t1251 124.206
R1640 VDDD.t1267 VDDD.t1916 124.206
R1641 VDDD.t1882 VDDD.t247 124.206
R1642 VDDD VDDD.t738 124.206
R1643 VDDD.t933 VDDD.t864 124.206
R1644 VDDD.t1333 VDDD.t35 124.206
R1645 VDDD.t1537 VDDD.t29 124.206
R1646 VDDD.t1945 VDDD.t959 124.206
R1647 VDDD.t1944 VDDD.t1190 124.206
R1648 VDDD.t676 VDDD.t1905 122.526
R1649 VDDD.t403 VDDD.t886 122.526
R1650 VDDD.t1361 VDDD.t1962 122.526
R1651 VDDD.t1189 VDDD.t465 122.526
R1652 VDDD.t839 VDDD 122.526
R1653 VDDD.t222 VDDD.t114 122.526
R1654 VDDD.t1101 VDDD.t79 122.526
R1655 VDDD.t447 VDDD 122.526
R1656 VDDD.t1316 VDDD.t1485 122.526
R1657 VDDD.t1506 VDDD.t1908 122.526
R1658 VDDD.n2088 VDDD.n2085 122.514
R1659 VDDD VDDD.t869 120.849
R1660 VDDD.t105 VDDD.t1253 120.849
R1661 VDDD.t333 VDDD.t1265 120.849
R1662 VDDD.t625 VDDD.t352 120.849
R1663 VDDD.n3156 VDDD.t2024 120.76
R1664 VDDD.n3602 VDDD.t1335 119.608
R1665 VDDD.n319 VDDD.t792 119.608
R1666 VDDD.n3642 VDDD.t166 119.608
R1667 VDDD.n3480 VDDD.t870 119.608
R1668 VDDD.n3493 VDDD.t1919 119.608
R1669 VDDD.n3497 VDDD.t1445 119.608
R1670 VDDD.n215 VDDD.t562 119.608
R1671 VDDD.n3340 VDDD.t1218 119.608
R1672 VDDD.n3332 VDDD.t249 119.608
R1673 VDDD.n3311 VDDD.t1714 119.608
R1674 VDDD.n388 VDDD.t14 119.608
R1675 VDDD.n464 VDDD.t901 119.608
R1676 VDDD.n3183 VDDD.t420 119.608
R1677 VDDD.n644 VDDD.t1566 119.608
R1678 VDDD.n687 VDDD.t1321 119.608
R1679 VDDD.n705 VDDD.t872 119.608
R1680 VDDD.n3268 VDDD.t777 119.608
R1681 VDDD.n757 VDDD.t1288 119.608
R1682 VDDD.n845 VDDD.t544 119.608
R1683 VDDD.n849 VDDD.t1559 119.608
R1684 VDDD.n892 VDDD.t1887 119.608
R1685 VDDD.n905 VDDD.t10 119.608
R1686 VDDD.n928 VDDD.t1934 119.608
R1687 VDDD.n932 VDDD.t446 119.608
R1688 VDDD.n1455 VDDD.t1416 119.608
R1689 VDDD.n1449 VDDD.t594 119.608
R1690 VDDD.n1149 VDDD.t1108 119.608
R1691 VDDD.n1384 VDDD.t1386 119.608
R1692 VDDD.n2814 VDDD.t695 119.608
R1693 VDDD.n2809 VDDD.t540 119.608
R1694 VDDD.n1276 VDDD.t1927 119.608
R1695 VDDD.n1289 VDDD.t1232 119.608
R1696 VDDD.n1309 VDDD.t1395 119.608
R1697 VDDD.n1310 VDDD.t107 119.608
R1698 VDDD.n2873 VDDD.t1972 119.608
R1699 VDDD.n2877 VDDD.t1313 119.608
R1700 VDDD.n1811 VDDD.t626 119.608
R1701 VDDD.n1706 VDDD.t1345 119.608
R1702 VDDD.n2589 VDDD.t1183 119.608
R1703 VDDD.n1575 VDDD.t550 119.608
R1704 VDDD.n2617 VDDD.t388 119.608
R1705 VDDD.n2620 VDDD.t74 119.608
R1706 VDDD.n1903 VDDD.t32 119.608
R1707 VDDD.n2348 VDDD.t758 119.608
R1708 VDDD.n2463 VDDD.t1191 119.608
R1709 VDDD.n2433 VDDD.t1946 119.608
R1710 VDDD.n1672 VDDD.t663 119.608
R1711 VDDD.n1885 VDDD.t614 119.608
R1712 VDDD.n2060 VDDD.t1279 119.608
R1713 VDDD.n2187 VDDD.t703 119.608
R1714 VDDD.n1997 VDDD.t1388 119.608
R1715 VDDD.n33 VDDD.t172 119.608
R1716 VDDD.n510 VDDD.t2005 119.257
R1717 VDDD.t1472 VDDD.t1710 119.171
R1718 VDDD.t619 VDDD.t813 119.171
R1719 VDDD.t858 VDDD.t719 119.171
R1720 VDDD.t1504 VDDD.t1385 119.171
R1721 VDDD.t1338 VDDD 119.171
R1722 VDDD.n236 VDDD.t2002 119.007
R1723 VDDD.n1597 VDDD.t2061 119.007
R1724 VDDD.n578 VDDD.t2103 118.919
R1725 VDDD.n786 VDDD.t2077 118.919
R1726 VDDD.n286 VDDD.t2028 118.853
R1727 VDDD.n497 VDDD.t1988 118.853
R1728 VDDD.n3302 VDDD.t2055 118.853
R1729 VDDD.n3347 VDDD.t1990 118.853
R1730 VDDD.n638 VDDD.t2113 118.853
R1731 VDDD.n806 VDDD.t2105 118.853
R1732 VDDD.n1337 VDDD.t2049 118.853
R1733 VDDD.n1656 VDDD.t2100 118.853
R1734 VDDD VDDD.t165 117.492
R1735 VDDD.t1474 VDDD.t215 117.492
R1736 VDDD VDDD.t900 117.492
R1737 VDDD.t1180 VDDD 117.492
R1738 VDDD.t1225 VDDD.t279 117.492
R1739 VDDD.n3257 VDDD.t2057 117.294
R1740 VDDD.n2957 VDDD.t2095 117.294
R1741 VDDD.n2218 VDDD.t2110 117.294
R1742 VDDD.n2301 VDDD.t2042 117.294
R1743 VDDD.n1345 VDDD.t296 116.341
R1744 VDDD.n1342 VDDD.t1679 116.341
R1745 VDDD.t3 VDDD.t793 115.814
R1746 VDDD VDDD.t440 115.814
R1747 VDDD.t755 VDDD.t642 115.814
R1748 VDDD.t1535 VDDD.t1579 115.814
R1749 VDDD.t1413 VDDD.t1883 115.814
R1750 VDDD.t207 VDDD 115.814
R1751 VDDD.t273 VDDD.t535 115.814
R1752 VDDD.t1715 VDDD.t537 115.814
R1753 VDDD.t860 VDDD 115.814
R1754 VDDD.t1186 VDDD 115.814
R1755 VDDD.t1627 VDDD 115.814
R1756 VDDD VDDD.t806 115.814
R1757 VDDD.t736 VDDD 115.814
R1758 VDDD.n2698 VDDD.t2003 115.109
R1759 VDDD.n256 VDDD.t1984 114.912
R1760 VDDD.t1937 VDDD.t676 112.457
R1761 VDDD.t1693 VDDD.t15 112.457
R1762 VDDD.t156 VDDD.t1922 112.457
R1763 VDDD.t834 VDDD.t789 112.457
R1764 VDDD.t1962 VDDD.t329 112.457
R1765 VDDD.t1859 VDDD.t1227 112.457
R1766 VDDD.t114 VDDD.t1519 112.457
R1767 VDDD.t1417 VDDD.t853 112.457
R1768 VDDD.t875 VDDD.t81 112.457
R1769 VDDD.t19 VDDD.t198 112.457
R1770 VDDD VDDD.t11 110.778
R1771 VDDD.t684 VDDD.t1267 110.778
R1772 VDDD.t1494 VDDD 110.778
R1773 VDDD.t864 VDDD.t1425 110.778
R1774 VDDD.t1758 VDDD.t1509 109.1
R1775 VDDD VDDD.t135 109.1
R1776 VDDD.t889 VDDD 109.1
R1777 VDDD.t761 VDDD 109.1
R1778 VDDD.t1261 VDDD.t1141 109.1
R1779 VDDD.t139 VDDD.t50 109.1
R1780 VDDD VDDD.t891 109.1
R1781 VDDD.t125 VDDD.t1096 109.1
R1782 VDDD VDDD.t1963 109.1
R1783 VDDD VDDD.t1965 109.1
R1784 VDDD VDDD.t367 109.1
R1785 VDDD VDDD.t780 109.1
R1786 VDDD.t1468 VDDD 109.1
R1787 VDDD.t551 VDDD 109.1
R1788 VDDD.t63 VDDD 109.1
R1789 VDDD.t1347 VDDD 109.1
R1790 VDDD.t475 VDDD.t1891 109.1
R1791 VDDD VDDD.t1448 109.1
R1792 VDDD VDDD.t177 107.421
R1793 VDDD.t129 VDDD 107.421
R1794 VDDD.t1330 VDDD.t1635 107.421
R1795 VDDD.t1957 VDDD.t1699 107.421
R1796 VDDD.t1959 VDDD.t190 107.421
R1797 VDDD.n2293 VDDD.n2022 106.559
R1798 VDDD.n2021 VDDD.n2020 106.559
R1799 VDDD VDDD.t1079 105.743
R1800 VDDD VDDD.t1812 105.743
R1801 VDDD VDDD.t1012 105.743
R1802 VDDD.t1949 VDDD.t146 105.743
R1803 VDDD VDDD.t629 105.743
R1804 VDDD.t573 VDDD 105.743
R1805 VDDD.t1085 VDDD 105.743
R1806 VDDD VDDD.t520 105.743
R1807 VDDD.t1775 VDDD 105.743
R1808 VDDD VDDD.t363 105.743
R1809 VDDD VDDD.t1127 105.743
R1810 VDDD VDDD.t1088 105.743
R1811 VDDD VDDD.t1074 105.743
R1812 VDDD VDDD.t1799 105.743
R1813 VDDD.t845 VDDD.t1615 104.064
R1814 VDDD.t1639 VDDD.t123 104.064
R1815 VDDD.t356 VDDD 104.064
R1816 VDDD.t1883 VDDD 104.064
R1817 VDDD.t660 VDDD.t233 104.064
R1818 VDDD.t148 VDDD.t1173 104.064
R1819 VDDD.t1340 VDDD.t1338 104.064
R1820 VDDD.t1446 VDDD.t0 104.064
R1821 VDDD VDDD.t563 102.385
R1822 VDDD.t533 VDDD.t584 102.385
R1823 VDDD.t502 VDDD.t587 102.385
R1824 VDDD.t1654 VDDD 102.385
R1825 VDDD VDDD.t175 102.385
R1826 VDDD.t1492 VDDD.t680 102.385
R1827 VDDD.t545 VDDD.t1587 102.385
R1828 VDDD.t531 VDDD.t1357 102.385
R1829 VDDD.t1400 VDDD.t1888 102.385
R1830 VDDD VDDD.t1607 102.385
R1831 VDDD.t770 VDDD.t27 102.385
R1832 VDDD.t1184 VDDD.t1513 102.385
R1833 VDDD.t1304 VDDD.t664 102.385
R1834 VDDD.n2492 VDDD.t1512 102.385
R1835 VDDD VDDD.t1381 102.385
R1836 VDDD VDDD.t1770 102.385
R1837 VDDD.t1784 VDDD.t1178 100.707
R1838 VDDD.t1674 VDDD.t1266 100.707
R1839 VDDD.t1213 VDDD.t1593 100.707
R1840 VDDD.t235 VDDD.t1377 100.707
R1841 VDDD.t1237 VDDD.t59 100.707
R1842 VDDD.t582 VDDD.t271 100.707
R1843 VDDD.t1668 VDDD.t143 100.707
R1844 VDDD.t823 VDDD.t1369 99.0288
R1845 VDDD.t1973 VDDD.t1371 99.0288
R1846 VDDD.t791 VDDD.t1282 99.0288
R1847 VDDD VDDD.t821 99.0288
R1848 VDDD VDDD.t595 99.0288
R1849 VDDD.t1009 VDDD.t1540 99.0288
R1850 VDDD.t852 VDDD.t1415 99.0288
R1851 VDDD.t1725 VDDD.t965 99.0288
R1852 VDDD VDDD.t1575 99.0288
R1853 VDDD.t1778 VDDD.t612 99.0288
R1854 VDDD.t1843 VDDD.t1901 97.3503
R1855 VDDD.t1911 VDDD.t784 95.6719
R1856 VDDD.t1553 VDDD.t1351 95.6719
R1857 VDDD.t1530 VDDD.t925 95.6719
R1858 VDDD.t569 VDDD.t1498 95.6719
R1859 VDDD VDDD.t917 95.6719
R1860 VDDD.t158 VDDD 95.6719
R1861 VDDD VDDD.t1561 95.6719
R1862 VDDD.n910 VDDD.t7 93.9934
R1863 VDDD.t1929 VDDD.n2739 93.9934
R1864 VDDD.n2740 VDDD.t1235 93.9934
R1865 VDDD.t443 VDDD.n2360 93.9934
R1866 VDDD.n278 VDDD.t344 93.81
R1867 VDDD.n321 VDDD.t468 93.81
R1868 VDDD.n3589 VDDD.t157 93.81
R1869 VDDD.n354 VDDD.t16 93.81
R1870 VDDD.n3487 VDDD.t1511 93.81
R1871 VDDD.n3490 VDDD.t1938 93.81
R1872 VDDD.n219 VDDD.t679 93.81
R1873 VDDD.n3378 VDDD.t748 93.81
R1874 VDDD.n3335 VDDD.t1272 93.81
R1875 VDDD.n3434 VDDD.t849 93.81
R1876 VDDD.n380 VDDD.t95 93.81
R1877 VDDD.n3289 VDDD.t951 93.81
R1878 VDDD.n3131 VDDD.t124 93.81
R1879 VDDD.n708 VDDD.t330 93.81
R1880 VDDD.n713 VDDD.t1206 93.81
R1881 VDDD.n588 VDDD.t1657 93.81
R1882 VDDD.n3219 VDDD.t270 93.81
R1883 VDDD.n763 VDDD.t812 93.81
R1884 VDDD.n850 VDDD.t1520 93.81
R1885 VDDD.n856 VDDD.t930 93.81
R1886 VDDD.n885 VDDD.t145 93.81
R1887 VDDD.n888 VDDD.t714 93.81
R1888 VDDD.n922 VDDD.t122 93.81
R1889 VDDD.n925 VDDD.t1917 93.81
R1890 VDDD.n1332 VDDD.t1910 93.81
R1891 VDDD.n1457 VDDD.t636 93.81
R1892 VDDD.n1375 VDDD.t661 93.81
R1893 VDDD.n1133 VDDD.t1696 93.81
R1894 VDDD.n2807 VDDD.t934 93.81
R1895 VDDD.n2803 VDDD.t1685 93.81
R1896 VDDD.n1272 VDDD.t787 93.81
R1897 VDDD.n1273 VDDD.t600 93.81
R1898 VDDD.n1314 VDDD.t592 93.81
R1899 VDDD.n1525 VDDD.t1518 93.81
R1900 VDDD.n2868 VDDD.t1543 93.81
R1901 VDDD.n2870 VDDD.t1427 93.81
R1902 VDDD.n1818 VDDD.t1424 93.81
R1903 VDDD.n1718 VDDD.t232 93.81
R1904 VDDD.n1590 VDDD.t1408 93.81
R1905 VDDD.n1587 VDDD.t773 93.81
R1906 VDDD.n2611 VDDD.t568 93.81
R1907 VDDD.n2613 VDDD.t429 93.81
R1908 VDDD.n1914 VDDD.t78 93.81
R1909 VDDD.n1915 VDDD.t1319 93.81
R1910 VDDD.n2437 VDDD.t1447 93.81
R1911 VDDD.n2429 VDDD.t1339 93.81
R1912 VDDD.n1667 VDDD.t1295 93.81
R1913 VDDD.n2391 VDDD.t1364 93.81
R1914 VDDD.n2064 VDDD.t809 93.81
R1915 VDDD.n2038 VDDD.t44 93.81
R1916 VDDD.n1967 VDDD.t384 93.81
R1917 VDDD.n28 VDDD.t1624 93.81
R1918 VDDD VDDD.t1508 92.315
R1919 VDDD.t1262 VDDD 92.315
R1920 VDDD VDDD.t187 92.315
R1921 VDDD.t1622 VDDD.t1257 92.315
R1922 VDDD.t1398 VDDD.t1099 92.315
R1923 VDDD.t1353 VDDD.t1656 92.315
R1924 VDDD.t432 VDDD.t1197 92.315
R1925 VDDD.t144 VDDD.t416 92.315
R1926 VDDD.t963 VDDD.t611 92.315
R1927 VDDD.t909 VDDD.t1542 92.315
R1928 VDDD.t941 VDDD.t1407 92.315
R1929 VDDD.t1374 VDDD.t567 92.315
R1930 VDDD.t1294 VDDD.t1731 92.315
R1931 VDDD VDDD.t1890 92.315
R1932 VDDD VDDD.t1583 90.6365
R1933 VDDD VDDD.t640 90.6365
R1934 VDDD.t187 VDDD.t517 90.6365
R1935 VDDD.t1595 VDDD 90.6365
R1936 VDDD.t1444 VDDD.t1920 88.9581
R1937 VDDD VDDD.t1322 88.9581
R1938 VDDD.t873 VDDD.t1320 88.9581
R1939 VDDD.t434 VDDD.t923 88.9581
R1940 VDDD.t1556 VDDD.t543 88.9581
R1941 VDDD.t358 VDDD.t339 88.9581
R1942 VDDD VDDD.t1605 88.9581
R1943 VDDD.t1881 VDDD.t281 88.9581
R1944 VDDD VDDD.t615 88.9581
R1945 VDDD.t1162 VDDD.t1695 87.2797
R1946 VDDD.t283 VDDD.t805 87.2797
R1947 VDDD.t542 VDDD.t291 87.2797
R1948 VDDD.t43 VDDD.t1118 87.2797
R1949 VDDD.t1589 VDDD.t1283 85.6012
R1950 VDDD.t359 VDDD.t1955 85.6012
R1951 VDDD.t742 VDDD.t1478 85.6012
R1952 VDDD.t854 VDDD.t621 85.6012
R1953 VDDD.t315 VDDD.t183 85.6012
R1954 VDDD.t1100 VDDD.t686 83.9228
R1955 VDDD.t1461 VDDD.t1621 83.9228
R1956 VDDD.t721 VDDD.t939 83.9228
R1957 VDDD.t414 VDDD.t967 83.9228
R1958 VDDD.n1795 VDDD.t1975 83.9228
R1959 VDDD.t686 VDDD.t841 82.2443
R1960 VDDD.t744 VDDD.t1461 82.2443
R1961 VDDD.t228 VDDD.t1650 82.2443
R1962 VDDD VDDD.t1192 82.2443
R1963 VDDD.t740 VDDD.t650 82.2443
R1964 VDDD.t25 VDDD 82.2443
R1965 VDDD.t706 VDDD.t311 82.2443
R1966 VDDD.t275 VDDD.t856 82.2443
R1967 VDDD.t1367 VDDD 80.5659
R1968 VDDD.t587 VDDD 80.5659
R1969 VDDD.n3293 VDDD.t1599 80.5659
R1970 VDDD VDDD.t880 80.5659
R1971 VDDD VDDD.t583 80.5659
R1972 VDDD VDDD.t410 80.5659
R1973 VDDD.t595 VDDD.n1482 80.5659
R1974 VDDD.t1383 VDDD.n1101 80.5659
R1975 VDDD.t1389 VDDD.t194 80.5659
R1976 VDDD.t1915 VDDD.t1517 80.5659
R1977 VDDD.t786 VDDD.t1194 80.5659
R1978 VDDD.t1393 VDDD.t77 80.5659
R1979 VDDD.t1381 VDDD.t1153 80.5659
R1980 VDDD.t528 VDDD.t815 78.8874
R1981 VDDD.t1713 VDDD.t1708 78.8874
R1982 VDDD.t680 VDDD.t248 78.8874
R1983 VDDD.t1217 VDDD.t545 78.8874
R1984 VDDD.t327 VDDD.t1637 78.8874
R1985 VDDD.t627 VDDD.t346 78.8874
R1986 VDDD.n3647 VDDD.t1138 77.209
R1987 VDDD.t1283 VDDD.t343 77.209
R1988 VDDD.n3100 VDDD.t1150 77.209
R1989 VDDD.t1909 VDDD.t742 77.209
R1990 VDDD.t1528 VDDD.t1308 75.5305
R1991 VDDD.t397 VDDD.t1162 75.5305
R1992 VDDD.t1118 VDDD.t1241 75.5305
R1993 VDDD.t83 VDDD 73.8521
R1994 VDDD VDDD.t92 73.8521
R1995 VDDD VDDD.t693 73.8521
R1996 VDDD.t178 VDDD 73.8521
R1997 VDDD.t1375 VDDD 73.8521
R1998 VDDD.t1192 VDDD 73.8521
R1999 VDDD.t795 VDDD 73.8521
R2000 VDDD.t142 VDDD.t963 73.8521
R2001 VDDD.n2861 VDDD.t1644 73.8521
R2002 VDDD.t1542 VDDD.t358 73.8521
R2003 VDDD.n2682 VDDD.t551 73.8521
R2004 VDDD.t567 VDDD.t1881 73.8521
R2005 VDDD.n2361 VDDD.t245 73.8521
R2006 VDDD.t778 VDDD 73.8521
R2007 VDDD.t797 VDDD.t1109 73.8521
R2008 VDDD.t841 VDDD.t1532 72.1736
R2009 VDDD.t960 VDDD.t744 72.1736
R2010 VDDD.t1306 VDDD.t1526 72.1736
R2011 VDDD.t430 VDDD.t1306 72.1736
R2012 VDDD.t725 VDDD.t721 70.4952
R2013 VDDD.t1351 VDDD.t725 70.4952
R2014 VDDD.t728 VDDD.t1353 70.4952
R2015 VDDD.t1405 VDDD.t728 70.4952
R2016 VDDD.t967 VDDD.t142 70.4952
R2017 VDDD.t419 VDDD.t1859 68.8168
R2018 VDDD.t1308 VDDD.t430 68.8168
R2019 VDDD.t955 VDDD 68.8168
R2020 VDDD.t1369 VDDD.t526 67.1383
R2021 VDDD.t1440 VDDD.t1973 67.1383
R2022 VDDD.n2861 VDDD.t860 67.1383
R2023 VDDD.t1109 VDDD.t736 67.1383
R2024 VDDD.t815 VDDD.t1273 65.4599
R2025 VDDD.t1939 VDDD.t1674 65.4599
R2026 VDDD.t445 VDDD.t755 65.4599
R2027 VDDD.t535 VDDD.t694 65.4599
R2028 VDDD.t350 VDDD.t627 65.4599
R2029 VDDD.t271 VDDD.t1463 65.4599
R2030 VDDD.t380 VDDD.t1668 65.4599
R2031 VDDD.t541 VDDD 65.4599
R2032 VDDD.t1470 VDDD 63.7814
R2033 VDDD.t343 VDDD.t889 63.7814
R2034 VDDD.t217 VDDD 63.7814
R2035 VDDD.t133 VDDD.n3293 63.7814
R2036 VDDD.t367 VDDD.t1909 63.7814
R2037 VDDD.t806 VDDD.n2492 63.7814
R2038 VDDD.n3602 VDDD.t1582 63.3219
R2039 VDDD.n278 VDDD.t1590 63.3219
R2040 VDDD.n319 VDDD.t216 63.3219
R2041 VDDD.n321 VDDD.t1475 63.3219
R2042 VDDD.n3642 VDDD.t1471 63.3219
R2043 VDDD.n3589 VDDD.t659 63.3219
R2044 VDDD.n354 VDDD.t1481 63.3219
R2045 VDDD.n3480 VDDD.t641 63.3219
R2046 VDDD.n3487 VDDD.t675 63.3219
R2047 VDDD.n3490 VDDD.t1586 63.3219
R2048 VDDD.n3493 VDDD.t1487 63.3219
R2049 VDDD.n3497 VDDD.t1584 63.3219
R2050 VDDD.n219 VDDD.t1592 63.3219
R2051 VDDD.n215 VDDD.t1867 63.3219
R2052 VDDD.n3340 VDDD.t1588 63.3219
R2053 VDDD.n3378 VDDD.t1399 63.3219
R2054 VDDD.n3335 VDDD.t1258 63.3219
R2055 VDDD.n3332 VDDD.t1493 63.3219
R2056 VDDD.n3434 VDDD.t1489 63.3219
R2057 VDDD.n3311 VDDD.t1473 63.3219
R2058 VDDD.n380 VDDD.t1869 63.3219
R2059 VDDD.n388 VDDD.t1865 63.3219
R2060 VDDD.n464 VDDD.t218 63.3219
R2061 VDDD.n3289 VDDD.t657 63.3219
R2062 VDDD.n3183 VDDD.t1228 63.3219
R2063 VDDD.n644 VDDD.t254 63.3219
R2064 VDDD.n3131 VDDD.t731 63.3219
R2065 VDDD.n687 VDDD.t1596 63.3219
R2066 VDDD.n705 VDDD.t1491 63.3219
R2067 VDDD.n708 VDDD.t1256 63.3219
R2068 VDDD.n713 VDDD.t645 63.3219
R2069 VDDD.n588 VDDD.t729 63.3219
R2070 VDDD.n3268 VDDD.t288 63.3219
R2071 VDDD.n3219 VDDD.t1252 63.3219
R2072 VDDD.n763 VDDD.t1260 63.3219
R2073 VDDD.n757 VDDD.t1477 63.3219
R2074 VDDD.n845 VDDD.t1900 63.3219
R2075 VDDD.n849 VDDD.t671 63.3219
R2076 VDDD.n850 VDDD.t673 63.3219
R2077 VDDD.n856 VDDD.t669 63.3219
R2078 VDDD.n885 VDDD.t1675 63.3219
R2079 VDDD.n888 VDDD.t1661 63.3219
R2080 VDDD.n892 VDDD.t260 63.3219
R2081 VDDD.n905 VDDD.t1667 63.3219
R2082 VDDD.n922 VDDD.t1594 63.3219
R2083 VDDD.n925 VDDD.t1254 63.3219
R2084 VDDD.n928 VDDD.t1871 63.3219
R2085 VDDD.n932 VDDD.t643 63.3219
R2086 VDDD.n1332 VDDD.t1479 63.3219
R2087 VDDD.n1455 VDDD.t1226 63.3219
R2088 VDDD.n1457 VDDD.t280 63.3219
R2089 VDDD.n1449 VDDD.t1677 63.3219
R2090 VDDD.n1149 VDDD.t306 63.3219
R2091 VDDD.n1375 VDDD.t316 63.3219
R2092 VDDD.n1384 VDDD.t338 63.3219
R2093 VDDD.n1133 VDDD.t398 63.3219
R2094 VDDD.n2814 VDDD.t274 63.3219
R2095 VDDD.n2809 VDDD.t264 63.3219
R2096 VDDD.n2807 VDDD.t334 63.3219
R2097 VDDD.n2803 VDDD.t1238 63.3219
R2098 VDDD.n1272 VDDD.t392 63.3219
R2099 VDDD.n1273 VDDD.t326 63.3219
R2100 VDDD.n1276 VDDD.t394 63.3219
R2101 VDDD.n1289 VDDD.t290 63.3219
R2102 VDDD.n1309 VDDD.t258 63.3219
R2103 VDDD.n1310 VDDD.t286 63.3219
R2104 VDDD.n1314 VDDD.t256 63.3219
R2105 VDDD.n1525 VDDD.t278 63.3219
R2106 VDDD.n2868 VDDD.t340 63.3219
R2107 VDDD.n2870 VDDD.t1681 63.3219
R2108 VDDD.n2873 VDDD.t300 63.3219
R2109 VDDD.n2877 VDDD.t262 63.3219
R2110 VDDD.n1811 VDDD.t733 63.3219
R2111 VDDD.n1818 VDDD.t310 63.3219
R2112 VDDD.n1706 VDDD.t400 63.3219
R2113 VDDD.n1718 VDDD.t308 63.3219
R2114 VDDD.n1590 VDDD.t272 63.3219
R2115 VDDD.n1587 VDDD.t322 63.3219
R2116 VDDD.n2589 VDDD.t402 63.3219
R2117 VDDD.n1575 VDDD.t320 63.3219
R2118 VDDD.n2611 VDDD.t282 63.3219
R2119 VDDD.n2613 VDDD.t336 63.3219
R2120 VDDD.n2617 VDDD.t302 63.3219
R2121 VDDD.n2620 VDDD.t1659 63.3219
R2122 VDDD.n1914 VDDD.t266 63.3219
R2123 VDDD.n1915 VDDD.t1673 63.3219
R2124 VDDD.n1903 VDDD.t1240 63.3219
R2125 VDDD.n2348 VDDD.t318 63.3219
R2126 VDDD.n2437 VDDD.t276 63.3219
R2127 VDDD.n2463 VDDD.t292 63.3219
R2128 VDDD.n2433 VDDD.t284 63.3219
R2129 VDDD.n2429 VDDD.t312 63.3219
R2130 VDDD.n1667 VDDD.t1669 63.3219
R2131 VDDD.n2391 VDDD.t314 63.3219
R2132 VDDD.n1672 VDDD.t1671 63.3219
R2133 VDDD.n1885 VDDD.t1665 63.3219
R2134 VDDD.n2060 VDDD.t294 63.3219
R2135 VDDD.n2064 VDDD.t332 63.3219
R2136 VDDD.n2038 VDDD.t1242 63.3219
R2137 VDDD.n2187 VDDD.t298 63.3219
R2138 VDDD.n1997 VDDD.t396 63.3219
R2139 VDDD.n1967 VDDD.t304 63.3219
R2140 VDDD.n28 VDDD.t639 63.3219
R2141 VDDD.n33 VDDD.t1397 63.3219
R2142 VDDD VDDD.t581 62.103
R2143 VDDD.t1708 VDDD.t528 62.103
R2144 VDDD.t1710 VDDD.t1713 62.103
R2145 VDDD.t1650 VDDD.t327 62.103
R2146 VDDD.t1637 VDDD.t1565 62.103
R2147 VDDD.t1266 VDDD.t144 62.103
R2148 VDDD.t121 VDDD.t1213 62.103
R2149 VDDD.t1724 VDDD 62.103
R2150 VDDD.t59 VDDD.t1684 62.103
R2151 VDDD.t1458 VDDD 62.103
R2152 VDDD.t346 VDDD.t740 62.103
R2153 VDDD.t1407 VDDD.t582 62.103
R2154 VDDD.t143 VDDD.t1294 62.103
R2155 VDDD VDDD.t1894 62.103
R2156 VDDD.t640 VDDD 60.4245
R2157 VDDD.n1482 VDDD.t955 60.4245
R2158 VDDD.t1500 VDDD.t414 60.4245
R2159 VDDD.t738 VDDD.n1101 60.4245
R2160 VDDD.t194 VDDD.t1631 60.4245
R2161 VDDD.t152 VDDD.t1389 60.4245
R2162 VDDD.n1795 VDDD.t348 60.4245
R2163 VDDD.t1153 VDDD.t1379 60.4245
R2164 VDDD.t887 VDDD.t850 58.7461
R2165 VDDD.t1635 VDDD.t228 58.7461
R2166 VDDD.t1955 VDDD.t365 58.7461
R2167 VDDD.t621 VDDD.t1494 58.7461
R2168 VDDD.t233 VDDD.t315 58.7461
R2169 VDDD.t311 VDDD.t1340 58.7461
R2170 VDDD.t0 VDDD.t275 58.7461
R2171 VDDD.t1903 VDDD.t1758 57.0676
R2172 VDDD.t1141 VDDD.t1935 57.0676
R2173 VDDD.t50 VDDD.t1328 57.0676
R2174 VDDD.t959 VDDD.t283 57.0676
R2175 VDDD.t291 VDDD.t1944 57.0676
R2176 VDDD.t1720 VDDD.t475 57.0676
R2177 VDDD.t1613 VDDD 55.3892
R2178 VDDD.t923 VDDD.t359 55.3892
R2179 VDDD.t654 VDDD.t1082 55.3892
R2180 VDDD.t487 VDDD.t1641 55.3892
R2181 VDDD.t173 VDDD.t674 53.7107
R2182 VDDD.t789 VDDD.t1285 53.7107
R2183 VDDD.t37 VDDD 53.7107
R2184 VDDD.t644 VDDD.t1482 53.7107
R2185 VDDD.t365 VDDD 53.7107
R2186 VDDD.t668 VDDD.t817 53.7107
R2187 VDDD.t1593 VDDD.t685 53.7107
R2188 VDDD.t1697 VDDD.t1417 53.7107
R2189 VDDD VDDD.t854 53.7107
R2190 VDDD.t110 VDDD.t1237 53.7107
R2191 VDDD.t805 VDDD.t875 53.7107
R2192 VDDD.t198 VDDD.t542 53.7107
R2193 VDDD.t969 VDDD.t1444 52.0323
R2194 VDDD.t1920 VDDD.t885 52.0323
R2195 VDDD VDDD.t952 52.0323
R2196 VDDD.t1942 VDDD.t502 52.0323
R2197 VDDD.t529 VDDD 52.0323
R2198 VDDD VDDD.t137 52.0323
R2199 VDDD.t1055 VDDD 52.0323
R2200 VDDD.t1947 VDDD 52.0323
R2201 VDDD.t1320 VDDD.t1619 52.0323
R2202 VDDD.t763 VDDD.t873 52.0323
R2203 VDDD VDDD.t65 52.0323
R2204 VDDD.t1577 VDDD 52.0323
R2205 VDDD VDDD.t1967 52.0323
R2206 VDDD.t1197 VDDD.t434 52.0323
R2207 VDDD.t543 VDDD.t715 52.0323
R2208 VDDD.t1102 VDDD.t1556 52.0323
R2209 VDDD.n909 VDDD.t795 52.0323
R2210 VDDD.t799 VDDD 52.0323
R2211 VDDD.t41 VDDD 52.0323
R2212 VDDD VDDD.t1523 52.0323
R2213 VDDD.t1631 VDDD 52.0323
R2214 VDDD VDDD.t1221 52.0323
R2215 VDDD.t1644 VDDD 52.0323
R2216 VDDD VDDD.t904 52.0323
R2217 VDDD.t589 VDDD.t101 52.0323
R2218 VDDD.t1739 VDDD 52.0323
R2219 VDDD.t1342 VDDD 52.0323
R2220 VDDD VDDD.t1633 52.0323
R2221 VDDD VDDD.t1223 52.0323
R2222 VDDD VDDD.t1646 52.0323
R2223 VDDD.t1872 VDDD.t408 52.0323
R2224 VDDD.t245 VDDD 52.0323
R2225 VDDD VDDD.t579 52.0323
R2226 VDDD VDDD.t631 52.0323
R2227 VDDD VDDD.t797 52.0323
R2228 VDDD.t633 VDDD 50.3539
R2229 VDDD.t850 VDDD 50.3539
R2230 VDDD.t86 VDDD 50.3539
R2231 VDDD.t1480 VDDD.t1693 50.3539
R2232 VDDD.t1922 VDDD.t658 50.3539
R2233 VDDD.t84 VDDD 50.3539
R2234 VDDD VDDD.t585 50.3539
R2235 VDDD.t423 VDDD 50.3539
R2236 VDDD.t611 VDDD.t181 50.3539
R2237 VDDD.t1575 VDDD 50.3539
R2238 VDDD.t1138 VDDD 48.6754
R2239 VDDD VDDD.t1793 48.6754
R2240 VDDD.t1812 VDDD 48.6754
R2241 VDDD.t1656 VDDD.t1403 48.6754
R2242 VDDD.t994 VDDD 48.6754
R2243 VDDD.t925 VDDD.t432 48.6754
R2244 VDDD.t1012 VDDD 48.6754
R2245 VDDD.t1502 VDDD.t569 48.6754
R2246 VDDD VDDD.t1085 48.6754
R2247 VDDD.t1770 VDDD 48.6754
R2248 VDDD.t1848 VDDD 46.997
R2249 VDDD.t1112 VDDD 46.997
R2250 VDDD.t215 VDDD.t467 45.3185
R2251 VDDD.t1924 VDDD.t1911 45.3185
R2252 VDDD.t784 VDDD.t217 45.3185
R2253 VDDD.t1599 VDDD 45.3185
R2254 VDDD.t717 VDDD.t1553 45.3185
R2255 VDDD.t635 VDDD.t1225 45.3185
R2256 VDDD.t1498 VDDD.t1725 45.3185
R2257 VDDD VDDD.t1383 45.3185
R2258 VDDD.t629 VDDD 45.3185
R2259 VDDD VDDD.t573 45.3185
R2260 VDDD.t1459 VDDD.t1778 45.3185
R2261 VDDD.t363 VDDD 45.3185
R2262 VDDD.t1905 VDDD.t403 43.6401
R2263 VDDD.t455 VDDD.t1784 43.6401
R2264 VDDD.t465 VDDD.t1361 43.6401
R2265 VDDD.t79 VDDD.t222 43.6401
R2266 VDDD.t1377 VDDD.t1316 43.6401
R2267 VDDD.t67 VDDD 43.6401
R2268 VDDD.t952 VDDD.t823 41.9616
R2269 VDDD.t15 VDDD.t88 41.9616
R2270 VDDD.t87 VDDD.t156 41.9616
R2271 VDDD.t1371 VDDD.t533 41.9616
R2272 VDDD.t1282 VDDD.t827 41.9616
R2273 VDDD.t1916 VDDD.t105 41.9616
R2274 VDDD.t1676 VDDD.t1009 41.9616
R2275 VDDD.t247 VDDD.t852 41.9616
R2276 VDDD.t1569 VDDD 41.9616
R2277 VDDD.t1265 VDDD.t933 41.9616
R2278 VDDD.t1975 VDDD 41.9616
R2279 VDDD.t29 VDDD.t770 41.9616
R2280 VDDD.n280 VDDD.t1284 41.5552
R2281 VDDD.n280 VDDD.t890 41.5552
R2282 VDDD.n349 VDDD.t1974 41.5552
R2283 VDDD.n349 VDDD.t534 41.5552
R2284 VDDD.n357 VDDD.t953 41.5552
R2285 VDDD.n357 VDDD.t1370 41.5552
R2286 VDDD.n3481 VDDD.t1301 41.5552
R2287 VDDD.n3481 VDDD.t888 41.5552
R2288 VDDD.n3484 VDDD.t1438 41.5552
R2289 VDDD.n3484 VDDD.t760 41.5552
R2290 VDDD.n227 VDDD.t1455 41.5552
R2291 VDDD.n227 VDDD.t136 41.5552
R2292 VDDD.n281 VDDD.t690 41.5552
R2293 VDDD.n281 VDDD.t762 41.5552
R2294 VDDD.n499 VDDD.t141 41.5552
R2295 VDDD.n499 VDDD.t892 41.5552
R2296 VDDD.n3343 VDDD.t546 41.5552
R2297 VDDD.n3343 VDDD.t532 41.5552
R2298 VDDD.n3329 VDDD.t138 41.5552
R2299 VDDD.n3329 VDDD.t681 41.5552
R2300 VDDD.n3297 VDDD.t530 41.5552
R2301 VDDD.n3297 VDDD.t1275 41.5552
R2302 VDDD.n375 VDDD.t1925 41.5552
R2303 VDDD.n375 VDDD.t785 41.5552
R2304 VDDD.n716 VDDD.t186 41.5552
R2305 VDDD.n716 VDDD.t783 41.5552
R2306 VDDD.n664 VDDD.t66 41.5552
R2307 VDDD.n664 VDDD.t1692 41.5552
R2308 VDDD.n722 VDDD.t1360 41.5552
R2309 VDDD.n722 VDDD.t1964 41.5552
R2310 VDDD.n580 VDDD.t1578 41.5552
R2311 VDDD.n580 VDDD.t1907 41.5552
R2312 VDDD.n3174 VDDD.t1968 41.5552
R2313 VDDD.n3174 VDDD.t699 41.5552
R2314 VDDD.n772 VDDD.t1700 41.5552
R2315 VDDD.n772 VDDD.t191 41.5552
R2316 VDDD.n859 VDDD.t221 41.5552
R2317 VDDD.n859 VDDD.t1522 41.5552
R2318 VDDD.n876 VDDD.t800 41.5552
R2319 VDDD.n876 VDDD.t441 41.5552
R2320 VDDD.n875 VDDD.t113 41.5552
R2321 VDDD.n875 VDDD.t1966 41.5552
R2322 VDDD.n881 VDDD.t42 41.5552
R2323 VDDD.n881 VDDD.t1898 41.5552
R2324 VDDD.n913 VDDD.t1524 41.5552
R2325 VDDD.n913 VDDD.t104 41.5552
R2326 VDDD.n919 VDDD.t189 41.5552
R2327 VDDD.n919 VDDD.t683 41.5552
R2328 VDDD.n1333 VDDD.t743 41.5552
R2329 VDDD.n1333 VDDD.t368 41.5552
R2330 VDDD.n1366 VDDD.t570 41.5552
R2331 VDDD.n1366 VDDD.t1726 41.5552
R2332 VDDD.n1339 VDDD.t1723 41.5552
R2333 VDDD.n1339 VDDD.t781 41.5552
R2334 VDDD.n1122 VDDD.t1632 41.5552
R2335 VDDD.n1122 VDDD.t1390 41.5552
R2336 VDDD.n1249 VDDD.t1645 41.5552
R2337 VDDD.n1249 VDDD.t861 41.5552
R2338 VDDD.n2846 VDDD.t1297 41.5552
R2339 VDDD.n2846 VDDD.t226 41.5552
R2340 VDDD.n1258 VDDD.t1222 41.5552
R2341 VDDD.n1258 VDDD.t208 41.5552
R2342 VDDD.n1264 VDDD.t159 41.5552
R2343 VDDD.n1264 VDDD.t574 41.5552
R2344 VDDD.n1267 VDDD.t6 41.5552
R2345 VDDD.n1267 VDDD.t1574 41.5552
R2346 VDDD.n1530 VDDD.t1914 41.5552
R2347 VDDD.n1530 VDDD.t362 41.5552
R2348 VDDD.n1532 VDDD.t918 41.5552
R2349 VDDD.n1532 VDDD.t630 41.5552
R2350 VDDD.n2862 VDDD.t905 41.5552
R2351 VDDD.n2862 VDDD.t709 41.5552
R2352 VDDD.n1825 VDDD.t1539 41.5552
R2353 VDDD.n1825 VDDD.t1469 41.5552
R2354 VDDD.n1732 VDDD.t1457 41.5552
R2355 VDDD.n1732 VDDD.t578 41.5552
R2356 VDDD.n1596 VDDD.t1634 41.5552
R2357 VDDD.n1596 VDDD.t1187 41.5552
R2358 VDDD.n1594 VDDD.t1224 41.5552
R2359 VDDD.n1594 VDDD.t1465 41.5552
R2360 VDDD.n2604 VDDD.t903 41.5552
R2361 VDDD.n2604 VDDD.t1628 41.5552
R2362 VDDD.n2605 VDDD.t1647 41.5552
R2363 VDDD.n2605 VDDD.t1718 41.5552
R2364 VDDD.n1931 VDDD.t1562 41.5552
R2365 VDDD.n1931 VDDD.t364 41.5552
R2366 VDDD.n1946 VDDD.t1392 41.5552
R2367 VDDD.n1946 VDDD.t576 41.5552
R2368 VDDD.n1660 VDDD.t1895 41.5552
R2369 VDDD.n1660 VDDD.t1348 41.5552
R2370 VDDD.n1661 VDDD.t580 41.5552
R2371 VDDD.n1661 VDDD.t109 41.5552
R2372 VDDD.n1640 VDDD.t826 41.5552
R2373 VDDD.n1640 VDDD.t40 41.5552
R2374 VDDD.n2406 VDDD.t1434 41.5552
R2375 VDDD.n2406 VDDD.t64 41.5552
R2376 VDDD.n2087 VDDD.t632 41.5552
R2377 VDDD.n2087 VDDD.t556 41.5552
R2378 VDDD.n2042 VDDD.t798 41.5552
R2379 VDDD.n2042 VDDD.t737 41.5552
R2380 VDDD.n1974 VDDD.t1689 41.5552
R2381 VDDD.n1974 VDDD.t1449 41.5552
R2382 VDDD.n16 VDDD.t99 41.5552
R2383 VDDD.n16 VDDD.t894 41.5552
R2384 VDDD.t179 VDDD.t660 40.2832
R2385 VDDD VDDD.t848 38.6047
R2386 VDDD.t137 VDDD.t1492 38.6047
R2387 VDDD.t1587 VDDD.t531 38.6047
R2388 VDDD.t269 VDDD 38.6047
R2389 VDDD.t1888 VDDD.t1666 38.6047
R2390 VDDD.t1884 VDDD.t1400 38.6047
R2391 VDDD.t1683 VDDD 38.6047
R2392 VDDD.t319 VDDD.t1184 38.6047
R2393 VDDD.t1513 VDDD.t469 38.6047
R2394 VDDD.t803 VDDD.t1304 38.6047
R2395 VDDD.t664 VDDD.t1664 38.6047
R2396 VDDD VDDD.t1180 36.9263
R2397 VDDD.t123 VDDD.t1548 36.9263
R2398 VDDD VDDD.t593 36.9263
R2399 VDDD.t1173 VDDD.t196 36.9263
R2400 VDDD.t1096 VDDD.t459 35.2479
R2401 VDDD.n3556 VDDD.n3555 34.6358
R2402 VDDD.n3086 VDDD.n3085 34.6358
R2403 VDDD.n3035 VDDD.n812 34.6358
R2404 VDDD.n1078 VDDD.n1077 34.6358
R2405 VDDD.n2913 VDDD.n2912 34.6358
R2406 VDDD.n2651 VDDD.n2650 34.6358
R2407 VDDD.n2452 VDDD.n2438 34.6358
R2408 VDDD.n2479 VDDD.n1647 34.6358
R2409 VDDD.n312 VDDD.n276 34.6358
R2410 VDDD.n318 VDDD.n274 34.6358
R2411 VDDD.n314 VDDD.n274 34.6358
R2412 VDDD.n3601 VDDD.n347 34.6358
R2413 VDDD.n3587 VDDD.n352 34.6358
R2414 VDDD.n3588 VDDD.n3587 34.6358
R2415 VDDD.n3591 VDDD.n3588 34.6358
R2416 VDDD.n3551 VDDD.n3550 34.6358
R2417 VDDD.n3547 VDDD.n3488 34.6358
R2418 VDDD.n3542 VDDD.n3541 34.6358
R2419 VDDD.n3371 VDDD.n3370 34.6358
R2420 VDDD.n3377 VDDD.n3376 34.6358
R2421 VDDD.n3384 VDDD.n3383 34.6358
R2422 VDDD.n3390 VDDD.n3389 34.6358
R2423 VDDD.n3425 VDDD.n3309 34.6358
R2424 VDDD.n3137 VDDD.n3136 34.6358
R2425 VDDD.n3128 VDDD.n654 34.6358
R2426 VDDD.n3133 VDDD.n3130 34.6358
R2427 VDDD.n743 VDDD.n742 34.6358
R2428 VDDD.n740 VDDD.n711 34.6358
R2429 VDDD.n736 VDDD.n735 34.6358
R2430 VDDD.n606 VDDD.n605 34.6358
R2431 VDDD.n603 VDDD.n586 34.6358
R2432 VDDD.n3270 VDDD.n570 34.6358
R2433 VDDD.n3043 VDDD.n768 34.6358
R2434 VDDD.n1082 VDDD.n840 34.6358
R2435 VDDD.n1064 VDDD.n1063 34.6358
R2436 VDDD.n1061 VDDD.n854 34.6358
R2437 VDDD.n1057 VDDD.n1056 34.6358
R2438 VDDD.n1054 VDDD.n861 34.6358
R2439 VDDD.n1028 VDDD.n1027 34.6358
R2440 VDDD.n1027 VDDD.n1026 34.6358
R2441 VDDD.n1020 VDDD.n1019 34.6358
R2442 VDDD.n1015 VDDD.n1014 34.6358
R2443 VDDD.n978 VDDD.n977 34.6358
R2444 VDDD.n973 VDDD.n972 34.6358
R2445 VDDD.n967 VDDD.n966 34.6358
R2446 VDDD.n963 VDDD.n929 34.6358
R2447 VDDD.n1500 VDDD.n1499 34.6358
R2448 VDDD.n1505 VDDD.n1329 34.6358
R2449 VDDD.n1505 VDDD.n1504 34.6358
R2450 VDDD.n1418 VDDD.n1362 34.6358
R2451 VDDD.n1435 VDDD.n1343 34.6358
R2452 VDDD.n2987 VDDD.n2986 34.6358
R2453 VDDD.n2830 VDDD.n2810 34.6358
R2454 VDDD.n2834 VDDD.n2833 34.6358
R2455 VDDD.n2840 VDDD.n2839 34.6358
R2456 VDDD.n2845 VDDD.n2844 34.6358
R2457 VDDD.n2772 VDDD.n1270 34.6358
R2458 VDDD.n2776 VDDD.n1270 34.6358
R2459 VDDD.n2763 VDDD.n2762 34.6358
R2460 VDDD.n2738 VDDD.n1295 34.6358
R2461 VDDD.n2725 VDDD.n1312 34.6358
R2462 VDDD.n1556 VDDD.n1527 34.6358
R2463 VDDD.n1556 VDDD.n1555 34.6358
R2464 VDDD.n2931 VDDD.n2866 34.6358
R2465 VDDD.n2927 VDDD.n2926 34.6358
R2466 VDDD.n2923 VDDD.n2871 34.6358
R2467 VDDD.n1857 VDDD.n1856 34.6358
R2468 VDDD.n1610 VDDD.n1593 34.6358
R2469 VDDD.n1614 VDDD.n1593 34.6358
R2470 VDDD.n1620 VDDD.n1619 34.6358
R2471 VDDD.n1625 VDDD.n1624 34.6358
R2472 VDDD.n2681 VDDD.n1572 34.6358
R2473 VDDD.n2669 VDDD.n2609 34.6358
R2474 VDDD.n2665 VDDD.n2664 34.6358
R2475 VDDD.n2661 VDDD.n2614 34.6358
R2476 VDDD.n1954 VDDD.n1927 34.6358
R2477 VDDD.n1954 VDDD.n1953 34.6358
R2478 VDDD.n2344 VDDD.n2343 34.6358
R2479 VDDD.n2359 VDDD.n1889 34.6358
R2480 VDDD.n2413 VDDD.n1663 34.6358
R2481 VDDD.n2409 VDDD.n2405 34.6358
R2482 VDDD.n2405 VDDD.n2404 34.6358
R2483 VDDD.n2398 VDDD.n2397 34.6358
R2484 VDDD.n2393 VDDD.n2390 34.6358
R2485 VDDD.n2364 VDDD.n2362 34.6358
R2486 VDDD.n3781 VDDD.n3780 34.6358
R2487 VDDD.n3776 VDDD.n3775 34.6358
R2488 VDDD.n3757 VDDD.n3756 34.6358
R2489 VDDD.n3757 VDDD.n20 34.6358
R2490 VDDD.n3773 VDDD.n20 34.6358
R2491 VDDD.n3754 VDDD.n29 34.6358
R2492 VDDD.n3748 VDDD.n31 34.6358
R2493 VDDD.n3749 VDDD.n3748 34.6358
R2494 VDDD.n3450 VDDD.n3449 34.3278
R2495 VDDD.n307 VDDD.n306 33.8829
R2496 VDDD.n3366 VDDD.n3365 33.8829
R2497 VDDD.n3395 VDDD.n3330 33.8829
R2498 VDDD.n3430 VDDD.n3305 33.8829
R2499 VDDD.n3038 VDDD.n3037 33.8829
R2500 VDDD.n1494 VDDD.n1334 33.8829
R2501 VDDD.n1853 VDDD.n1817 33.8829
R2502 VDDD.n531 VDDD.n530 33.6462
R2503 VDDD.n1402 VDDD.n1373 33.6462
R2504 VDDD.n1404 VDDD.n1403 33.6462
R2505 VDDD.n1412 VDDD.n1411 33.6462
R2506 VDDD.n1876 VDDD.n1875 33.6462
R2507 VDDD.n1865 VDDD.n1864 33.6462
R2508 VDDD.t900 VDDD 33.5694
R2509 VDDD.t1546 VDDD.t1330 33.5694
R2510 VDDD.t1699 VDDD.t421 33.5694
R2511 VDDD.t190 VDDD.t1957 33.5694
R2512 VDDD.t442 VDDD.t1660 33.5694
R2513 VDDD VDDD.t1496 33.5694
R2514 VDDD.t321 VDDD.t1188 33.5694
R2515 VDDD.t405 VDDD.t313 33.5694
R2516 VDDD.n1356 VDDD.n1346 33.5064
R2517 VDDD.n330 VDDD.n329 33.1299
R2518 VDDD.n1454 VDDD.n1452 33.1299
R2519 VDDD.n2476 VDDD.n2475 33.1299
R2520 VDDD.n2368 VDDD.n2367 33.1299
R2521 VDDD.n1000 VDDD.n999 32.7534
R2522 VDDD.n2600 VDDD.n2597 32.7534
R2523 VDDD.n2678 VDDD.n1573 32.7534
R2524 VDDD.n2456 VDDD.n2455 32.7534
R2525 VDDD.n1022 VDDD.n883 32.377
R2526 VDDD.n2777 VDDD.n2776 32.377
R2527 VDDD.n1555 VDDD.n1554 32.377
R2528 VDDD.n2934 VDDD.n2933 32.377
R2529 VDDD.n2932 VDDD.n2931 32.377
R2530 VDDD.n1616 VDDD.n1615 32.377
R2531 VDDD.n2672 VDDD.n2671 32.377
R2532 VDDD.n2670 VDDD.n2669 32.377
R2533 VDDD.n1953 VDDD.n1952 32.377
R2534 VDDD.n2400 VDDD.n1665 32.377
R2535 VDDD.n3774 VDDD.n3773 32.377
R2536 VDDD.n3031 VDDD.n3030 32.377
R2537 VDDD.n1086 VDDD.n1085 32.377
R2538 VDDD.n992 VDDD.n991 32.377
R2539 VDDD.n2909 VDDD.n2879 32.377
R2540 VDDD.n2647 VDDD.n2622 32.377
R2541 VDDD.n314 VDDD.n313 32.0005
R2542 VDDD.n3543 VDDD.n3542 32.0005
R2543 VDDD.n3140 VDDD.n647 32.0005
R2544 VDDD.n742 VDDD.n741 32.0005
R2545 VDDD.n1063 VDDD.n1062 32.0005
R2546 VDDD.n971 VDDD.n970 32.0005
R2547 VDDD.n1504 VDDD.n1330 32.0005
R2548 VDDD.n2994 VDDD.n2993 32.0005
R2549 VDDD.n2838 VDDD.n2805 32.0005
R2550 VDDD.n2764 VDDD.n2763 32.0005
R2551 VDDD.n2721 VDDD.n1312 32.0005
R2552 VDDD.n2919 VDDD.n2918 32.0005
R2553 VDDD.n2657 VDDD.n2656 32.0005
R2554 VDDD.n2343 VDDD.n2342 32.0005
R2555 VDDD.n3750 VDDD.n3749 32.0005
R2556 VDDD.t1874 VDDD.t1937 31.891
R2557 VDDD.t1176 VDDD.t203 31.891
R2558 VDDD.t329 VDDD.t881 31.891
R2559 VDDD.t1519 VDDD.t411 31.891
R2560 VDDD.t1245 VDDD.t213 31.891
R2561 VDDD VDDD.t547 31.891
R2562 VDDD.n3124 VDDD.n657 31.624
R2563 VDDD.n1805 VDDD.n1684 31.4519
R2564 VDDD.n3427 VDDD.n3426 31.2476
R2565 VDDD.n599 VDDD.n598 31.2476
R2566 VDDD.n837 VDDD.n828 30.8711
R2567 VDDD.n2988 VDDD.n2987 30.8711
R2568 VDDD.n1417 VDDD.n1415 30.7205
R2569 VDDD.n1861 VDDD.n1814 30.7205
R2570 VDDD VDDD.t1488 30.2125
R2571 VDDD.t557 VDDD.t713 30.2125
R2572 VDDD.t7 VDDD 30.2125
R2573 VDDD.t772 VDDD.t1648 30.2125
R2574 VDDD.t161 VDDD.t1363 30.2125
R2575 VDDD.n3568 VDDD.n3567 30.1181
R2576 VDDD.n3147 VDDD.n3146 30.1181
R2577 VDDD.n1012 VDDD.n1011 30.1181
R2578 VDDD.n2917 VDDD.n2916 30.1181
R2579 VDDD.n2591 VDDD.n2590 30.1181
R2580 VDDD.n2655 VDDD.n2654 30.1181
R2581 VDDD.n2464 VDDD.n2462 30.1181
R2582 VDDD.n2469 VDDD.n2468 30.1181
R2583 VDDD.n2388 VDDD.n2387 30.1181
R2584 VDDD.n3744 VDDD.n3743 30.1181
R2585 VDDD.n3530 VDDD.n3529 29.7417
R2586 VDDD.n3370 VDDD.n3341 29.7417
R2587 VDDD.n3372 VDDD.n3338 29.7417
R2588 VDDD.n3385 VDDD.n3333 29.7417
R2589 VDDD.n3391 VDDD.n3390 29.7417
R2590 VDDD.n3082 VDDD.n688 29.7417
R2591 VDDD.n1074 VDDD.n846 29.7417
R2592 VDDD.n907 VDDD.n906 29.7417
R2593 VDDD.n2595 VDDD.n2594 29.7417
R2594 VDDD.n2371 VDDD.n2370 29.7417
R2595 VDDD.n465 VDDD.n463 29.3652
R2596 VDDD.n1800 VDDD.n1687 29.2576
R2597 VDDD.n1396 VDDD.n1395 28.9887
R2598 VDDD.t759 VDDD.t1367 28.5341
R2599 VDDD.t793 VDDD.t834 28.5341
R2600 VDDD VDDD.t976 28.5341
R2601 VDDD.t880 VDDD.t782 28.5341
R2602 VDDD.t1951 VDDD.t211 28.5341
R2603 VDDD VDDD.t927 28.5341
R2604 VDDD.t410 VDDD.t1521 28.5341
R2605 VDDD.t1706 VDDD.t188 28.5341
R2606 VDDD.t853 VDDD.t1413 28.5341
R2607 VDDD.t828 VDDD 28.5341
R2608 VDDD VDDD.t150 28.5341
R2609 VDDD.t1296 VDDD.t1452 28.5341
R2610 VDDD.t1024 VDDD 28.5341
R2611 VDDD.n1345 VDDD.t829 28.4453
R2612 VDDD.n1342 VDDD.t242 28.4453
R2613 VDDD.n3129 VDDD.n3128 27.8593
R2614 VDDD.n595 VDDD.n570 27.8593
R2615 VDDD.n771 VDDD.n768 27.8593
R2616 VDDD.n3027 VDDD.n820 27.8593
R2617 VDDD.n502 VDDD.t22 27.5805
R2618 VDDD.n502 VDDD.t1248 27.5805
R2619 VDDD.n543 VDDD.t24 27.5805
R2620 VDDD.n543 VDDD.t460 27.5805
R2621 VDDD.n514 VDDD.t1598 27.5805
R2622 VDDD.n514 VDDD.t128 27.5805
R2623 VDDD.n512 VDDD.t126 27.5805
R2624 VDDD.n512 VDDD.t1602 27.5805
R2625 VDDD.n517 VDDD.t1181 27.5805
R2626 VDDD.n517 VDDD.t130 27.5805
R2627 VDDD.n520 VDDD.t820 27.5805
R2628 VDDD.n368 VDDD.t822 27.5805
R2629 VDDD.n368 VDDD.t1600 27.5805
R2630 VDDD.n523 VDDD.t462 27.5805
R2631 VDDD.n523 VDDD.t458 27.5805
R2632 VDDD.n369 VDDD.t134 27.5805
R2633 VDDD.n369 VDDD.t1179 27.5805
R2634 VDDD.n817 VDDD.t360 27.5805
R2635 VDDD.n817 VDDD.t435 27.5805
R2636 VDDD.n819 VDDD.t433 27.5805
R2637 VDDD.n819 VDDD.t1531 27.5805
R2638 VDDD.n827 VDDD.t437 27.5805
R2639 VDDD.n827 VDDD.t1527 27.5805
R2640 VDDD.n839 VDDD.t431 27.5805
R2641 VDDD.n839 VDDD.t1529 27.5805
R2642 VDDD.n1372 VDDD.t964 27.5805
R2643 VDDD.n1376 VDDD.t180 27.5805
R2644 VDDD.n1376 VDDD.t234 27.5805
R2645 VDDD.n1379 VDDD.t184 27.5805
R2646 VDDD.n1379 VDDD.t236 27.5805
R2647 VDDD.n1380 VDDD.t1317 27.5805
R2648 VDDD.n1380 VDDD.t1507 27.5805
R2649 VDDD.n1370 VDDD.t1501 27.5805
R2650 VDDD.n1370 VDDD.t968 27.5805
R2651 VDDD.n1409 VDDD.t966 27.5805
R2652 VDDD.n1409 VDDD.t238 27.5805
R2653 VDDD.n1363 VDDD.t1503 27.5805
R2654 VDDD.n1363 VDDD.t1499 27.5805
R2655 VDDD.n1416 VDDD.t1555 27.5805
R2656 VDDD.n1416 VDDD.t1315 27.5805
R2657 VDDD.n1352 VDDD.t1495 27.5805
R2658 VDDD.n1352 VDDD.t1497 27.5805
R2659 VDDD.n1688 VDDD.t1608 27.5805
R2660 VDDD.n1688 VDDD.t1976 27.5805
R2661 VDDD.n1686 VDDD.t349 27.5805
R2662 VDDD.n1686 VDDD.t1610 27.5805
R2663 VDDD.n1685 VDDD.t351 27.5805
R2664 VDDD.n1683 VDDD.t347 27.5805
R2665 VDDD.n1683 VDDD.t651 27.5805
R2666 VDDD.n1808 VDDD.t647 27.5805
R2667 VDDD.n1808 VDDD.t769 27.5805
R2668 VDDD.n1812 VDDD.t653 27.5805
R2669 VDDD.n1812 VDDD.t649 27.5805
R2670 VDDD.n1813 VDDD.t353 27.5805
R2671 VDDD.n1813 VDDD.t36 27.5805
R2672 VDDD.n1816 VDDD.t30 27.5805
R2673 VDDD.n1816 VDDD.t28 27.5805
R2674 VDDD.n1736 VDDD.t767 27.5805
R2675 VDDD.n1736 VDDD.t765 27.5805
R2676 VDDD.n3559 VDDD.n3558 27.4829
R2677 VDDD.n1044 VDDD.n872 27.4829
R2678 VDDD.n1031 VDDD.n879 27.4829
R2679 VDDD.n2992 VDDD.n1127 27.4829
R2680 VDDD.n1608 VDDD.n1607 27.4829
R2681 VDDD.n2407 VDDD.n1663 27.4829
R2682 VDDD.n3786 VDDD.n3785 27.0566
R2683 VDDD.n733 VDDD.n718 27.0566
R2684 VDDD.n1848 VDDD.n1819 27.0566
R2685 VDDD.n2448 VDDD.n2438 27.0566
R2686 VDDD.t1372 VDDD.t824 26.8556
R2687 VDDD VDDD.t127 26.8556
R2688 VDDD VDDD.t295 26.8556
R2689 VDDD.t1394 VDDD.t285 26.8556
R2690 VDDD.t393 VDDD.t1231 26.8556
R2691 VDDD.t309 VDDD 26.8556
R2692 VDDD.t757 VDDD.t1239 26.8556
R2693 VDDD.n3527 VDDD.n3498 26.7859
R2694 VDDD.n3008 VDDD.n3007 26.7299
R2695 VDDD.n3308 VDDD.t1709 26.5955
R2696 VDDD.n3308 VDDD.t1711 26.5955
R2697 VDDD.n520 VDDD.t132 26.5955
R2698 VDDD.n646 VDDD.t1636 26.5955
R2699 VDDD.n646 VDDD.t1651 26.5955
R2700 VDDD.n649 VDDD.t1551 26.5955
R2701 VDDD.n649 VDDD.t1547 26.5955
R2702 VDDD.n650 VDDD.t1549 26.5955
R2703 VDDD.n650 VDDD.t1545 26.5955
R2704 VDDD.n656 VDDD.t212 26.5955
R2705 VDDD.n656 VDDD.t474 26.5955
R2706 VDDD.n653 VDDD.t210 26.5955
R2707 VDDD.n653 VDDD.t1640 26.5955
R2708 VDDD.n585 VDDD.t1352 26.5955
R2709 VDDD.n585 VDDD.t718 26.5955
R2710 VDDD.n589 VDDD.t1404 26.5955
R2711 VDDD.n589 VDDD.t1354 26.5955
R2712 VDDD.n592 VDDD.t1406 26.5955
R2713 VDDD.n592 VDDD.t720 26.5955
R2714 VDDD.n767 VDDD.t424 26.5955
R2715 VDDD.n767 VDDD.t1443 26.5955
R2716 VDDD.n770 VDDD.t422 26.5955
R2717 VDDD.n770 VDDD.t1958 26.5955
R2718 VDDD.n773 VDDD.t1960 26.5955
R2719 VDDD.n773 VDDD.t1200 26.5955
R2720 VDDD.n814 VDDD.t928 26.5955
R2721 VDDD.n814 VDDD.t1956 26.5955
R2722 VDDD.n818 VDDD.t924 26.5955
R2723 VDDD.n818 VDDD.t1198 26.5955
R2724 VDDD.n1372 VDDD.t182 26.5955
R2725 VDDD.n1112 VDDD.t1576 26.5955
R2726 VDDD.n1112 VDDD.t1570 26.5955
R2727 VDDD.n1115 VDDD.t1572 26.5955
R2728 VDDD.n1115 VDDD.t197 26.5955
R2729 VDDD.n1119 VDDD.t149 26.5955
R2730 VDDD.n1119 VDDD.t193 26.5955
R2731 VDDD.n1123 VDDD.t151 26.5955
R2732 VDDD.n1123 VDDD.t195 26.5955
R2733 VDDD.n1126 VDDD.t153 26.5955
R2734 VDDD.n1126 VDDD.t1250 26.5955
R2735 VDDD.n1685 VDDD.t1978 26.5955
R2736 VDDD.n3158 VDDD.n3157 26.3341
R2737 VDDD.n2701 VDDD.n2700 26.3341
R2738 VDDD.n3145 VDDD.n3144 25.977
R2739 VDDD.n604 VDDD.n603 25.977
R2740 VDDD.n2743 VDDD.n2742 25.224
R2741 VDDD.n2735 VDDD.n1296 25.224
R2742 VDDD.n2358 VDDD.n2357 25.224
R2743 VDDD.n3399 VDDD.n3398 25.1912
R2744 VDDD.n3291 VDDD.n371 25.1912
R2745 VDDD.n990 VDDD.n911 25.1912
R2746 VDDD.n1484 VDDD.n1483 25.1912
R2747 VDDD.n3418 VDDD.n3313 25.1912
R2748 VDDD.n469 VDDD.n373 25.1912
R2749 VDDD.n3098 VDDD.n668 25.1912
R2750 VDDD.n1044 VDDD.n1043 25.1912
R2751 VDDD.n1032 VDDD.n1031 25.1912
R2752 VDDD.n3006 VDDD.n1113 25.1912
R2753 VDDD.n2998 VDDD.n1120 25.1912
R2754 VDDD.n2986 VDDD.n1129 25.1912
R2755 VDDD.n2785 VDDD.n2784 25.1912
R2756 VDDD.n1793 VDDD.n1690 25.1912
R2757 VDDD.n1607 VDDD.n1595 25.1912
R2758 VDDD.n3728 VDDD.n38 25.1912
R2759 VDDD.n138 VDDD.n130 25.1912
R2760 VDDD.t1000 VDDD.t1617 25.1772
R2761 VDDD.t642 VDDD.t1535 25.1772
R2762 VDDD.t537 VDDD.t273 25.1772
R2763 VDDD.n1398 VDDD.n1397 24.8691
R2764 VDDD.n1801 VDDD.n1800 24.8691
R2765 VDDD.n3563 VDDD.n3482 24.8476
R2766 VDDD.n3534 VDDD.n3495 24.8476
R2767 VDDD.n460 VDDD.n376 24.8476
R2768 VDDD.n3090 VDDD.n3089 24.8476
R2769 VDDD.n3081 VDDD.n3080 24.8476
R2770 VDDD.n3028 VDDD.n3027 24.8476
R2771 VDDD.n1073 VDDD.n1072 24.8476
R2772 VDDD.n996 VDDD.n908 24.8476
R2773 VDDD.n959 VDDD.n958 24.8476
R2774 VDDD.n2820 VDDD.n2819 24.8476
R2775 VDDD.n2826 VDDD.n2825 24.8476
R2776 VDDD.n3741 VDDD.n34 24.8476
R2777 VDDD.n3046 VDDD.n3045 24.5271
R2778 VDDD.n2741 VDDD.n1293 24.5079
R2779 VDDD.n1547 VDDD.n1533 24.5079
R2780 VDDD.n535 VDDD.n534 24.5077
R2781 VDDD.n3785 VDDD.n15 23.7181
R2782 VDDD.n306 VDDD.n305 23.7181
R2783 VDDD.n3579 VDDD.n269 23.7181
R2784 VDDD.n3446 VDDD.n3445 23.7181
R2785 VDDD.n676 VDDD.n668 23.7181
R2786 VDDD.n1494 VDDD.n1493 23.7181
R2787 VDDD.n1303 VDDD.n1295 23.7181
R2788 VDDD.n1697 VDDD.n1690 23.7181
R2789 VDDD.n1935 VDDD.n1930 23.7181
R2790 VDDD.n1896 VDDD.n1889 23.7181
R2791 VDDD.n2491 VDDD.n1647 23.7181
R2792 VDDD.n1993 VDDD.n1981 23.7181
R2793 VDDD.n2020 VDDD.n1981 23.7181
R2794 VDDD.n3781 VDDD.n15 23.7181
R2795 VDDD.n3715 VDDD.n38 23.7181
R2796 VDDD.n139 VDDD.n138 23.7181
R2797 VDDD.t937 VDDD.t1474 23.4987
R2798 VDDD.t939 VDDD 23.4987
R2799 VDDD VDDD.t1706 23.4987
R2800 VDDD.t1253 VDDD.t1534 23.4987
R2801 VDDD.t279 VDDD.t1430 23.4987
R2802 VDDD.t1452 VDDD 23.4987
R2803 VDDD.t1291 VDDD.t333 23.4987
R2804 VDDD.t1971 VDDD.t710 23.4987
R2805 VDDD.t648 VDDD.t625 23.4987
R2806 VDDD.t387 VDDD.t1719 23.4987
R2807 VDDD VDDD.t1512 23.4987
R2808 VDDD.n327 VDDD.n326 23.3417
R2809 VDDD.n3430 VDDD.n3429 23.3417
R2810 VDDD.n838 VDDD.n837 23.3417
R2811 VDDD.n966 VDDD.n965 23.3417
R2812 VDDD.n1463 VDDD.n1462 23.3417
R2813 VDDD.n2833 VDDD.n2832 23.3417
R2814 VDDD.n2745 VDDD.n2744 23.3417
R2815 VDDD.n2734 VDDD.n2733 23.3417
R2816 VDDD.n1854 VDDD.n1853 23.3417
R2817 VDDD.n1902 VDDD.n1900 23.3417
R2818 VDDD.n2457 VDDD.n2435 23.3417
R2819 VDDD.n2474 VDDD.n2430 23.3417
R2820 VDDD.n2905 VDDD.n2904 23.3088
R2821 VDDD.n2643 VDDD.n2642 23.3088
R2822 VDDD.n606 VDDD.n583 22.9652
R2823 VDDD.n330 VDDD.n270 22.9652
R2824 VDDD.n3551 VDDD.n3485 22.9652
R2825 VDDD.n735 VDDD.n734 22.9652
R2826 VDDD.n1056 VDDD.n1055 22.9652
R2827 VDDD.n979 VDDD.n978 22.9652
R2828 VDDD.n1468 VDDD.n1452 22.9652
R2829 VDDD.n2847 VDDD.n2845 22.9652
R2830 VDDD.n2780 VDDD.n2779 22.9652
R2831 VDDD.n1552 VDDD.n1531 22.9652
R2832 VDDD.n2939 VDDD.n2938 22.9652
R2833 VDDD.n2677 VDDD.n2676 22.9652
R2834 VDDD.n1948 VDDD.n1947 22.9652
R2835 VDDD.n2414 VDDD.n2413 22.9652
R2836 VDDD.n3776 VDDD.n17 22.9652
R2837 VDDD.n3737 VDDD.n3736 22.9652
R2838 VDDD.n1415 VDDD.n1364 22.6748
R2839 VDDD.n1862 VDDD.n1861 22.6748
R2840 VDDD.n3426 VDDD.n3425 22.2123
R2841 VDDD.n1940 VDDD.n1887 22.2123
R2842 VDDD.n3452 VDDD.n3451 22.1096
R2843 VDDD.n3603 VDDD.n3601 22.0807
R2844 VDDD.n3037 VDDD.n3036 21.8358
R2845 VDDD.t813 VDDD.t1472 21.8203
R2846 VDDD VDDD.t1951 21.8203
R2847 VDDD.t723 VDDD.t858 21.8203
R2848 VDDD VDDD.t776 21.8203
R2849 VDDD.t1485 VDDD.t1506 21.8203
R2850 VDDD.t1908 VDDD.t1504 21.8203
R2851 VDDD.t1680 VDDD.t406 21.8203
R2852 VDDD.t335 VDDD.t945 21.8203
R2853 VDDD.n3597 VDDD.n347 21.4593
R2854 VDDD.n3580 VDDD.n3579 21.4593
R2855 VDDD.n3567 VDDD.n3565 21.4593
R2856 VDDD.n3559 VDDD.n3482 21.4593
R2857 VDDD.n3555 VDDD.n3485 21.4593
R2858 VDDD.n3530 VDDD.n3495 21.4593
R2859 VDDD.n3445 VDDD.n3299 21.4593
R2860 VDDD.n3396 VDDD.n3395 21.4593
R2861 VDDD.n462 VDDD.n461 21.4593
R2862 VDDD.n3082 VDDD.n3081 21.4593
R2863 VDDD.n734 VDDD.n733 21.4593
R2864 VDDD.n1074 VDDD.n1073 21.4593
R2865 VDDD.n1055 VDDD.n1054 21.4593
R2866 VDDD.n999 VDDD.n998 21.4593
R2867 VDDD.n992 VDDD.n908 21.4593
R2868 VDDD.n2784 VDDD.n1265 21.4593
R2869 VDDD.n2749 VDDD.n1290 21.4593
R2870 VDDD.n2729 VDDD.n1307 21.4593
R2871 VDDD.n1548 VDDD.n1547 21.4593
R2872 VDDD.n2938 VDDD.n2863 21.4593
R2873 VDDD.n2916 VDDD.n2875 21.4593
R2874 VDDD.n2600 VDDD.n2599 21.4593
R2875 VDDD.n2678 VDDD.n2677 21.4593
R2876 VDDD.n2676 VDDD.n2606 21.4593
R2877 VDDD.n2654 VDDD.n2618 21.4593
R2878 VDDD.n1945 VDDD.n1930 21.4593
R2879 VDDD.n2352 VDDD.n2351 21.4593
R2880 VDDD.n2462 VDDD.n2461 21.4593
R2881 VDDD.n2470 VDDD.n2469 21.4593
R2882 VDDD.n2367 VDDD.n1886 21.4593
R2883 VDDD.n3780 VDDD.n17 21.4593
R2884 VDDD.n3737 VDDD.n34 21.4593
R2885 VDDD.n3270 VDDD.n3269 21.2404
R2886 VDDD.n3452 VDDD.n370 21.2369
R2887 VDDD.n456 VDDD.n455 20.7064
R2888 VDDD.n3158 VDDD.n3155 20.4852
R2889 VDDD.n3245 VDDD.n3172 20.4852
R2890 VDDD.n320 VDDD.n318 20.3299
R2891 VDDD.n3597 VDDD.n3596 20.3299
R2892 VDDD.n3581 VDDD.n3580 20.3299
R2893 VDDD.n3538 VDDD.n3537 20.3299
R2894 VDDD.n3421 VDDD.n3309 20.3299
R2895 VDDD.n465 VDDD.n373 20.3299
R2896 VDDD.n707 VDDD.n706 20.3299
R2897 VDDD.n1068 VDDD.n1067 20.3299
R2898 VDDD.n1456 VDDD.n1329 20.3299
R2899 VDDD.n2762 VDDD.n1277 20.3299
R2900 VDDD.n2726 VDDD.n2725 20.3299
R2901 VDDD.n2918 VDDD.n2917 20.3299
R2902 VDDD.n2656 VDDD.n2655 20.3299
R2903 VDDD.n2344 VDDD.n1904 20.3299
R2904 VDDD.n2468 VDDD.n2432 20.3299
R2905 VDDD.n2464 VDDD.n2432 20.3299
R2906 VDDD.n3744 VDDD.n31 20.3299
R2907 VDDD.t2 VDDD.t688 20.1418
R2908 VDDD.t747 VDDD.t1271 20.1418
R2909 VDDD.t810 VDDD.t1882 20.1418
R2910 VDDD.t352 VDDD.t1333 20.1418
R2911 VDDD.t35 VDDD.t1537 20.1418
R2912 VDDD.t547 VDDD.t902 20.1418
R2913 VDDD.t702 VDDD 20.1418
R2914 VDDD.n1356 VDDD.n1355 19.9534
R2915 VDDD.n1806 VDDD.n1805 19.7491
R2916 VDDD.n455 VDDD.n454 19.633
R2917 VDDD.n2911 VDDD.n2910 19.577
R2918 VDDD.n2649 VDDD.n2648 19.577
R2919 VDDD.n3806 VDDD.n3805 19.2067
R2920 VDDD.n3661 VDDD.n222 19.2067
R2921 VDDD.n1760 VDDD.n1759 19.2067
R2922 VDDD.n2125 VDDD.n2124 19.2067
R2923 VDDD.n2319 VDDD.n2318 19.2067
R2924 VDDD.n95 VDDD.n94 19.2067
R2925 VDDD.n198 VDDD.n197 19.2067
R2926 VDDD.n979 VDDD.n917 19.2005
R2927 VDDD.n2847 VDDD.n1251 19.2005
R2928 VDDD.n3031 VDDD.n816 18.824
R2929 VDDD.n1085 VDDD.n1084 18.824
R2930 VDDD.n1078 VDDD.n842 18.824
R2931 VDDD.n1430 VDDD.n1429 18.824
R2932 VDDD.n1436 VDDD.n1435 18.824
R2933 VDDD.n3244 VDDD.n3242 18.7591
R2934 VDDD.n409 VDDD.n393 18.7474
R2935 VDDD.n308 VDDD.n279 18.4476
R2936 VDDD.n3550 VDDD.n3549 18.4476
R2937 VDDD.n3133 VDDD.n3132 18.4476
R2938 VDDD.n736 VDDD.n715 18.4476
R2939 VDDD.n1057 VDDD.n858 18.4476
R2940 VDDD.n957 VDDD.n956 18.4476
R2941 VDDD.n1498 VDDD.n1497 18.4476
R2942 VDDD.n1395 VDDD.n1382 18.4476
R2943 VDDD.n2824 VDDD.n2813 18.4476
R2944 VDDD.n2926 VDDD.n2925 18.4476
R2945 VDDD.n1849 VDDD.n1848 18.4476
R2946 VDDD.n2664 VDDD.n2663 18.4476
R2947 VDDD.n3595 VDDD.n350 18.0711
R2948 VDDD.n3583 VDDD.n3582 18.0711
R2949 VDDD.n3372 VDDD.n3371 18.0711
R2950 VDDD.n3389 VDDD.n3333 18.0711
R2951 VDDD.n1026 VDDD.n883 18.0711
R2952 VDDD.n977 VDDD.n920 18.0711
R2953 VDDD.n1418 VDDD.n1417 18.0711
R2954 VDDD.n1125 VDDD.n1124 18.0711
R2955 VDDD.n2844 VDDD.n2801 18.0711
R2956 VDDD.n2779 VDDD.n2778 18.0711
R2957 VDDD.n1553 VDDD.n1552 18.0711
R2958 VDDD.n2933 VDDD.n2932 18.0711
R2959 VDDD.n1857 VDDD.n1814 18.0711
R2960 VDDD.n1615 VDDD.n1614 18.0711
R2961 VDDD.n2671 VDDD.n2670 18.0711
R2962 VDDD.n1948 VDDD.n1928 18.0711
R2963 VDDD.n2404 VDDD.n1665 18.0711
R2964 VDDD.n3775 VDDD.n3774 18.0711
R2965 VDDD.n611 VDDD.n610 18.0382
R2966 VDDD.n1469 VDDD.n1468 18.0382
R2967 VDDD.n3736 VDDD.n3735 18.0382
R2968 VDDD.n3450 VDDD.n3296 18.0369
R2969 VDDD.n1219 VDDD.n1218 17.9678
R2970 VDDD.n544 VDDD.n542 17.9537
R2971 VDDD.n1397 VDDD.n1396 17.9205
R2972 VDDD.n3421 VDDD.n3420 17.6946
R2973 VDDD.n1013 VDDD.n1012 17.6946
R2974 VDDD.n2590 VDDD.n1578 17.6946
R2975 VDDD.n2389 VDDD.n2388 17.6946
R2976 VDDD.n245 VDDD.n242 17.612
R2977 VDDD.n420 VDDD.n391 17.612
R2978 VDDD.n3700 VDDD.n3699 17.612
R2979 VDDD.n147 VDDD.n146 17.612
R2980 VDDD.n1408 VDDD.n1368 17.5548
R2981 VDDD.n3827 VDDD.n1 17.3413
R2982 VDDD.n3045 VDDD.n3044 17.3181
R2983 VDDD.n1385 VDDD.n1382 17.0992
R2984 VDDD.t1334 VDDD 16.785
R2985 VDDD.t1764 VDDD.t1652 16.785
R2986 VDDD.t457 VDDD.t1761 16.785
R2987 VDDD.t1190 VDDD.t1945 16.785
R2988 VDDD.n3245 VDDD.n3244 16.7729
R2989 VDDD.n1199 VDDD.n1198 16.6847
R2990 VDDD.n2536 VDDD.n2535 16.6847
R2991 VDDD.n2271 VDDD.n2270 16.6847
R2992 VDDD.n3644 VDDD.n270 16.5652
R2993 VDDD.n1445 VDDD.n1438 16.5652
R2994 VDDD.n279 VDDD.n276 16.1887
R2995 VDDD.n599 VDDD.n591 16.1887
R2996 VDDD.n596 VDDD.n595 16.1887
R2997 VDDD.n1499 VDDD.n1498 16.1887
R2998 VDDD.n1850 VDDD.n1849 16.1887
R2999 VDDD.n2455 VDDD.n2454 16.1887
R3000 VDDD.n2454 VDDD.n2453 16.1887
R3001 VDDD.n2477 VDDD.n2476 16.1887
R3002 VDDD.n2478 VDDD.n2477 16.1887
R3003 VDDD.n3086 VDDD.n684 16.1887
R3004 VDDD.n2165 VDDD.n2163 16.139
R3005 VDDD.n2016 VDDD.n1986 16.139
R3006 VDDD.n3196 VDDD.n3195 15.8683
R3007 VDDD.n3716 VDDD.n3715 15.8683
R3008 VDDD.n3706 VDDD.n48 15.8683
R3009 VDDD.n3138 VDDD.n3137 15.8123
R3010 VDDD.n591 VDDD.n590 15.8123
R3011 VDDD.n1431 VDDD.n1430 15.8123
R3012 VDDD.n1483 VDDD.n1436 15.8123
R3013 VDDD.n1124 VDDD.n1120 15.8123
R3014 VDDD.n2778 VDDD.n2777 15.8123
R3015 VDDD.n2751 VDDD.n1277 15.8123
R3016 VDDD.n2727 VDDD.n2726 15.8123
R3017 VDDD.n1554 VDDD.n1553 15.8123
R3018 VDDD.n1952 VDDD.n1928 15.8123
R3019 VDDD.n2349 VDDD.n1904 15.8123
R3020 VDDD.n1403 VDDD.n1402 15.7262
R3021 VDDD.n1398 VDDD.n1378 15.7262
R3022 VDDD.n3449 VDDD.n3448 15.6579
R3023 VDDD.n3291 VDDD.n3290 15.5335
R3024 VDDD.n1796 VDDD.n1689 15.4774
R3025 VDDD.n1477 VDDD.n1437 15.4029
R3026 VDDD.n3435 VDDD.n3433 15.2745
R3027 VDDD.t328 VDDD.t473 15.1065
R3028 VDDD.t730 VDDD.t1544 15.1065
R3029 VDDD.t1897 VDDD.t1953 15.1065
R3030 VDDD.t598 VDDD.t682 15.1065
R3031 VDDD.t617 VDDD.t1870 15.1065
R3032 VDDD VDDD.t192 15.1065
R3033 VDDD.t225 VDDD.t746 15.1065
R3034 VDDD.t263 VDDD.t1428 15.1065
R3035 VDDD.t1423 VDDD 15.1065
R3036 VDDD.t910 VDDD.t1464 15.1065
R3037 VDDD.t1433 VDDD.t571 15.1065
R3038 VDDD.n3242 VDDD.n3241 15.101
R3039 VDDD.n2556 VDDD.n2555 14.9
R3040 VDDD.n2291 VDDD.n2290 14.9
R3041 VDDD.n816 VDDD.n815 14.6829
R3042 VDDD.n1786 VDDD.n1785 14.6246
R3043 VDDD.n1179 VDDD.n1178 14.5851
R3044 VDDD.n2516 VDDD.n2515 14.5851
R3045 VDDD.n2251 VDDD.n2250 14.5851
R3046 VDDD.n1084 VDDD.n1083 14.3064
R3047 VDDD.n947 VDDD.n944 14.2735
R3048 VDDD.n2859 VDDD.n2858 14.2735
R3049 VDDD.n2894 VDDD.n2893 14.2735
R3050 VDDD.n2635 VDDD.n2634 14.2735
R3051 VDDD.n2491 VDDD.n2490 14.2735
R3052 VDDD.n3706 VDDD.n47 14.2735
R3053 VDDD.n140 VDDD.n139 14.2735
R3054 VDDD.n2188 VDDD.n2186 14.2308
R3055 VDDD.n548 VDDD.n507 14.2027
R3056 VDDD.n2084 VDDD.n2080 14.2027
R3057 VDDD.n2149 VDDD.n2022 13.8955
R3058 VDDD.n3464 VDDD.n3463 13.8514
R3059 VDDD.t75 VDDD.t129 13.4281
R3060 VDDD.t1199 VDDD.n811 13.4281
R3061 VDDD.t376 VDDD.t1292 13.4281
R3062 VDDD.t1349 VDDD.t257 13.4281
R3063 VDDD.t106 VDDD.t205 13.4281
R3064 VDDD.t917 VDDD.t361 13.4281
R3065 VDDD.t1233 VDDD.t1263 13.4281
R3066 VDDD.t289 VDDD.t559 13.4281
R3067 VDDD.t597 VDDD.t1926 13.4281
R3068 VDDD.t1573 VDDD.t158 13.4281
R3069 VDDD.t908 VDDD.t299 13.4281
R3070 VDDD.t1312 VDDD.t878 13.4281
R3071 VDDD.t732 VDDD.t652 13.4281
R3072 VDDD.t1373 VDDD.t301 13.4281
R3073 VDDD.t73 VDDD.t1862 13.4281
R3074 VDDD.t374 VDDD.t1411 13.4281
R3075 VDDD.t1662 VDDD.t317 13.4281
R3076 VDDD.t31 VDDD.t1203 13.4281
R3077 VDDD.t1561 VDDD.t575 13.4281
R3078 VDDD.t554 VDDD.t1804 13.4281
R3079 VDDD.n3398 VDDD.n3396 13.177
R3080 VDDD.n461 VDDD.n460 13.177
R3081 VDDD.n3089 VDDD.n683 13.177
R3082 VDDD.n841 VDDD.n840 13.177
R3083 VDDD.n2746 VDDD.n1290 13.177
R3084 VDDD.n2732 VDDD.n1307 13.177
R3085 VDDD.n2910 VDDD.n2909 13.177
R3086 VDDD.n2648 VDDD.n2647 13.177
R3087 VDDD.n2353 VDDD.n2352 13.177
R3088 VDDD.n2461 VDDD.n2460 13.177
R3089 VDDD.n2471 VDDD.n2470 13.177
R3090 VDDD.n1378 VDDD.n1377 13.1662
R3091 VDDD.n2940 VDDD.n1248 12.9273
R3092 VDDD.n267 VDDD.n266 12.8005
R3093 VDDD.n301 VDDD.n300 12.8005
R3094 VDDD.n3288 VDDD.n479 12.8005
R3095 VDDD.n404 VDDD.n397 12.8005
R3096 VDDD.n3361 VDDD.n3360 12.8005
R3097 VDDD.n3136 VDDD.n651 12.8005
R3098 VDDD.n809 VDDD.n780 12.8005
R3099 VDDD.n3036 VDDD.n3035 12.8005
R3100 VDDD.n2163 VDDD.n2022 12.8005
R3101 VDDD.n2020 VDDD.n1986 12.8005
R3102 VDDD.n256 VDDD.n255 12.4487
R3103 VDDD.n2698 VDDD.n2697 12.4487
R3104 VDDD.n1807 VDDD.n1806 12.4348
R3105 VDDD.n3565 VDDD.n3564 12.424
R3106 VDDD.n3144 VDDD.n647 12.424
R3107 VDDD.n1355 VDDD.n1353 12.424
R3108 VDDD.n2993 VDDD.n2992 12.424
R3109 VDDD.n1481 VDDD.n1438 12.0476
R3110 VDDD.n3009 VDDD.n3008 12.0476
R3111 VDDD.n3091 VDDD.n3090 12.0147
R3112 VDDD.n2819 VDDD.n2818 12.0147
R3113 VDDD.n3010 VDDD.n3009 11.818
R3114 VDDD.t1940 VDDD.t1886 11.7496
R3115 VDDD VDDD.t1314 11.7496
R3116 VDDD.t1209 VDDD.t916 11.7496
R3117 VDDD.t701 VDDD.t915 11.7496
R3118 VDDD.t160 VDDD.t1435 11.7496
R3119 VDDD.t727 VDDD.t868 11.7496
R3120 VDDD.t1421 VDDD.t863 11.7496
R3121 VDDD.t1182 VDDD.t163 11.7496
R3122 VDDD.t1733 VDDD.t1626 11.7496
R3123 VDDD.t749 VDDD.t454 11.7496
R3124 VDDD.t1204 VDDD.t453 11.7496
R3125 VDDD.t1735 VDDD.t662 11.7496
R3126 VDDD.n548 VDDD.n503 11.6711
R3127 VDDD.n609 VDDD.n583 11.6711
R3128 VDDD.n328 VDDD.n327 11.2946
R3129 VDDD.n3140 VDDD.n3139 11.2946
R3130 VDDD.n1087 VDDD.n838 11.2946
R3131 VDDD.n1464 VDDD.n1463 11.2946
R3132 VDDD.n2924 VDDD.n2923 11.2946
R3133 VDDD.n2662 VDDD.n2661 11.2946
R3134 VDDD.n2460 VDDD.n2435 11.2946
R3135 VDDD.n2471 VDDD.n2430 11.2946
R3136 VDDD.n3644 VDDD.n3643 11.1998
R3137 VDDD.n998 VDDD.n997 10.9181
R3138 VDDD.n2599 VDDD.n2598 10.9181
R3139 VDDD.n2363 VDDD.n1886 10.9181
R3140 VDDD.n2089 VDDD.n2088 10.848
R3141 VDDD.n1481 VDDD.n1437 10.5417
R3142 VDDD.n2940 VDDD.n2939 10.5417
R3143 VDDD.n2085 VDDD.n2084 10.5417
R3144 VDDD.n531 VDDD.n518 10.2405
R3145 VDDD.n1404 VDDD.n1371 10.2405
R3146 VDDD.n1367 VDDD.n1364 10.2405
R3147 VDDD.n3124 VDDD.n3123 10.2212
R3148 VDDD.t1918 VDDD.t1585 10.0712
R3149 VDDD.t140 VDDD.t1036 10.0712
R3150 VDDD.t1255 VDDD.t871 10.0712
R3151 VDDD.t209 VDDD.t1690 10.0712
R3152 VDDD.t672 VDDD.t1558 10.0712
R3153 VDDD.t103 VDDD.t986 10.0712
R3154 VDDD.t17 VDDD.t425 10.0712
R3155 VDDD.t413 VDDD.t1467 10.0712
R3156 VDDD.t4 VDDD.t91 10.0712
R3157 VDDD.t227 VDDD.t921 10.0712
R3158 VDDD VDDD.t1977 10.0712
R3159 VDDD.t1686 VDDD.t768 10.0712
R3160 VDDD.t514 VDDD.t1538 10.0712
R3161 VDDD.t1928 VDDD.t1460 10.0712
R3162 VDDD.t108 VDDD.t1121 10.0712
R3163 VDDD.n3429 VDDD.n3428 9.78874
R3164 VDDD.n3029 VDDD.n3028 9.78874
R3165 VDDD.n2780 VDDD.n1265 9.78874
R3166 VDDD.n2744 VDDD.n2743 9.78874
R3167 VDDD.n2735 VDDD.n2734 9.78874
R3168 VDDD.n1548 VDDD.n1531 9.78874
R3169 VDDD.n1947 VDDD.n1945 9.78874
R3170 VDDD.n2357 VDDD.n1900 9.78874
R3171 VDDD.n3810 VDDD.n3809 9.73273
R3172 VDDD.n3811 VDDD.n3810 9.73273
R3173 VDDD.n3815 VDDD.n3814 9.73273
R3174 VDDD.n3816 VDDD.n3815 9.73273
R3175 VDDD.n3816 VDDD.n3 9.73273
R3176 VDDD.n3820 VDDD.n3 9.73273
R3177 VDDD.n3821 VDDD.n3820 9.73273
R3178 VDDD.n3823 VDDD.n3821 9.73273
R3179 VDDD.n3790 VDDD.n3789 9.73273
R3180 VDDD.n3791 VDDD.n3790 9.73273
R3181 VDDD.n3795 VDDD.n3794 9.73273
R3182 VDDD.n3796 VDDD.n3795 9.73273
R3183 VDDD.n3796 VDDD.n10 9.73273
R3184 VDDD.n3800 VDDD.n10 9.73273
R3185 VDDD.n3801 VDDD.n3800 9.73273
R3186 VDDD.n3802 VDDD.n3801 9.73273
R3187 VDDD.n3611 VDDD.n345 9.73273
R3188 VDDD.n3630 VDDD.n338 9.73273
R3189 VDDD.n3636 VDDD.n3635 9.73273
R3190 VDDD.n239 VDDD.n238 9.73273
R3191 VDDD.n3674 VDDD.n217 9.73273
R3192 VDDD.n3670 VDDD.n217 9.73273
R3193 VDDD.n3668 VDDD.n3667 9.73273
R3194 VDDD.n3664 VDDD.n3663 9.73273
R3195 VDDD.n3655 VDDD.n3654 9.73273
R3196 VDDD.n3649 VDDD.n3648 9.73273
R3197 VDDD.n3648 VDDD.n229 9.73273
R3198 VDDD.n3512 VDDD.n3509 9.73273
R3199 VDDD.n424 VDDD.n423 9.73273
R3200 VDDD.n432 VDDD.n429 9.73273
R3201 VDDD.n432 VDDD.n431 9.73273
R3202 VDDD.n448 VDDD.n381 9.73273
R3203 VDDD.n451 VDDD.n450 9.73273
R3204 VDDD.n729 VDDD.n728 9.73273
R3205 VDDD.n728 VDDD.n727 9.73273
R3206 VDDD.n3101 VDDD.n667 9.73273
R3207 VDDD.n3101 VDDD.n666 9.73273
R3208 VDDD.n3105 VDDD.n666 9.73273
R3209 VDDD.n3106 VDDD.n3105 9.73273
R3210 VDDD.n3110 VDDD.n3109 9.73273
R3211 VDDD.n3234 VDDD.n3175 9.73273
R3212 VDDD.n3230 VDDD.n3175 9.73273
R3213 VDDD.n3228 VDDD.n3227 9.73273
R3214 VDDD.n3227 VDDD.n3177 9.73273
R3215 VDDD.n3223 VDDD.n3177 9.73273
R3216 VDDD.n3213 VDDD.n3212 9.73273
R3217 VDDD.n3209 VDDD.n3208 9.73273
R3218 VDDD.n3206 VDDD.n3184 9.73273
R3219 VDDD.n3202 VDDD.n3201 9.73273
R3220 VDDD.n3062 VDDD.n3061 9.73273
R3221 VDDD.n3058 VDDD.n3057 9.73273
R3222 VDDD.n3055 VDDD.n761 9.73273
R3223 VDDD.n3051 VDDD.n3050 9.73273
R3224 VDDD.n3050 VDDD.n3049 9.73273
R3225 VDDD.n2973 VDDD.n2972 9.73273
R3226 VDDD.n2972 VDDD.n1136 9.73273
R3227 VDDD.n1231 VDDD.n1152 9.73273
R3228 VDDD.n1229 VDDD.n1228 9.73273
R3229 VDDD.n1223 VDDD.n1222 9.73273
R3230 VDDD.n1844 VDDD.n1843 9.73273
R3231 VDDD.n1843 VDDD.n1842 9.73273
R3232 VDDD.n1839 VDDD.n1838 9.73273
R3233 VDDD.n1838 VDDD.n1837 9.73273
R3234 VDDD.n1756 VDDD.n1755 9.73273
R3235 VDDD.n1750 VDDD.n1749 9.73273
R3236 VDDD.n1747 VDDD.n1733 9.73273
R3237 VDDD.n1779 VDDD.n1778 9.73273
R3238 VDDD.n1775 VDDD.n1774 9.73273
R3239 VDDD.n1774 VDDD.n1773 9.73273
R3240 VDDD.n1773 VDDD.n1710 9.73273
R3241 VDDD.n1726 VDDD.n1725 9.73273
R3242 VDDD.n2446 VDDD.n2445 9.73273
R3243 VDDD.n2576 VDDD.n1639 9.73273
R3244 VDDD.n2574 VDDD.n1641 9.73273
R3245 VDDD.n2132 VDDD.n2130 9.73273
R3246 VDDD.n2136 VDDD.n2135 9.73273
R3247 VDDD.n2106 VDDD.n2069 9.73273
R3248 VDDD.n2113 VDDD.n2067 9.73273
R3249 VDDD.n2114 VDDD.n2113 9.73273
R3250 VDDD.n2115 VDDD.n2114 9.73273
R3251 VDDD.n2119 VDDD.n2118 9.73273
R3252 VDDD.n2169 VDDD.n2168 9.73273
R3253 VDDD.n2171 VDDD.n2169 9.73273
R3254 VDDD.n2175 VDDD.n2039 9.73273
R3255 VDDD.n2178 VDDD.n2177 9.73273
R3256 VDDD.n2182 VDDD.n2181 9.73273
R3257 VDDD.n2183 VDDD.n2182 9.73273
R3258 VDDD.n2196 VDDD.n2032 9.73273
R3259 VDDD.n2013 VDDD.n2012 9.73273
R3260 VDDD.n2007 VDDD.n2006 9.73273
R3261 VDDD.n2006 VDDD.n2003 9.73273
R3262 VDDD.n2001 VDDD.n2000 9.73273
R3263 VDDD.n2323 VDDD.n2322 9.73273
R3264 VDDD.n2313 VDDD.n2312 9.73273
R3265 VDDD.n2307 VDDD.n2306 9.73273
R3266 VDDD.n91 VDDD.n90 9.73273
R3267 VDDD.n90 VDDD.n89 9.73273
R3268 VDDD.n86 VDDD.n85 9.73273
R3269 VDDD.n85 VDDD.n84 9.73273
R3270 VDDD.n84 VDDD.n76 9.73273
R3271 VDDD.n80 VDDD.n76 9.73273
R3272 VDDD.n80 VDDD.n79 9.73273
R3273 VDDD.n79 VDDD.n78 9.73273
R3274 VDDD.n67 VDDD.n60 9.73273
R3275 VDDD.n108 VDDD.n67 9.73273
R3276 VDDD.n106 VDDD.n105 9.73273
R3277 VDDD.n105 VDDD.n68 9.73273
R3278 VDDD.n101 VDDD.n68 9.73273
R3279 VDDD.n101 VDDD.n100 9.73273
R3280 VDDD.n100 VDDD.n99 9.73273
R3281 VDDD.n99 VDDD.n70 9.73273
R3282 VDDD.n194 VDDD.n193 9.73273
R3283 VDDD.n193 VDDD.n192 9.73273
R3284 VDDD.n189 VDDD.n188 9.73273
R3285 VDDD.n188 VDDD.n187 9.73273
R3286 VDDD.n187 VDDD.n176 9.73273
R3287 VDDD.n183 VDDD.n176 9.73273
R3288 VDDD.n183 VDDD.n182 9.73273
R3289 VDDD.n182 VDDD.n181 9.73273
R3290 VDDD.n151 VDDD.n150 9.73273
R3291 VDDD.n152 VDDD.n151 9.73273
R3292 VDDD.n156 VDDD.n155 9.73273
R3293 VDDD.n157 VDDD.n156 9.73273
R3294 VDDD.n157 VDDD.n120 9.73273
R3295 VDDD.n170 VDDD.n120 9.73273
R3296 VDDD.n171 VDDD.n170 9.73273
R3297 VDDD.n200 VDDD.n171 9.73273
R3298 VDDD.n1743 VDDD.n1742 9.71972
R3299 VDDD.n131 VDDD 9.6274
R3300 VDDD.n3832 VDDD.n3831 9.60526
R3301 VDDD.n3451 VDDD.n3296 9.6005
R3302 VDDD.n3650 VDDD.n3649 9.52116
R3303 VDDD.n3106 VDDD.n665 9.52116
R3304 VDDD.n1834 VDDD.n1826 9.52116
R3305 VDDD.n1748 VDDD.n1747 9.52116
R3306 VDDD.n2575 VDDD.n2574 9.52116
R3307 VDDD.n2308 VDDD.n2307 9.52116
R3308 VDDD.n1796 VDDD.n1687 9.50907
R3309 VDDD.n2701 VDDD.n1568 9.49016
R3310 VDDD.n313 VDDD.n312 9.41227
R3311 VDDD.n3596 VDDD.n3595 9.41227
R3312 VDDD.n3582 VDDD.n3581 9.41227
R3313 VDDD.n3568 VDDD.n269 9.41227
R3314 VDDD.n3543 VDDD.n3488 9.41227
R3315 VDDD.n3376 VDDD.n3338 9.41227
R3316 VDDD.n3385 VDDD.n3384 9.41227
R3317 VDDD.n741 VDDD.n740 9.41227
R3318 VDDD.n597 VDDD.n596 9.41227
R3319 VDDD.n1062 VDDD.n1061 9.41227
R3320 VDDD.n1019 VDDD.n886 9.41227
R3321 VDDD.n1014 VDDD.n1013 9.41227
R3322 VDDD.n972 VDDD.n971 9.41227
R3323 VDDD.n1500 VDDD.n1330 9.41227
R3324 VDDD.n1344 VDDD.n1343 9.41227
R3325 VDDD.n2839 VDDD.n2838 9.41227
R3326 VDDD.n2768 VDDD.n1274 9.41227
R3327 VDDD.n2720 VDDD.n2719 9.41227
R3328 VDDD.n2919 VDDD.n2871 9.41227
R3329 VDDD.n1621 VDDD.n1620 9.41227
R3330 VDDD.n1625 VDDD.n1578 9.41227
R3331 VDDD.n2657 VDDD.n2614 9.41227
R3332 VDDD.n1916 VDDD.n1906 9.41227
R3333 VDDD.n2397 VDDD.n1668 9.41227
R3334 VDDD.n2390 VDDD.n2389 9.41227
R3335 VDDD.n3750 VDDD.n29 9.41227
R3336 VDDD.n3632 VDDD.n336 9.30959
R3337 VDDD.n3508 VDDD.n3507 9.30959
R3338 VDDD.n267 VDDD.n232 9.3005
R3339 VDDD.n267 VDDD.n231 9.3005
R3340 VDDD.n267 VDDD.n230 9.3005
R3341 VDDD.n251 VDDD.n250 9.3005
R3342 VDDD.n248 VDDD.n235 9.3005
R3343 VDDD.n245 VDDD.n244 9.3005
R3344 VDDD.n243 VDDD.n242 9.3005
R3345 VDDD.n239 VDDD.n211 9.3005
R3346 VDDD.n238 VDDD.n212 9.3005
R3347 VDDD.n3677 VDDD.n3676 9.3005
R3348 VDDD.n3674 VDDD.n3673 9.3005
R3349 VDDD.n3672 VDDD.n217 9.3005
R3350 VDDD.n3671 VDDD.n3670 9.3005
R3351 VDDD.n3668 VDDD.n218 9.3005
R3352 VDDD.n3667 VDDD.n3666 9.3005
R3353 VDDD.n3665 VDDD.n3664 9.3005
R3354 VDDD.n3663 VDDD.n221 9.3005
R3355 VDDD.n3661 VDDD.n3660 9.3005
R3356 VDDD.n3659 VDDD.n222 9.3005
R3357 VDDD.n3658 VDDD.n3657 9.3005
R3358 VDDD.n3655 VDDD.n223 9.3005
R3359 VDDD.n3654 VDDD.n3653 9.3005
R3360 VDDD.n3652 VDDD.n3651 9.3005
R3361 VDDD.n3649 VDDD.n226 9.3005
R3362 VDDD.n3648 VDDD.n228 9.3005
R3363 VDDD.n3505 VDDD.n229 9.3005
R3364 VDDD.n3507 VDDD.n3506 9.3005
R3365 VDDD.n3509 VDDD.n3503 9.3005
R3366 VDDD.n3513 VDDD.n3512 9.3005
R3367 VDDD.n3515 VDDD.n3498 9.3005
R3368 VDDD.n3527 VDDD.n3526 9.3005
R3369 VDDD.n3531 VDDD.n3530 9.3005
R3370 VDDD.n3532 VDDD.n3495 9.3005
R3371 VDDD.n3534 VDDD.n3533 9.3005
R3372 VDDD.n3536 VDDD.n3494 9.3005
R3373 VDDD.n3537 VDDD.n3492 9.3005
R3374 VDDD.n3539 VDDD.n3538 9.3005
R3375 VDDD.n3541 VDDD.n3540 9.3005
R3376 VDDD.n3542 VDDD.n3489 9.3005
R3377 VDDD.n3544 VDDD.n3543 9.3005
R3378 VDDD.n3545 VDDD.n3488 9.3005
R3379 VDDD.n3547 VDDD.n3546 9.3005
R3380 VDDD.n3550 VDDD.n3486 9.3005
R3381 VDDD.n3552 VDDD.n3551 9.3005
R3382 VDDD.n3553 VDDD.n3485 9.3005
R3383 VDDD.n3555 VDDD.n3554 9.3005
R3384 VDDD.n3556 VDDD.n3483 9.3005
R3385 VDDD.n3560 VDDD.n3559 9.3005
R3386 VDDD.n3561 VDDD.n3482 9.3005
R3387 VDDD.n3563 VDDD.n3562 9.3005
R3388 VDDD.n3567 VDDD.n3566 9.3005
R3389 VDDD.n3569 VDDD.n3568 9.3005
R3390 VDDD.n3475 VDDD.n269 9.3005
R3391 VDDD.n3579 VDDD.n3578 9.3005
R3392 VDDD.n3580 VDDD.n358 9.3005
R3393 VDDD.n3581 VDDD.n356 9.3005
R3394 VDDD.n3582 VDDD.n353 9.3005
R3395 VDDD.n3584 VDDD.n3583 9.3005
R3396 VDDD.n3585 VDDD.n352 9.3005
R3397 VDDD.n3587 VDDD.n3586 9.3005
R3398 VDDD.n3588 VDDD.n351 9.3005
R3399 VDDD.n3592 VDDD.n3591 9.3005
R3400 VDDD.n3593 VDDD.n350 9.3005
R3401 VDDD.n3595 VDDD.n3594 9.3005
R3402 VDDD.n3596 VDDD.n348 9.3005
R3403 VDDD.n3598 VDDD.n3597 9.3005
R3404 VDDD.n3599 VDDD.n347 9.3005
R3405 VDDD.n3601 VDDD.n3600 9.3005
R3406 VDDD.n3604 VDDD.n346 9.3005
R3407 VDDD.n3608 VDDD.n3607 9.3005
R3408 VDDD.n3609 VDDD.n345 9.3005
R3409 VDDD.n3611 VDDD.n3610 9.3005
R3410 VDDD.n3616 VDDD.n3615 9.3005
R3411 VDDD.n3619 VDDD.n338 9.3005
R3412 VDDD.n3630 VDDD.n3629 9.3005
R3413 VDDD.n3633 VDDD.n3632 9.3005
R3414 VDDD.n3635 VDDD.n3634 9.3005
R3415 VDDD.n3636 VDDD.n335 9.3005
R3416 VDDD.n3639 VDDD.n3638 9.3005
R3417 VDDD.n3641 VDDD.n3640 9.3005
R3418 VDDD.n3644 VDDD.n333 9.3005
R3419 VDDD.n332 VDDD.n270 9.3005
R3420 VDDD.n331 VDDD.n330 9.3005
R3421 VDDD.n328 VDDD.n271 9.3005
R3422 VDDD.n326 VDDD.n325 9.3005
R3423 VDDD.n324 VDDD.n323 9.3005
R3424 VDDD.n320 VDDD.n273 9.3005
R3425 VDDD.n318 VDDD.n317 9.3005
R3426 VDDD.n316 VDDD.n274 9.3005
R3427 VDDD.n315 VDDD.n314 9.3005
R3428 VDDD.n313 VDDD.n275 9.3005
R3429 VDDD.n312 VDDD.n311 9.3005
R3430 VDDD.n310 VDDD.n276 9.3005
R3431 VDDD.n309 VDDD.n308 9.3005
R3432 VDDD.n306 VDDD.n277 9.3005
R3433 VDDD.n406 VDDD.n397 9.3005
R3434 VDDD.n407 VDDD.n397 9.3005
R3435 VDDD.n409 VDDD.n408 9.3005
R3436 VDDD.n412 VDDD.n392 9.3005
R3437 VDDD.n417 VDDD.n416 9.3005
R3438 VDDD.n418 VDDD.n391 9.3005
R3439 VDDD.n420 VDDD.n419 9.3005
R3440 VDDD.n423 VDDD.n390 9.3005
R3441 VDDD.n425 VDDD.n424 9.3005
R3442 VDDD.n427 VDDD.n426 9.3005
R3443 VDDD.n429 VDDD.n387 9.3005
R3444 VDDD.n433 VDDD.n432 9.3005
R3445 VDDD.n431 VDDD.n386 9.3005
R3446 VDDD.n439 VDDD.n381 9.3005
R3447 VDDD.n448 VDDD.n447 9.3005
R3448 VDDD.n450 VDDD.n379 9.3005
R3449 VDDD.n452 VDDD.n451 9.3005
R3450 VDDD.n454 VDDD.n453 9.3005
R3451 VDDD.n455 VDDD.n377 9.3005
R3452 VDDD.n457 VDDD.n456 9.3005
R3453 VDDD.n458 VDDD.n376 9.3005
R3454 VDDD.n460 VDDD.n459 9.3005
R3455 VDDD.n462 VDDD.n374 9.3005
R3456 VDDD.n466 VDDD.n465 9.3005
R3457 VDDD.n467 VDDD.n373 9.3005
R3458 VDDD.n469 VDDD.n468 9.3005
R3459 VDDD.n472 VDDD.n372 9.3005
R3460 VDDD.n476 VDDD.n475 9.3005
R3461 VDDD.n477 VDDD.n371 9.3005
R3462 VDDD.n3291 VDDD.n478 9.3005
R3463 VDDD.n3286 VDDD.n479 9.3005
R3464 VDDD.n488 VDDD.n479 9.3005
R3465 VDDD.n493 VDDD.n479 9.3005
R3466 VDDD.n557 VDDD.n479 9.3005
R3467 VDDD.n556 VDDD.n555 9.3005
R3468 VDDD.n553 VDDD.n495 9.3005
R3469 VDDD.n552 VDDD.n551 9.3005
R3470 VDDD.n550 VDDD.n549 9.3005
R3471 VDDD.n548 VDDD.n547 9.3005
R3472 VDDD.n545 VDDD.n544 9.3005
R3473 VDDD.n541 VDDD.n508 9.3005
R3474 VDDD.n539 VDDD.n538 9.3005
R3475 VDDD.n537 VDDD.n513 9.3005
R3476 VDDD.n536 VDDD.n535 9.3005
R3477 VDDD.n534 VDDD.n533 9.3005
R3478 VDDD.n532 VDDD.n531 9.3005
R3479 VDDD.n530 VDDD.n519 9.3005
R3480 VDDD.n529 VDDD.n528 9.3005
R3481 VDDD.n527 VDDD.n526 9.3005
R3482 VDDD.n524 VDDD.n366 9.3005
R3483 VDDD.n3466 VDDD.n3465 9.3005
R3484 VDDD.n3462 VDDD.n3461 9.3005
R3485 VDDD.n3453 VDDD.n3452 9.3005
R3486 VDDD.n3445 VDDD.n3444 9.3005
R3487 VDDD.n3442 VDDD.n3441 9.3005
R3488 VDDD.n3440 VDDD.n3300 9.3005
R3489 VDDD.n3439 VDDD.n3438 9.3005
R3490 VDDD.n3437 VDDD.n3436 9.3005
R3491 VDDD.n3433 VDDD.n3432 9.3005
R3492 VDDD.n3431 VDDD.n3430 9.3005
R3493 VDDD.n3427 VDDD.n3306 9.3005
R3494 VDDD.n3426 VDDD.n3307 9.3005
R3495 VDDD.n3425 VDDD.n3424 9.3005
R3496 VDDD.n3423 VDDD.n3309 9.3005
R3497 VDDD.n3422 VDDD.n3421 9.3005
R3498 VDDD.n3420 VDDD.n3312 9.3005
R3499 VDDD.n3418 VDDD.n3417 9.3005
R3500 VDDD.n3322 VDDD.n3313 9.3005
R3501 VDDD.n3409 VDDD.n3408 9.3005
R3502 VDDD.n3406 VDDD.n3323 9.3005
R3503 VDDD.n3405 VDDD.n3404 9.3005
R3504 VDDD.n3403 VDDD.n3402 9.3005
R3505 VDDD.n3399 VDDD.n3327 9.3005
R3506 VDDD.n3398 VDDD.n3328 9.3005
R3507 VDDD.n3395 VDDD.n3394 9.3005
R3508 VDDD.n3393 VDDD.n3392 9.3005
R3509 VDDD.n3390 VDDD.n3331 9.3005
R3510 VDDD.n3389 VDDD.n3388 9.3005
R3511 VDDD.n3387 VDDD.n3333 9.3005
R3512 VDDD.n3386 VDDD.n3385 9.3005
R3513 VDDD.n3384 VDDD.n3334 9.3005
R3514 VDDD.n3383 VDDD.n3382 9.3005
R3515 VDDD.n3381 VDDD.n3380 9.3005
R3516 VDDD.n3377 VDDD.n3337 9.3005
R3517 VDDD.n3376 VDDD.n3375 9.3005
R3518 VDDD.n3374 VDDD.n3338 9.3005
R3519 VDDD.n3373 VDDD.n3372 9.3005
R3520 VDDD.n3371 VDDD.n3339 9.3005
R3521 VDDD.n3370 VDDD.n3369 9.3005
R3522 VDDD.n3368 VDDD.n3367 9.3005
R3523 VDDD.n3365 VDDD.n3342 9.3005
R3524 VDDD.n678 VDDD.n668 9.3005
R3525 VDDD.n3098 VDDD.n3097 9.3005
R3526 VDDD.n3096 VDDD.n3095 9.3005
R3527 VDDD.n3094 VDDD.n3093 9.3005
R3528 VDDD.n3092 VDDD.n3091 9.3005
R3529 VDDD.n3090 VDDD.n682 9.3005
R3530 VDDD.n3089 VDDD.n3088 9.3005
R3531 VDDD.n3087 VDDD.n3086 9.3005
R3532 VDDD.n3085 VDDD.n3084 9.3005
R3533 VDDD.n3083 VDDD.n3082 9.3005
R3534 VDDD.n3081 VDDD.n686 9.3005
R3535 VDDD.n3080 VDDD.n3079 9.3005
R3536 VDDD.n697 VDDD.n690 9.3005
R3537 VDDD.n706 VDDD.n704 9.3005
R3538 VDDD.n707 VDDD.n695 9.3005
R3539 VDDD.n744 VDDD.n743 9.3005
R3540 VDDD.n742 VDDD.n696 9.3005
R3541 VDDD.n741 VDDD.n710 9.3005
R3542 VDDD.n740 VDDD.n739 9.3005
R3543 VDDD.n738 VDDD.n711 9.3005
R3544 VDDD.n737 VDDD.n736 9.3005
R3545 VDDD.n735 VDDD.n712 9.3005
R3546 VDDD.n734 VDDD.n717 9.3005
R3547 VDDD.n733 VDDD.n732 9.3005
R3548 VDDD.n731 VDDD.n718 9.3005
R3549 VDDD.n730 VDDD.n729 9.3005
R3550 VDDD.n728 VDDD.n719 9.3005
R3551 VDDD.n727 VDDD.n726 9.3005
R3552 VDDD.n725 VDDD.n667 9.3005
R3553 VDDD.n3102 VDDD.n3101 9.3005
R3554 VDDD.n3103 VDDD.n666 9.3005
R3555 VDDD.n3105 VDDD.n3104 9.3005
R3556 VDDD.n3107 VDDD.n3106 9.3005
R3557 VDDD.n3109 VDDD.n3108 9.3005
R3558 VDDD.n3111 VDDD.n3110 9.3005
R3559 VDDD.n3123 VDDD.n3122 9.3005
R3560 VDDD.n3125 VDDD.n3124 9.3005
R3561 VDDD.n3126 VDDD.n654 9.3005
R3562 VDDD.n3128 VDDD.n3127 9.3005
R3563 VDDD.n3130 VDDD.n652 9.3005
R3564 VDDD.n3134 VDDD.n3133 9.3005
R3565 VDDD.n3136 VDDD.n3135 9.3005
R3566 VDDD.n3137 VDDD.n648 9.3005
R3567 VDDD.n3141 VDDD.n3140 9.3005
R3568 VDDD.n3142 VDDD.n647 9.3005
R3569 VDDD.n3144 VDDD.n3143 9.3005
R3570 VDDD.n3145 VDDD.n645 9.3005
R3571 VDDD.n3146 VDDD.n643 9.3005
R3572 VDDD.n3148 VDDD.n3147 9.3005
R3573 VDDD.n3150 VDDD.n636 9.3005
R3574 VDDD.n3152 VDDD.n3151 9.3005
R3575 VDDD.n3154 VDDD.n3153 9.3005
R3576 VDDD.n3159 VDDD.n3158 9.3005
R3577 VDDD.n3169 VDDD.n3168 9.3005
R3578 VDDD.n618 VDDD.n617 9.3005
R3579 VDDD.n615 VDDD.n614 9.3005
R3580 VDDD.n613 VDDD.n581 9.3005
R3581 VDDD.n612 VDDD.n611 9.3005
R3582 VDDD.n609 VDDD.n608 9.3005
R3583 VDDD.n607 VDDD.n606 9.3005
R3584 VDDD.n605 VDDD.n584 9.3005
R3585 VDDD.n603 VDDD.n602 9.3005
R3586 VDDD.n601 VDDD.n586 9.3005
R3587 VDDD.n600 VDDD.n599 9.3005
R3588 VDDD.n597 VDDD.n587 9.3005
R3589 VDDD.n596 VDDD.n593 9.3005
R3590 VDDD.n595 VDDD.n594 9.3005
R3591 VDDD.n570 VDDD.n568 9.3005
R3592 VDDD.n3271 VDDD.n3270 9.3005
R3593 VDDD.n3267 VDDD.n3266 9.3005
R3594 VDDD.n3259 VDDD.n3258 9.3005
R3595 VDDD.n3255 VDDD.n573 9.3005
R3596 VDDD.n3254 VDDD.n3253 9.3005
R3597 VDDD.n3252 VDDD.n3251 9.3005
R3598 VDDD.n3249 VDDD.n575 9.3005
R3599 VDDD.n3248 VDDD.n3247 9.3005
R3600 VDDD.n3246 VDDD.n3245 9.3005
R3601 VDDD.n3238 VDDD.n3237 9.3005
R3602 VDDD.n3234 VDDD.n3233 9.3005
R3603 VDDD.n3232 VDDD.n3175 9.3005
R3604 VDDD.n3231 VDDD.n3230 9.3005
R3605 VDDD.n3228 VDDD.n3176 9.3005
R3606 VDDD.n3227 VDDD.n3226 9.3005
R3607 VDDD.n3225 VDDD.n3177 9.3005
R3608 VDDD.n3224 VDDD.n3223 9.3005
R3609 VDDD.n3221 VDDD.n3178 9.3005
R3610 VDDD.n3218 VDDD.n3217 9.3005
R3611 VDDD.n3216 VDDD.n3215 9.3005
R3612 VDDD.n3213 VDDD.n3180 9.3005
R3613 VDDD.n3212 VDDD.n3211 9.3005
R3614 VDDD.n3210 VDDD.n3209 9.3005
R3615 VDDD.n3208 VDDD.n3182 9.3005
R3616 VDDD.n3206 VDDD.n3205 9.3005
R3617 VDDD.n3204 VDDD.n3184 9.3005
R3618 VDDD.n3203 VDDD.n3202 9.3005
R3619 VDDD.n3201 VDDD.n3185 9.3005
R3620 VDDD.n3199 VDDD.n3198 9.3005
R3621 VDDD.n3197 VDDD.n3196 9.3005
R3622 VDDD.n809 VDDD.n783 9.3005
R3623 VDDD.n809 VDDD.n808 9.3005
R3624 VDDD.n801 VDDD.n800 9.3005
R3625 VDDD.n798 VDDD.n785 9.3005
R3626 VDDD.n796 VDDD.n795 9.3005
R3627 VDDD.n794 VDDD.n793 9.3005
R3628 VDDD.n791 VDDD.n753 9.3005
R3629 VDDD.n789 VDDD.n754 9.3005
R3630 VDDD.n3063 VDDD.n3062 9.3005
R3631 VDDD.n3061 VDDD.n3060 9.3005
R3632 VDDD.n3059 VDDD.n3058 9.3005
R3633 VDDD.n3057 VDDD.n760 9.3005
R3634 VDDD.n3055 VDDD.n3054 9.3005
R3635 VDDD.n3053 VDDD.n761 9.3005
R3636 VDDD.n3052 VDDD.n3051 9.3005
R3637 VDDD.n3050 VDDD.n762 9.3005
R3638 VDDD.n3049 VDDD.n3048 9.3005
R3639 VDDD.n3047 VDDD.n3046 9.3005
R3640 VDDD.n3045 VDDD.n766 9.3005
R3641 VDDD.n3043 VDDD.n3042 9.3005
R3642 VDDD.n3041 VDDD.n768 9.3005
R3643 VDDD.n3040 VDDD.n3039 9.3005
R3644 VDDD.n3037 VDDD.n769 9.3005
R3645 VDDD.n3035 VDDD.n3034 9.3005
R3646 VDDD.n3033 VDDD.n812 9.3005
R3647 VDDD.n3032 VDDD.n3031 9.3005
R3648 VDDD.n3029 VDDD.n813 9.3005
R3649 VDDD.n3027 VDDD.n3026 9.3005
R3650 VDDD.n830 VDDD.n829 9.3005
R3651 VDDD.n837 VDDD.n836 9.3005
R3652 VDDD.n1088 VDDD.n1087 9.3005
R3653 VDDD.n1085 VDDD.n826 9.3005
R3654 VDDD.n1082 VDDD.n1081 9.3005
R3655 VDDD.n1080 VDDD.n840 9.3005
R3656 VDDD.n1079 VDDD.n1078 9.3005
R3657 VDDD.n1077 VDDD.n1076 9.3005
R3658 VDDD.n1075 VDDD.n1074 9.3005
R3659 VDDD.n1073 VDDD.n844 9.3005
R3660 VDDD.n1072 VDDD.n1071 9.3005
R3661 VDDD.n1070 VDDD.n1069 9.3005
R3662 VDDD.n1068 VDDD.n848 9.3005
R3663 VDDD.n1067 VDDD.n1066 9.3005
R3664 VDDD.n1065 VDDD.n1064 9.3005
R3665 VDDD.n1063 VDDD.n852 9.3005
R3666 VDDD.n1062 VDDD.n853 9.3005
R3667 VDDD.n1061 VDDD.n1060 9.3005
R3668 VDDD.n1059 VDDD.n854 9.3005
R3669 VDDD.n1058 VDDD.n1057 9.3005
R3670 VDDD.n1056 VDDD.n855 9.3005
R3671 VDDD.n1055 VDDD.n860 9.3005
R3672 VDDD.n1054 VDDD.n1053 9.3005
R3673 VDDD.n871 VDDD.n861 9.3005
R3674 VDDD.n1045 VDDD.n1044 9.3005
R3675 VDDD.n1043 VDDD.n1042 9.3005
R3676 VDDD.n1041 VDDD.n1040 9.3005
R3677 VDDD.n1038 VDDD.n874 9.3005
R3678 VDDD.n1037 VDDD.n1036 9.3005
R3679 VDDD.n1035 VDDD.n1034 9.3005
R3680 VDDD.n1032 VDDD.n878 9.3005
R3681 VDDD.n1031 VDDD.n1030 9.3005
R3682 VDDD.n1029 VDDD.n1028 9.3005
R3683 VDDD.n1027 VDDD.n880 9.3005
R3684 VDDD.n1026 VDDD.n1025 9.3005
R3685 VDDD.n1024 VDDD.n883 9.3005
R3686 VDDD.n1023 VDDD.n1022 9.3005
R3687 VDDD.n1020 VDDD.n884 9.3005
R3688 VDDD.n1019 VDDD.n1018 9.3005
R3689 VDDD.n1017 VDDD.n886 9.3005
R3690 VDDD.n1016 VDDD.n1015 9.3005
R3691 VDDD.n1014 VDDD.n887 9.3005
R3692 VDDD.n1013 VDDD.n890 9.3005
R3693 VDDD.n1012 VDDD.n891 9.3005
R3694 VDDD.n1011 VDDD.n1010 9.3005
R3695 VDDD.n906 VDDD.n903 9.3005
R3696 VDDD.n1002 VDDD.n1001 9.3005
R3697 VDDD.n999 VDDD.n904 9.3005
R3698 VDDD.n996 VDDD.n995 9.3005
R3699 VDDD.n994 VDDD.n908 9.3005
R3700 VDDD.n993 VDDD.n992 9.3005
R3701 VDDD.n990 VDDD.n989 9.3005
R3702 VDDD.n988 VDDD.n911 9.3005
R3703 VDDD.n987 VDDD.n986 9.3005
R3704 VDDD.n985 VDDD.n912 9.3005
R3705 VDDD.n983 VDDD.n982 9.3005
R3706 VDDD.n981 VDDD.n917 9.3005
R3707 VDDD.n980 VDDD.n979 9.3005
R3708 VDDD.n978 VDDD.n918 9.3005
R3709 VDDD.n977 VDDD.n976 9.3005
R3710 VDDD.n975 VDDD.n920 9.3005
R3711 VDDD.n974 VDDD.n973 9.3005
R3712 VDDD.n972 VDDD.n921 9.3005
R3713 VDDD.n971 VDDD.n924 9.3005
R3714 VDDD.n970 VDDD.n969 9.3005
R3715 VDDD.n968 VDDD.n967 9.3005
R3716 VDDD.n966 VDDD.n927 9.3005
R3717 VDDD.n963 VDDD.n962 9.3005
R3718 VDDD.n961 VDDD.n929 9.3005
R3719 VDDD.n960 VDDD.n959 9.3005
R3720 VDDD.n958 VDDD.n930 9.3005
R3721 VDDD.n957 VDDD.n933 9.3005
R3722 VDDD.n956 VDDD.n934 9.3005
R3723 VDDD.n954 VDDD.n953 9.3005
R3724 VDDD.n952 VDDD.n951 9.3005
R3725 VDDD.n949 VDDD.n936 9.3005
R3726 VDDD.n947 VDDD.n946 9.3005
R3727 VDDD.n1447 VDDD.n1438 9.3005
R3728 VDDD.n1481 VDDD.n1480 9.3005
R3729 VDDD.n1479 VDDD.n1437 9.3005
R3730 VDDD.n1478 VDDD.n1477 9.3005
R3731 VDDD.n1473 VDDD.n1448 9.3005
R3732 VDDD.n1472 VDDD.n1471 9.3005
R3733 VDDD.n1470 VDDD.n1469 9.3005
R3734 VDDD.n1468 VDDD.n1467 9.3005
R3735 VDDD.n1466 VDDD.n1452 9.3005
R3736 VDDD.n1465 VDDD.n1464 9.3005
R3737 VDDD.n1462 VDDD.n1453 9.3005
R3738 VDDD.n1460 VDDD.n1459 9.3005
R3739 VDDD.n1456 VDDD.n1325 9.3005
R3740 VDDD.n1329 VDDD.n1326 9.3005
R3741 VDDD.n1506 VDDD.n1505 9.3005
R3742 VDDD.n1504 VDDD.n1503 9.3005
R3743 VDDD.n1502 VDDD.n1330 9.3005
R3744 VDDD.n1501 VDDD.n1500 9.3005
R3745 VDDD.n1499 VDDD.n1331 9.3005
R3746 VDDD.n1497 VDDD.n1496 9.3005
R3747 VDDD.n1495 VDDD.n1494 9.3005
R3748 VDDD.n1491 VDDD.n1490 9.3005
R3749 VDDD.n1489 VDDD.n1336 9.3005
R3750 VDDD.n1487 VDDD.n1486 9.3005
R3751 VDDD.n1485 VDDD.n1484 9.3005
R3752 VDDD.n1483 VDDD.n1341 9.3005
R3753 VDDD.n1435 VDDD.n1434 9.3005
R3754 VDDD.n1433 VDDD.n1343 9.3005
R3755 VDDD.n1432 VDDD.n1431 9.3005
R3756 VDDD.n1429 VDDD.n1428 9.3005
R3757 VDDD.n1357 VDDD.n1356 9.3005
R3758 VDDD.n1362 VDDD.n1361 9.3005
R3759 VDDD.n1419 VDDD.n1418 9.3005
R3760 VDDD.n1417 VDDD.n1351 9.3005
R3761 VDDD.n1415 VDDD.n1414 9.3005
R3762 VDDD.n1413 VDDD.n1412 9.3005
R3763 VDDD.n1411 VDDD.n1365 9.3005
R3764 VDDD.n1408 VDDD.n1407 9.3005
R3765 VDDD.n1406 VDDD.n1368 9.3005
R3766 VDDD.n1405 VDDD.n1404 9.3005
R3767 VDDD.n1403 VDDD.n1369 9.3005
R3768 VDDD.n1402 VDDD.n1401 9.3005
R3769 VDDD.n1400 VDDD.n1373 9.3005
R3770 VDDD.n1399 VDDD.n1398 9.3005
R3771 VDDD.n1396 VDDD.n1381 9.3005
R3772 VDDD.n1395 VDDD.n1394 9.3005
R3773 VDDD.n1393 VDDD.n1382 9.3005
R3774 VDDD.n1392 VDDD.n1391 9.3005
R3775 VDDD.n1388 VDDD.n1383 9.3005
R3776 VDDD.n1386 VDDD.n1099 9.3005
R3777 VDDD.n3012 VDDD.n3011 9.3005
R3778 VDDD.n3009 VDDD.n1102 9.3005
R3779 VDDD.n3008 VDDD.n1111 9.3005
R3780 VDDD.n3006 VDDD.n3005 9.3005
R3781 VDDD.n3004 VDDD.n1113 9.3005
R3782 VDDD.n3003 VDDD.n3002 9.3005
R3783 VDDD.n3001 VDDD.n1114 9.3005
R3784 VDDD.n2998 VDDD.n2997 9.3005
R3785 VDDD.n2996 VDDD.n1120 9.3005
R3786 VDDD.n2995 VDDD.n2994 9.3005
R3787 VDDD.n2993 VDDD.n1121 9.3005
R3788 VDDD.n2992 VDDD.n2991 9.3005
R3789 VDDD.n2990 VDDD.n2989 9.3005
R3790 VDDD.n2987 VDDD.n1128 9.3005
R3791 VDDD.n2986 VDDD.n2985 9.3005
R3792 VDDD.n2984 VDDD.n1129 9.3005
R3793 VDDD.n2983 VDDD.n2982 9.3005
R3794 VDDD.n2980 VDDD.n1130 9.3005
R3795 VDDD.n2978 VDDD.n2977 9.3005
R3796 VDDD.n2976 VDDD.n2975 9.3005
R3797 VDDD.n2973 VDDD.n1135 9.3005
R3798 VDDD.n2972 VDDD.n2971 9.3005
R3799 VDDD.n1138 VDDD.n1136 9.3005
R3800 VDDD.n1152 VDDD.n1147 9.3005
R3801 VDDD.n1232 VDDD.n1231 9.3005
R3802 VDDD.n1229 VDDD.n1148 9.3005
R3803 VDDD.n1228 VDDD.n1227 9.3005
R3804 VDDD.n1226 VDDD.n1225 9.3005
R3805 VDDD.n1223 VDDD.n1154 9.3005
R3806 VDDD.n1222 VDDD.n1221 9.3005
R3807 VDDD.n1220 VDDD.n1219 9.3005
R3808 VDDD.n1218 VDDD.n1217 9.3005
R3809 VDDD.n1216 VDDD.n1215 9.3005
R3810 VDDD.n1214 VDDD.n1158 9.3005
R3811 VDDD.n1213 VDDD.n1212 9.3005
R3812 VDDD.n1211 VDDD.n1210 9.3005
R3813 VDDD.n1209 VDDD.n1160 9.3005
R3814 VDDD.n1208 VDDD.n1207 9.3005
R3815 VDDD.n1206 VDDD.n1161 9.3005
R3816 VDDD.n1205 VDDD.n1204 9.3005
R3817 VDDD.n1203 VDDD.n1162 9.3005
R3818 VDDD.n1202 VDDD.n1201 9.3005
R3819 VDDD.n1200 VDDD.n1199 9.3005
R3820 VDDD.n1198 VDDD.n1197 9.3005
R3821 VDDD.n1196 VDDD.n1195 9.3005
R3822 VDDD.n1194 VDDD.n1165 9.3005
R3823 VDDD.n1193 VDDD.n1192 9.3005
R3824 VDDD.n1191 VDDD.n1190 9.3005
R3825 VDDD.n1189 VDDD.n1167 9.3005
R3826 VDDD.n1188 VDDD.n1187 9.3005
R3827 VDDD.n1186 VDDD.n1168 9.3005
R3828 VDDD.n1185 VDDD.n1184 9.3005
R3829 VDDD.n1183 VDDD.n1169 9.3005
R3830 VDDD.n1182 VDDD.n1181 9.3005
R3831 VDDD.n1180 VDDD.n1179 9.3005
R3832 VDDD.n1305 VDDD.n1295 9.3005
R3833 VDDD.n2738 VDDD.n2737 9.3005
R3834 VDDD.n2736 VDDD.n2735 9.3005
R3835 VDDD.n2734 VDDD.n1306 9.3005
R3836 VDDD.n2732 VDDD.n2731 9.3005
R3837 VDDD.n2730 VDDD.n2729 9.3005
R3838 VDDD.n2727 VDDD.n1308 9.3005
R3839 VDDD.n2726 VDDD.n1311 9.3005
R3840 VDDD.n2725 VDDD.n2724 9.3005
R3841 VDDD.n2723 VDDD.n1312 9.3005
R3842 VDDD.n2722 VDDD.n2721 9.3005
R3843 VDDD.n2720 VDDD.n1313 9.3005
R3844 VDDD.n2719 VDDD.n2718 9.3005
R3845 VDDD.n1524 VDDD.n1523 9.3005
R3846 VDDD.n1527 VDDD.n1520 9.3005
R3847 VDDD.n1557 VDDD.n1556 9.3005
R3848 VDDD.n1555 VDDD.n1521 9.3005
R3849 VDDD.n1554 VDDD.n1528 9.3005
R3850 VDDD.n1553 VDDD.n1529 9.3005
R3851 VDDD.n1552 VDDD.n1551 9.3005
R3852 VDDD.n1550 VDDD.n1531 9.3005
R3853 VDDD.n1549 VDDD.n1548 9.3005
R3854 VDDD.n1547 VDDD.n1546 9.3005
R3855 VDDD.n1545 VDDD.n1533 9.3005
R3856 VDDD.n1544 VDDD.n1543 9.3005
R3857 VDDD.n1542 VDDD.n1534 9.3005
R3858 VDDD.n1541 VDDD.n1540 9.3005
R3859 VDDD.n1539 VDDD.n1537 9.3005
R3860 VDDD.n1538 VDDD.n1293 9.3005
R3861 VDDD.n2741 VDDD.n1294 9.3005
R3862 VDDD.n2743 VDDD.n1292 9.3005
R3863 VDDD.n2744 VDDD.n1291 9.3005
R3864 VDDD.n2747 VDDD.n2746 9.3005
R3865 VDDD.n2749 VDDD.n2748 9.3005
R3866 VDDD.n2752 VDDD.n2751 9.3005
R3867 VDDD.n1285 VDDD.n1277 9.3005
R3868 VDDD.n2762 VDDD.n2761 9.3005
R3869 VDDD.n2763 VDDD.n1275 9.3005
R3870 VDDD.n2765 VDDD.n2764 9.3005
R3871 VDDD.n2766 VDDD.n1274 9.3005
R3872 VDDD.n2768 VDDD.n2767 9.3005
R3873 VDDD.n2770 VDDD.n1271 9.3005
R3874 VDDD.n2773 VDDD.n2772 9.3005
R3875 VDDD.n2774 VDDD.n1270 9.3005
R3876 VDDD.n2776 VDDD.n2775 9.3005
R3877 VDDD.n2777 VDDD.n1269 9.3005
R3878 VDDD.n2778 VDDD.n1268 9.3005
R3879 VDDD.n2779 VDDD.n1266 9.3005
R3880 VDDD.n2781 VDDD.n2780 9.3005
R3881 VDDD.n2782 VDDD.n1265 9.3005
R3882 VDDD.n2784 VDDD.n2783 9.3005
R3883 VDDD.n2785 VDDD.n1260 9.3005
R3884 VDDD.n2788 VDDD.n2787 9.3005
R3885 VDDD.n2789 VDDD.n1259 9.3005
R3886 VDDD.n2791 VDDD.n2790 9.3005
R3887 VDDD.n2794 VDDD.n2793 9.3005
R3888 VDDD.n2858 VDDD.n2857 9.3005
R3889 VDDD.n2859 VDDD.n1252 9.3005
R3890 VDDD.n2849 VDDD.n1251 9.3005
R3891 VDDD.n2848 VDDD.n2847 9.3005
R3892 VDDD.n2845 VDDD.n2800 9.3005
R3893 VDDD.n2844 VDDD.n2843 9.3005
R3894 VDDD.n2842 VDDD.n2801 9.3005
R3895 VDDD.n2841 VDDD.n2840 9.3005
R3896 VDDD.n2839 VDDD.n2802 9.3005
R3897 VDDD.n2838 VDDD.n2837 9.3005
R3898 VDDD.n2836 VDDD.n2805 9.3005
R3899 VDDD.n2835 VDDD.n2834 9.3005
R3900 VDDD.n2833 VDDD.n2806 9.3005
R3901 VDDD.n2830 VDDD.n2829 9.3005
R3902 VDDD.n2828 VDDD.n2810 9.3005
R3903 VDDD.n2827 VDDD.n2826 9.3005
R3904 VDDD.n2825 VDDD.n2811 9.3005
R3905 VDDD.n2824 VDDD.n2823 9.3005
R3906 VDDD.n2822 VDDD.n2813 9.3005
R3907 VDDD.n2821 VDDD.n2820 9.3005
R3908 VDDD.n2819 VDDD.n2815 9.3005
R3909 VDDD.n2818 VDDD.n1241 9.3005
R3910 VDDD.n2959 VDDD.n2958 9.3005
R3911 VDDD.n2956 VDDD.n2955 9.3005
R3912 VDDD.n2948 VDDD.n1244 9.3005
R3913 VDDD.n2947 VDDD.n2946 9.3005
R3914 VDDD.n2944 VDDD.n1246 9.3005
R3915 VDDD.n2943 VDDD.n2942 9.3005
R3916 VDDD.n2941 VDDD.n2940 9.3005
R3917 VDDD.n2939 VDDD.n1250 9.3005
R3918 VDDD.n2938 VDDD.n2937 9.3005
R3919 VDDD.n2936 VDDD.n2863 9.3005
R3920 VDDD.n2935 VDDD.n2934 9.3005
R3921 VDDD.n2933 VDDD.n2864 9.3005
R3922 VDDD.n2932 VDDD.n2865 9.3005
R3923 VDDD.n2931 VDDD.n2930 9.3005
R3924 VDDD.n2929 VDDD.n2866 9.3005
R3925 VDDD.n2928 VDDD.n2927 9.3005
R3926 VDDD.n2926 VDDD.n2867 9.3005
R3927 VDDD.n2923 VDDD.n2922 9.3005
R3928 VDDD.n2921 VDDD.n2871 9.3005
R3929 VDDD.n2920 VDDD.n2919 9.3005
R3930 VDDD.n2918 VDDD.n2872 9.3005
R3931 VDDD.n2917 VDDD.n2874 9.3005
R3932 VDDD.n2916 VDDD.n2915 9.3005
R3933 VDDD.n2914 VDDD.n2913 9.3005
R3934 VDDD.n2912 VDDD.n2876 9.3005
R3935 VDDD.n2909 VDDD.n2908 9.3005
R3936 VDDD.n2907 VDDD.n2906 9.3005
R3937 VDDD.n2904 VDDD.n2903 9.3005
R3938 VDDD.n2902 VDDD.n2901 9.3005
R3939 VDDD.n2900 VDDD.n2899 9.3005
R3940 VDDD.n2898 VDDD.n2882 9.3005
R3941 VDDD.n2897 VDDD.n2896 9.3005
R3942 VDDD.n2894 VDDD.n2883 9.3005
R3943 VDDD.n1699 VDDD.n1690 9.3005
R3944 VDDD.n1793 VDDD.n1700 9.3005
R3945 VDDD.n1790 VDDD.n1789 9.3005
R3946 VDDD.n1788 VDDD.n1701 9.3005
R3947 VDDD.n1787 VDDD.n1786 9.3005
R3948 VDDD.n1784 VDDD.n1783 9.3005
R3949 VDDD.n1782 VDDD.n1781 9.3005
R3950 VDDD.n1779 VDDD.n1705 9.3005
R3951 VDDD.n1778 VDDD.n1777 9.3005
R3952 VDDD.n1776 VDDD.n1775 9.3005
R3953 VDDD.n1774 VDDD.n1708 9.3005
R3954 VDDD.n1773 VDDD.n1772 9.3005
R3955 VDDD.n1711 VDDD.n1710 9.3005
R3956 VDDD.n1725 VDDD.n1724 9.3005
R3957 VDDD.n1726 VDDD.n1716 9.3005
R3958 VDDD.n1763 VDDD.n1762 9.3005
R3959 VDDD.n1760 VDDD.n1717 9.3005
R3960 VDDD.n1759 VDDD.n1758 9.3005
R3961 VDDD.n1757 VDDD.n1756 9.3005
R3962 VDDD.n1755 VDDD.n1729 9.3005
R3963 VDDD.n1753 VDDD.n1752 9.3005
R3964 VDDD.n1751 VDDD.n1750 9.3005
R3965 VDDD.n1749 VDDD.n1731 9.3005
R3966 VDDD.n1747 VDDD.n1746 9.3005
R3967 VDDD.n1745 VDDD.n1733 9.3005
R3968 VDDD.n1744 VDDD.n1743 9.3005
R3969 VDDD.n1742 VDDD.n1734 9.3005
R3970 VDDD.n1740 VDDD.n1739 9.3005
R3971 VDDD.n1738 VDDD.n1689 9.3005
R3972 VDDD.n1797 VDDD.n1796 9.3005
R3973 VDDD.n1798 VDDD.n1687 9.3005
R3974 VDDD.n1800 VDDD.n1799 9.3005
R3975 VDDD.n1803 VDDD.n1802 9.3005
R3976 VDDD.n1805 VDDD.n1804 9.3005
R3977 VDDD.n1877 VDDD.n1876 9.3005
R3978 VDDD.n1875 VDDD.n1874 9.3005
R3979 VDDD.n1866 VDDD.n1865 9.3005
R3980 VDDD.n1864 VDDD.n1810 9.3005
R3981 VDDD.n1861 VDDD.n1860 9.3005
R3982 VDDD.n1859 VDDD.n1814 9.3005
R3983 VDDD.n1858 VDDD.n1857 9.3005
R3984 VDDD.n1856 VDDD.n1815 9.3005
R3985 VDDD.n1853 VDDD.n1852 9.3005
R3986 VDDD.n1851 VDDD.n1850 9.3005
R3987 VDDD.n1848 VDDD.n1847 9.3005
R3988 VDDD.n1846 VDDD.n1819 9.3005
R3989 VDDD.n1845 VDDD.n1844 9.3005
R3990 VDDD.n1843 VDDD.n1820 9.3005
R3991 VDDD.n1842 VDDD.n1841 9.3005
R3992 VDDD.n1840 VDDD.n1839 9.3005
R3993 VDDD.n1838 VDDD.n1823 9.3005
R3994 VDDD.n1837 VDDD.n1836 9.3005
R3995 VDDD.n1835 VDDD.n1834 9.3005
R3996 VDDD.n1832 VDDD.n1831 9.3005
R3997 VDDD.n2702 VDDD.n2701 9.3005
R3998 VDDD.n2692 VDDD.n2691 9.3005
R3999 VDDD.n2693 VDDD.n2692 9.3005
R4000 VDDD.n1600 VDDD.n1599 9.3005
R4001 VDDD.n1604 VDDD.n1603 9.3005
R4002 VDDD.n1605 VDDD.n1595 9.3005
R4003 VDDD.n1607 VDDD.n1606 9.3005
R4004 VDDD.n1611 VDDD.n1610 9.3005
R4005 VDDD.n1612 VDDD.n1593 9.3005
R4006 VDDD.n1614 VDDD.n1613 9.3005
R4007 VDDD.n1615 VDDD.n1592 9.3005
R4008 VDDD.n1617 VDDD.n1616 9.3005
R4009 VDDD.n1619 VDDD.n1618 9.3005
R4010 VDDD.n1620 VDDD.n1589 9.3005
R4011 VDDD.n1622 VDDD.n1621 9.3005
R4012 VDDD.n1624 VDDD.n1623 9.3005
R4013 VDDD.n1626 VDDD.n1625 9.3005
R4014 VDDD.n1627 VDDD.n1578 9.3005
R4015 VDDD.n2590 VDDD.n2588 9.3005
R4016 VDDD.n2592 VDDD.n2591 9.3005
R4017 VDDD.n2594 VDDD.n2593 9.3005
R4018 VDDD.n2596 VDDD.n1574 9.3005
R4019 VDDD.n2601 VDDD.n2600 9.3005
R4020 VDDD.n2602 VDDD.n1572 9.3005
R4021 VDDD.n2681 VDDD.n2680 9.3005
R4022 VDDD.n2679 VDDD.n2678 9.3005
R4023 VDDD.n2677 VDDD.n2603 9.3005
R4024 VDDD.n2676 VDDD.n2675 9.3005
R4025 VDDD.n2674 VDDD.n2606 9.3005
R4026 VDDD.n2673 VDDD.n2672 9.3005
R4027 VDDD.n2671 VDDD.n2607 9.3005
R4028 VDDD.n2670 VDDD.n2608 9.3005
R4029 VDDD.n2669 VDDD.n2668 9.3005
R4030 VDDD.n2667 VDDD.n2609 9.3005
R4031 VDDD.n2666 VDDD.n2665 9.3005
R4032 VDDD.n2664 VDDD.n2610 9.3005
R4033 VDDD.n2661 VDDD.n2660 9.3005
R4034 VDDD.n2659 VDDD.n2614 9.3005
R4035 VDDD.n2658 VDDD.n2657 9.3005
R4036 VDDD.n2656 VDDD.n2615 9.3005
R4037 VDDD.n2655 VDDD.n2616 9.3005
R4038 VDDD.n2654 VDDD.n2653 9.3005
R4039 VDDD.n2652 VDDD.n2651 9.3005
R4040 VDDD.n2650 VDDD.n2619 9.3005
R4041 VDDD.n2647 VDDD.n2646 9.3005
R4042 VDDD.n2645 VDDD.n2644 9.3005
R4043 VDDD.n2642 VDDD.n2641 9.3005
R4044 VDDD.n2640 VDDD.n2639 9.3005
R4045 VDDD.n2638 VDDD.n2637 9.3005
R4046 VDDD.n2636 VDDD.n2635 9.3005
R4047 VDDD.n1898 VDDD.n1889 9.3005
R4048 VDDD.n2359 VDDD.n1899 9.3005
R4049 VDDD.n2357 VDDD.n2356 9.3005
R4050 VDDD.n2355 VDDD.n1900 9.3005
R4051 VDDD.n2354 VDDD.n2353 9.3005
R4052 VDDD.n2351 VDDD.n1901 9.3005
R4053 VDDD.n2349 VDDD.n2347 9.3005
R4054 VDDD.n2346 VDDD.n1904 9.3005
R4055 VDDD.n2345 VDDD.n2344 9.3005
R4056 VDDD.n2343 VDDD.n1905 9.3005
R4057 VDDD.n2342 VDDD.n2341 9.3005
R4058 VDDD.n2340 VDDD.n1906 9.3005
R4059 VDDD.n1916 VDDD.n1907 9.3005
R4060 VDDD.n1925 VDDD.n1924 9.3005
R4061 VDDD.n1927 VDDD.n1912 9.3005
R4062 VDDD.n1955 VDDD.n1954 9.3005
R4063 VDDD.n1953 VDDD.n1913 9.3005
R4064 VDDD.n1952 VDDD.n1951 9.3005
R4065 VDDD.n1950 VDDD.n1928 9.3005
R4066 VDDD.n1949 VDDD.n1948 9.3005
R4067 VDDD.n1947 VDDD.n1929 9.3005
R4068 VDDD.n1945 VDDD.n1944 9.3005
R4069 VDDD.n1943 VDDD.n1930 9.3005
R4070 VDDD.n2362 VDDD.n1888 9.3005
R4071 VDDD.n2365 VDDD.n2364 9.3005
R4072 VDDD.n2367 VDDD.n2366 9.3005
R4073 VDDD.n2369 VDDD.n1884 9.3005
R4074 VDDD.n2372 VDDD.n2371 9.3005
R4075 VDDD.n2387 VDDD.n2386 9.3005
R4076 VDDD.n2388 VDDD.n1671 9.3005
R4077 VDDD.n2389 VDDD.n1670 9.3005
R4078 VDDD.n2390 VDDD.n1669 9.3005
R4079 VDDD.n2394 VDDD.n2393 9.3005
R4080 VDDD.n2395 VDDD.n1668 9.3005
R4081 VDDD.n2397 VDDD.n2396 9.3005
R4082 VDDD.n2398 VDDD.n1666 9.3005
R4083 VDDD.n2401 VDDD.n2400 9.3005
R4084 VDDD.n2402 VDDD.n1665 9.3005
R4085 VDDD.n2404 VDDD.n2403 9.3005
R4086 VDDD.n2405 VDDD.n1664 9.3005
R4087 VDDD.n2410 VDDD.n2409 9.3005
R4088 VDDD.n2411 VDDD.n1663 9.3005
R4089 VDDD.n2413 VDDD.n2412 9.3005
R4090 VDDD.n2414 VDDD.n1658 9.3005
R4091 VDDD.n2415 VDDD.n2414 9.3005
R4092 VDDD.n2417 VDDD.n2416 9.3005
R4093 VDDD.n2418 VDDD.n1654 9.3005
R4094 VDDD.n2421 VDDD.n2420 9.3005
R4095 VDDD.n2490 VDDD.n2489 9.3005
R4096 VDDD.n2491 VDDD.n1648 9.3005
R4097 VDDD.n2481 VDDD.n1647 9.3005
R4098 VDDD.n2480 VDDD.n2479 9.3005
R4099 VDDD.n2476 VDDD.n2428 9.3005
R4100 VDDD.n2474 VDDD.n2473 9.3005
R4101 VDDD.n2472 VDDD.n2471 9.3005
R4102 VDDD.n2469 VDDD.n2431 9.3005
R4103 VDDD.n2468 VDDD.n2467 9.3005
R4104 VDDD.n2466 VDDD.n2432 9.3005
R4105 VDDD.n2465 VDDD.n2464 9.3005
R4106 VDDD.n2462 VDDD.n2434 9.3005
R4107 VDDD.n2460 VDDD.n2459 9.3005
R4108 VDDD.n2458 VDDD.n2457 9.3005
R4109 VDDD.n2455 VDDD.n2436 9.3005
R4110 VDDD.n2452 VDDD.n2451 9.3005
R4111 VDDD.n2450 VDDD.n2438 9.3005
R4112 VDDD.n2449 VDDD.n2448 9.3005
R4113 VDDD.n2446 VDDD.n2439 9.3005
R4114 VDDD.n2445 VDDD.n2444 9.3005
R4115 VDDD.n2443 VDDD.n2442 9.3005
R4116 VDDD.n1639 VDDD.n1637 9.3005
R4117 VDDD.n2577 VDDD.n2576 9.3005
R4118 VDDD.n2574 VDDD.n2573 9.3005
R4119 VDDD.n2566 VDDD.n1641 9.3005
R4120 VDDD.n2565 VDDD.n2564 9.3005
R4121 VDDD.n2562 VDDD.n1643 9.3005
R4122 VDDD.n2561 VDDD.n2560 9.3005
R4123 VDDD.n2559 VDDD.n2558 9.3005
R4124 VDDD.n2556 VDDD.n1646 9.3005
R4125 VDDD.n2556 VDDD.n1645 9.3005
R4126 VDDD.n2555 VDDD.n2554 9.3005
R4127 VDDD.n2553 VDDD.n2552 9.3005
R4128 VDDD.n2551 VDDD.n2495 9.3005
R4129 VDDD.n2550 VDDD.n2549 9.3005
R4130 VDDD.n2548 VDDD.n2547 9.3005
R4131 VDDD.n2546 VDDD.n2497 9.3005
R4132 VDDD.n2545 VDDD.n2544 9.3005
R4133 VDDD.n2543 VDDD.n2498 9.3005
R4134 VDDD.n2542 VDDD.n2541 9.3005
R4135 VDDD.n2540 VDDD.n2499 9.3005
R4136 VDDD.n2539 VDDD.n2538 9.3005
R4137 VDDD.n2537 VDDD.n2536 9.3005
R4138 VDDD.n2535 VDDD.n2534 9.3005
R4139 VDDD.n2533 VDDD.n2532 9.3005
R4140 VDDD.n2531 VDDD.n2502 9.3005
R4141 VDDD.n2530 VDDD.n2529 9.3005
R4142 VDDD.n2528 VDDD.n2527 9.3005
R4143 VDDD.n2526 VDDD.n2504 9.3005
R4144 VDDD.n2525 VDDD.n2524 9.3005
R4145 VDDD.n2523 VDDD.n2505 9.3005
R4146 VDDD.n2522 VDDD.n2521 9.3005
R4147 VDDD.n2520 VDDD.n2506 9.3005
R4148 VDDD.n2519 VDDD.n2518 9.3005
R4149 VDDD.n2517 VDDD.n2516 9.3005
R4150 VDDD.n1995 VDDD.n1981 9.3005
R4151 VDDD.n2020 VDDD.n2019 9.3005
R4152 VDDD.n2017 VDDD.n2016 9.3005
R4153 VDDD.n2013 VDDD.n1996 9.3005
R4154 VDDD.n2012 VDDD.n2011 9.3005
R4155 VDDD.n2010 VDDD.n2009 9.3005
R4156 VDDD.n2007 VDDD.n1999 9.3005
R4157 VDDD.n2006 VDDD.n2005 9.3005
R4158 VDDD.n2004 VDDD.n2003 9.3005
R4159 VDDD.n2001 VDDD.n1963 9.3005
R4160 VDDD.n2000 VDDD.n1964 9.3005
R4161 VDDD.n2324 VDDD.n2323 9.3005
R4162 VDDD.n2322 VDDD.n2321 9.3005
R4163 VDDD.n2320 VDDD.n2319 9.3005
R4164 VDDD.n2318 VDDD.n2317 9.3005
R4165 VDDD.n2316 VDDD.n2315 9.3005
R4166 VDDD.n2313 VDDD.n1971 9.3005
R4167 VDDD.n2312 VDDD.n2311 9.3005
R4168 VDDD.n2310 VDDD.n2309 9.3005
R4169 VDDD.n2307 VDDD.n1973 9.3005
R4170 VDDD.n2306 VDDD.n2305 9.3005
R4171 VDDD.n2304 VDDD.n1975 9.3005
R4172 VDDD.n2303 VDDD.n2302 9.3005
R4173 VDDD.n2300 VDDD.n1976 9.3005
R4174 VDDD.n2299 VDDD.n2298 9.3005
R4175 VDDD.n2297 VDDD.n2296 9.3005
R4176 VDDD.n2295 VDDD.n1979 9.3005
R4177 VDDD.n2081 VDDD.n1980 9.3005
R4178 VDDD.n2082 VDDD.n2074 9.3005
R4179 VDDD.n2084 VDDD.n2083 9.3005
R4180 VDDD.n2091 VDDD.n2090 9.3005
R4181 VDDD.n2093 VDDD.n2069 9.3005
R4182 VDDD.n2106 VDDD.n2105 9.3005
R4183 VDDD.n2110 VDDD.n2109 9.3005
R4184 VDDD.n2111 VDDD.n2067 9.3005
R4185 VDDD.n2113 VDDD.n2112 9.3005
R4186 VDDD.n2114 VDDD.n2066 9.3005
R4187 VDDD.n2116 VDDD.n2115 9.3005
R4188 VDDD.n2118 VDDD.n2117 9.3005
R4189 VDDD.n2119 VDDD.n2063 9.3005
R4190 VDDD.n2122 VDDD.n2121 9.3005
R4191 VDDD.n2124 VDDD.n2123 9.3005
R4192 VDDD.n2126 VDDD.n2125 9.3005
R4193 VDDD.n2128 VDDD.n2127 9.3005
R4194 VDDD.n2130 VDDD.n2059 9.3005
R4195 VDDD.n2133 VDDD.n2132 9.3005
R4196 VDDD.n2135 VDDD.n2134 9.3005
R4197 VDDD.n2136 VDDD.n2057 9.3005
R4198 VDDD.n2139 VDDD.n2138 9.3005
R4199 VDDD.n2141 VDDD.n2140 9.3005
R4200 VDDD.n2144 VDDD.n2143 9.3005
R4201 VDDD.n2146 VDDD.n2145 9.3005
R4202 VDDD.n2147 VDDD.n2049 9.3005
R4203 VDDD.n2150 VDDD.n2149 9.3005
R4204 VDDD.n2050 VDDD.n2022 9.3005
R4205 VDDD.n2163 VDDD.n2159 9.3005
R4206 VDDD.n2166 VDDD.n2165 9.3005
R4207 VDDD.n2168 VDDD.n2167 9.3005
R4208 VDDD.n2169 VDDD.n2040 9.3005
R4209 VDDD.n2172 VDDD.n2171 9.3005
R4210 VDDD.n2173 VDDD.n2039 9.3005
R4211 VDDD.n2175 VDDD.n2174 9.3005
R4212 VDDD.n2177 VDDD.n2037 9.3005
R4213 VDDD.n2179 VDDD.n2178 9.3005
R4214 VDDD.n2181 VDDD.n2180 9.3005
R4215 VDDD.n2182 VDDD.n2035 9.3005
R4216 VDDD.n2184 VDDD.n2183 9.3005
R4217 VDDD.n2186 VDDD.n2185 9.3005
R4218 VDDD.n2189 VDDD.n2033 9.3005
R4219 VDDD.n2193 VDDD.n2192 9.3005
R4220 VDDD.n2194 VDDD.n2032 9.3005
R4221 VDDD.n2196 VDDD.n2195 9.3005
R4222 VDDD.n2201 VDDD.n2200 9.3005
R4223 VDDD.n2204 VDDD.n2028 9.3005
R4224 VDDD.n2216 VDDD.n2215 9.3005
R4225 VDDD.n2220 VDDD.n2219 9.3005
R4226 VDDD.n2221 VDDD.n2026 9.3005
R4227 VDDD.n2223 VDDD.n2222 9.3005
R4228 VDDD.n2224 VDDD.n2025 9.3005
R4229 VDDD.n2227 VDDD.n2226 9.3005
R4230 VDDD.n2291 VDDD.n2228 9.3005
R4231 VDDD.n2291 VDDD.n2024 9.3005
R4232 VDDD.n2290 VDDD.n2289 9.3005
R4233 VDDD.n2288 VDDD.n2287 9.3005
R4234 VDDD.n2286 VDDD.n2230 9.3005
R4235 VDDD.n2285 VDDD.n2284 9.3005
R4236 VDDD.n2283 VDDD.n2282 9.3005
R4237 VDDD.n2281 VDDD.n2232 9.3005
R4238 VDDD.n2280 VDDD.n2279 9.3005
R4239 VDDD.n2278 VDDD.n2233 9.3005
R4240 VDDD.n2277 VDDD.n2276 9.3005
R4241 VDDD.n2275 VDDD.n2234 9.3005
R4242 VDDD.n2274 VDDD.n2273 9.3005
R4243 VDDD.n2272 VDDD.n2271 9.3005
R4244 VDDD.n2270 VDDD.n2269 9.3005
R4245 VDDD.n2268 VDDD.n2267 9.3005
R4246 VDDD.n2266 VDDD.n2237 9.3005
R4247 VDDD.n2265 VDDD.n2264 9.3005
R4248 VDDD.n2263 VDDD.n2262 9.3005
R4249 VDDD.n2261 VDDD.n2239 9.3005
R4250 VDDD.n2260 VDDD.n2259 9.3005
R4251 VDDD.n2258 VDDD.n2240 9.3005
R4252 VDDD.n2257 VDDD.n2256 9.3005
R4253 VDDD.n2255 VDDD.n2241 9.3005
R4254 VDDD.n2254 VDDD.n2253 9.3005
R4255 VDDD.n2252 VDDD.n2251 9.3005
R4256 VDDD.n135 VDDD.n134 9.3005
R4257 VDDD.n136 VDDD.n130 9.3005
R4258 VDDD.n138 VDDD.n137 9.3005
R4259 VDDD.n139 VDDD.n128 9.3005
R4260 VDDD.n140 VDDD.n127 9.3005
R4261 VDDD.n144 VDDD.n143 9.3005
R4262 VDDD.n146 VDDD.n145 9.3005
R4263 VDDD.n148 VDDD.n147 9.3005
R4264 VDDD.n150 VDDD.n149 9.3005
R4265 VDDD.n151 VDDD.n124 9.3005
R4266 VDDD.n153 VDDD.n152 9.3005
R4267 VDDD.n155 VDDD.n154 9.3005
R4268 VDDD.n156 VDDD.n122 9.3005
R4269 VDDD.n158 VDDD.n157 9.3005
R4270 VDDD.n159 VDDD.n120 9.3005
R4271 VDDD.n170 VDDD.n169 9.3005
R4272 VDDD.n171 VDDD.n118 9.3005
R4273 VDDD.n201 VDDD.n200 9.3005
R4274 VDDD.n198 VDDD.n119 9.3005
R4275 VDDD.n197 VDDD.n196 9.3005
R4276 VDDD.n195 VDDD.n194 9.3005
R4277 VDDD.n193 VDDD.n173 9.3005
R4278 VDDD.n192 VDDD.n191 9.3005
R4279 VDDD.n190 VDDD.n189 9.3005
R4280 VDDD.n188 VDDD.n175 9.3005
R4281 VDDD.n187 VDDD.n186 9.3005
R4282 VDDD.n185 VDDD.n176 9.3005
R4283 VDDD.n184 VDDD.n183 9.3005
R4284 VDDD.n182 VDDD.n177 9.3005
R4285 VDDD.n181 VDDD.n180 9.3005
R4286 VDDD.n179 VDDD.n48 9.3005
R4287 VDDD.n3706 VDDD.n3705 9.3005
R4288 VDDD.n3704 VDDD.n47 9.3005
R4289 VDDD.n3703 VDDD.n3702 9.3005
R4290 VDDD.n3700 VDDD.n49 9.3005
R4291 VDDD.n3699 VDDD.n3698 9.3005
R4292 VDDD.n61 VDDD.n60 9.3005
R4293 VDDD.n67 VDDD.n66 9.3005
R4294 VDDD.n109 VDDD.n108 9.3005
R4295 VDDD.n106 VDDD.n59 9.3005
R4296 VDDD.n105 VDDD.n104 9.3005
R4297 VDDD.n103 VDDD.n68 9.3005
R4298 VDDD.n102 VDDD.n101 9.3005
R4299 VDDD.n100 VDDD.n69 9.3005
R4300 VDDD.n99 VDDD.n98 9.3005
R4301 VDDD.n97 VDDD.n70 9.3005
R4302 VDDD.n96 VDDD.n95 9.3005
R4303 VDDD.n94 VDDD.n93 9.3005
R4304 VDDD.n92 VDDD.n91 9.3005
R4305 VDDD.n90 VDDD.n73 9.3005
R4306 VDDD.n89 VDDD.n88 9.3005
R4307 VDDD.n87 VDDD.n86 9.3005
R4308 VDDD.n85 VDDD.n75 9.3005
R4309 VDDD.n84 VDDD.n83 9.3005
R4310 VDDD.n82 VDDD.n76 9.3005
R4311 VDDD.n81 VDDD.n80 9.3005
R4312 VDDD.n79 VDDD.n77 9.3005
R4313 VDDD.n78 VDDD.n45 9.3005
R4314 VDDD.n3717 VDDD.n3716 9.3005
R4315 VDDD.n3715 VDDD.n3714 9.3005
R4316 VDDD.n3726 VDDD.n38 9.3005
R4317 VDDD.n3728 VDDD.n3727 9.3005
R4318 VDDD.n3731 VDDD.n37 9.3005
R4319 VDDD.n3733 VDDD.n3732 9.3005
R4320 VDDD.n3735 VDDD.n3734 9.3005
R4321 VDDD.n3736 VDDD.n35 9.3005
R4322 VDDD.n3738 VDDD.n3737 9.3005
R4323 VDDD.n3739 VDDD.n34 9.3005
R4324 VDDD.n3741 VDDD.n3740 9.3005
R4325 VDDD.n3743 VDDD.n32 9.3005
R4326 VDDD.n3745 VDDD.n3744 9.3005
R4327 VDDD.n3746 VDDD.n31 9.3005
R4328 VDDD.n3748 VDDD.n3747 9.3005
R4329 VDDD.n3749 VDDD.n30 9.3005
R4330 VDDD.n3751 VDDD.n3750 9.3005
R4331 VDDD.n3752 VDDD.n29 9.3005
R4332 VDDD.n3754 VDDD.n3753 9.3005
R4333 VDDD.n3756 VDDD.n27 9.3005
R4334 VDDD.n3758 VDDD.n3757 9.3005
R4335 VDDD.n3759 VDDD.n20 9.3005
R4336 VDDD.n3773 VDDD.n3772 9.3005
R4337 VDDD.n3774 VDDD.n19 9.3005
R4338 VDDD.n3775 VDDD.n18 9.3005
R4339 VDDD.n3777 VDDD.n3776 9.3005
R4340 VDDD.n3778 VDDD.n17 9.3005
R4341 VDDD.n3780 VDDD.n3779 9.3005
R4342 VDDD.n3782 VDDD.n3781 9.3005
R4343 VDDD.n3783 VDDD.n15 9.3005
R4344 VDDD.n3785 VDDD.n3784 9.3005
R4345 VDDD.n3787 VDDD.n3786 9.3005
R4346 VDDD.n3789 VDDD.n3788 9.3005
R4347 VDDD.n3790 VDDD.n13 9.3005
R4348 VDDD.n3792 VDDD.n3791 9.3005
R4349 VDDD.n3794 VDDD.n3793 9.3005
R4350 VDDD.n3795 VDDD.n11 9.3005
R4351 VDDD.n3797 VDDD.n3796 9.3005
R4352 VDDD.n3798 VDDD.n10 9.3005
R4353 VDDD.n3800 VDDD.n3799 9.3005
R4354 VDDD.n3801 VDDD.n9 9.3005
R4355 VDDD.n3803 VDDD.n3802 9.3005
R4356 VDDD.n3805 VDDD.n3804 9.3005
R4357 VDDD.n3807 VDDD.n3806 9.3005
R4358 VDDD.n3809 VDDD.n3808 9.3005
R4359 VDDD.n3810 VDDD.n6 9.3005
R4360 VDDD.n3812 VDDD.n3811 9.3005
R4361 VDDD.n3814 VDDD.n3813 9.3005
R4362 VDDD.n3815 VDDD.n4 9.3005
R4363 VDDD.n3817 VDDD.n3816 9.3005
R4364 VDDD.n3818 VDDD.n3 9.3005
R4365 VDDD.n3820 VDDD.n3819 9.3005
R4366 VDDD.n3821 VDDD.n2 9.3005
R4367 VDDD.n3824 VDDD.n3823 9.3005
R4368 VDDD.n3825 VDDD.n1 9.3005
R4369 VDDD.n3827 VDDD.n3826 9.3005
R4370 VDDD.n3830 VDDD.n0 9.3005
R4371 VDDD.n3200 VDDD.n3199 9.20381
R4372 VDDD.n1225 VDDD.n1153 9.20381
R4373 VDDD.n2138 VDDD.n2137 9.20381
R4374 VDDD.n3809 VDDD.n7 9.09802
R4375 VDDD.n3823 VDDD.n3822 9.09802
R4376 VDDD.n3789 VDDD.n14 9.09802
R4377 VDDD.n3802 VDDD.n8 9.09802
R4378 VDDD.n3607 VDDD.n3605 9.09802
R4379 VDDD.n3615 VDDD.n3614 9.09802
R4380 VDDD.n3632 VDDD.n3631 9.09802
R4381 VDDD.n3638 VDDD.n334 9.09802
R4382 VDDD.n3663 VDDD.n3662 9.09802
R4383 VDDD.n3657 VDDD.n224 9.09802
R4384 VDDD.n3507 VDDD.n3504 9.09802
R4385 VDDD.n451 VDDD.n378 9.09802
R4386 VDDD.n3110 VDDD.n658 9.09802
R4387 VDDD.n3223 VDDD.n3222 9.09802
R4388 VDDD.n3215 VDDD.n3179 9.09802
R4389 VDDD.n3199 VDDD.n3187 9.09802
R4390 VDDD.n790 VDDD.n789 9.09802
R4391 VDDD.n3049 VDDD.n765 9.09802
R4392 VDDD.n2974 VDDD.n2973 9.09802
R4393 VDDD.n1225 VDDD.n1224 9.09802
R4394 VDDD.n1222 VDDD.n1156 9.09802
R4395 VDDD.n1844 VDDD.n1821 9.09802
R4396 VDDD.n1756 VDDD.n1728 9.09802
R4397 VDDD.n1781 VDDD.n1704 9.09802
R4398 VDDD.n1762 VDDD.n1761 9.09802
R4399 VDDD.n2447 VDDD.n2446 9.09802
R4400 VDDD.n2128 VDDD.n2061 9.09802
R4401 VDDD.n2138 VDDD.n2056 9.09802
R4402 VDDD.n2086 VDDD.n2069 9.09802
R4403 VDDD.n2121 VDDD.n2062 9.09802
R4404 VDDD.n2183 VDDD.n2034 9.09802
R4405 VDDD.n2192 VDDD.n2190 9.09802
R4406 VDDD.n2200 VDDD.n2199 9.09802
R4407 VDDD.n2322 VDDD.n1969 9.09802
R4408 VDDD.n2315 VDDD.n1970 9.09802
R4409 VDDD.n91 VDDD.n72 9.09802
R4410 VDDD.n78 VDDD.n46 9.09802
R4411 VDDD.n60 VDDD.n52 9.09802
R4412 VDDD.n71 VDDD.n70 9.09802
R4413 VDDD.n194 VDDD.n172 9.09802
R4414 VDDD.n181 VDDD.n178 9.09802
R4415 VDDD.n150 VDDD.n125 9.09802
R4416 VDDD.n200 VDDD.n199 9.09802
R4417 VDDD.n323 VDDD.n272 9.03579
R4418 VDDD.n3549 VDDD.n3548 9.03579
R4419 VDDD.n3365 VDDD.n3364 9.03579
R4420 VDDD.n3147 VDDD.n642 9.03579
R4421 VDDD.n715 VDDD.n714 9.03579
R4422 VDDD.n858 VDDD.n857 9.03579
R4423 VDDD.n1011 VDDD.n893 9.03579
R4424 VDDD.n931 VDDD.n929 9.03579
R4425 VDDD.n1461 VDDD.n1460 9.03579
R4426 VDDD.n2812 VDDD.n2810 9.03579
R4427 VDDD.n1855 VDDD.n1854 9.03579
R4428 VDDD.n2591 VDDD.n1576 9.03579
R4429 VDDD.n2387 VDDD.n1673 9.03579
R4430 VDDD.n3743 VDDD.n3742 9.03579
R4431 VDDD.n1740 VDDD.n1737 9.02345
R4432 VDDD.n3157 VDDD.n3156 8.9761
R4433 VDDD.n2700 VDDD.n2699 8.9761
R4434 VDDD.n542 VDDD.n511 8.81089
R4435 VDDD.n1411 VDDD.n1410 8.77764
R4436 VDDD.n1802 VDDD.n1801 8.77764
R4437 VDDD.n1865 VDDD.n1809 8.77764
R4438 VDDD.n605 VDDD.n604 8.65932
R4439 VDDD.n983 VDDD.n917 8.62646
R4440 VDDD.n1741 VDDD.n1740 8.49886
R4441 VDDD.t869 VDDD.n3646 8.39273
R4442 VDDD.t165 VDDD.n3645 8.39273
R4443 VDDD.t837 VDDD.t1243 8.39273
R4444 VDDD.t591 VDDD.t277 8.39273
R4445 VDDD.t391 VDDD.t599 8.39273
R4446 VDDD.t1318 VDDD.t265 8.39273
R4447 VDDD.n3676 VDDD.n216 8.35752
R4448 VDDD.n427 VDDD.n389 8.35752
R4449 VDDD.n3208 VDDD.n3207 8.35752
R4450 VDDD.n3062 VDDD.n758 8.35752
R4451 VDDD.n2129 VDDD.n2128 8.35752
R4452 VDDD.n2009 VDDD.n1998 8.35752
R4453 VDDD.n2878 VDDD.n2875 8.28285
R4454 VDDD.n2621 VDDD.n2618 8.28285
R4455 VDDD.n3436 VDDD.n3435 8.18368
R4456 VDDD.n1743 VDDD.n1735 8.04017
R4457 VDDD.n2564 VDDD.n1641 7.75995
R4458 VDDD.n2143 VDDD.n2141 7.75995
R4459 VDDD.n2216 VDDD.n2028 7.75995
R4460 VDDD.n2306 VDDD.n1975 7.75995
R4461 VDDD.n3656 VDDD.n3655 7.72281
R4462 VDDD.n729 VDDD.n721 7.72281
R4463 VDDD.n3230 VDDD.n3229 7.72281
R4464 VDDD.n1754 VDDD.n1753 7.72281
R4465 VDDD.n2442 VDDD.n2440 7.72281
R4466 VDDD.n2107 VDDD.n2106 7.72281
R4467 VDDD.n2314 VDDD.n2313 7.72281
R4468 VDDD.n3139 VDDD.n3138 7.52991
R4469 VDDD.n2699 VDDD.n2698 7.39867
R4470 VDDD.n305 VDDD.n282 7.15344
R4471 VDDD.n3548 VDDD.n3547 7.15344
R4472 VDDD.n714 VDDD.n711 7.15344
R4473 VDDD.n610 VDDD.n609 7.15344
R4474 VDDD.n857 VDDD.n854 7.15344
R4475 VDDD.n872 VDDD.n861 7.15344
R4476 VDDD.n958 VDDD.n957 7.15344
R4477 VDDD.n2989 VDDD.n1127 7.15344
R4478 VDDD.n2825 VDDD.n2824 7.15344
R4479 VDDD.n2859 VDDD.n1251 7.15344
R4480 VDDD.n2164 VDDD.n2041 7.0881
R4481 VDDD.n3130 VDDD.n3129 6.77697
R4482 VDDD.n3039 VDDD.n771 6.77697
R4483 VDDD.n829 VDDD.n820 6.77697
R4484 VDDD.n2764 VDDD.n1274 6.77697
R4485 VDDD.n2721 VDDD.n2720 6.77697
R4486 VDDD.n2342 VDDD.n1906 6.77697
R4487 VDDD.n3155 VDDD.n3154 6.73838
R4488 VDDD.n3248 VDDD.n3172 6.73838
R4489 VDDD.t584 VDDD 6.71428
R4490 VDDD VDDD.t619 6.71428
R4491 VDDD.t1357 VDDD 6.71428
R4492 VDDD.n3290 VDDD.n3288 6.67526
R4493 VDDD.n3237 VDDD.n3173 6.66496
R4494 VDDD.n1834 VDDD.n1833 6.66496
R4495 VDDD.n530 VDDD.n529 6.58769
R4496 VDDD.n3669 VDDD.n3668 6.55918
R4497 VDDD.n430 VDDD.n381 6.55918
R4498 VDDD.n3215 VDDD.n3214 6.55918
R4499 VDDD.n3056 VDDD.n3055 6.55918
R4500 VDDD.n1725 VDDD.n1719 6.55918
R4501 VDDD.n2120 VDDD.n2119 6.55918
R4502 VDDD.n2178 VDDD.n2036 6.55918
R4503 VDDD.n2002 VDDD.n2001 6.55918
R4504 VDDD.n1940 VDDD.n1939 6.46951
R4505 VDDD.n2557 VDDD.n2556 6.46951
R4506 VDDD.n2291 VDDD.n2023 6.46951
R4507 VDDD.n3536 VDDD.n3535 6.4005
R4508 VDDD.n697 VDDD.n689 6.4005
R4509 VDDD.n1069 VDDD.n847 6.4005
R4510 VDDD.n882 VDDD.n879 6.4005
R4511 VDDD.n965 VDDD.n964 6.4005
R4512 VDDD.n2832 VDDD.n2831 6.4005
R4513 VDDD.n2934 VDDD.n2863 6.4005
R4514 VDDD.n2692 VDDD.n1569 6.4005
R4515 VDDD.n1609 VDDD.n1608 6.4005
R4516 VDDD.n2672 VDDD.n2606 6.4005
R4517 VDDD.n2408 VDDD.n2407 6.4005
R4518 VDDD.n1863 VDDD.n1862 6.21764
R4519 VDDD.n3607 VDDD.n3606 6.03025
R4520 VDDD.n3638 VDDD.n3637 6.03025
R4521 VDDD.n240 VDDD.n239 6.03025
R4522 VDDD.n423 VDDD.n422 6.03025
R4523 VDDD.n3186 VDDD.n3184 6.03025
R4524 VDDD.n1231 VDDD.n1230 6.03025
R4525 VDDD.n1780 VDDD.n1779 6.03025
R4526 VDDD.n2192 VDDD.n2191 6.03025
R4527 VDDD.n2014 VDDD.n2013 6.03025
R4528 VDDD.n355 VDDD.n352 6.02403
R4529 VDDD.n3591 VDDD.n3590 6.02403
R4530 VDDD.n3541 VDDD.n3491 6.02403
R4531 VDDD.n3380 VDDD.n3336 6.02403
R4532 VDDD.n3380 VDDD.n3379 6.02403
R4533 VDDD.n743 VDDD.n709 6.02403
R4534 VDDD.n1064 VDDD.n851 6.02403
R4535 VDDD.n1022 VDDD.n1021 6.02403
R4536 VDDD.n970 VDDD.n926 6.02403
R4537 VDDD.n2808 VDDD.n2805 6.02403
R4538 VDDD.n2772 VDDD.n2771 6.02403
R4539 VDDD.n2770 VDDD.n2769 6.02403
R4540 VDDD.n1524 VDDD.n1315 6.02403
R4541 VDDD.n1527 VDDD.n1526 6.02403
R4542 VDDD.n2869 VDDD.n2866 6.02403
R4543 VDDD.n1616 VDDD.n1591 6.02403
R4544 VDDD.n2612 VDDD.n2609 6.02403
R4545 VDDD.n1927 VDDD.n1926 6.02403
R4546 VDDD.n1925 VDDD.n1917 6.02403
R4547 VDDD.n2400 VDDD.n2399 6.02403
R4548 VDDD.n3756 VDDD.n3755 6.02403
R4549 VDDD.n1410 VDDD.n1408 5.85193
R4550 VDDD.n1215 VDDD.n1214 5.66204
R4551 VDDD.n1214 VDDD.n1213 5.66204
R4552 VDDD.n1210 VDDD.n1209 5.66204
R4553 VDDD.n1209 VDDD.n1208 5.66204
R4554 VDDD.n1208 VDDD.n1161 5.66204
R4555 VDDD.n1204 VDDD.n1161 5.66204
R4556 VDDD.n1204 VDDD.n1203 5.66204
R4557 VDDD.n1203 VDDD.n1202 5.66204
R4558 VDDD.n1195 VDDD.n1194 5.66204
R4559 VDDD.n1194 VDDD.n1193 5.66204
R4560 VDDD.n1190 VDDD.n1189 5.66204
R4561 VDDD.n1189 VDDD.n1188 5.66204
R4562 VDDD.n1188 VDDD.n1168 5.66204
R4563 VDDD.n1184 VDDD.n1168 5.66204
R4564 VDDD.n1184 VDDD.n1183 5.66204
R4565 VDDD.n1183 VDDD.n1182 5.66204
R4566 VDDD.n2552 VDDD.n2551 5.66204
R4567 VDDD.n2551 VDDD.n2550 5.66204
R4568 VDDD.n2547 VDDD.n2546 5.66204
R4569 VDDD.n2546 VDDD.n2545 5.66204
R4570 VDDD.n2545 VDDD.n2498 5.66204
R4571 VDDD.n2541 VDDD.n2498 5.66204
R4572 VDDD.n2541 VDDD.n2540 5.66204
R4573 VDDD.n2540 VDDD.n2539 5.66204
R4574 VDDD.n2532 VDDD.n2531 5.66204
R4575 VDDD.n2531 VDDD.n2530 5.66204
R4576 VDDD.n2527 VDDD.n2526 5.66204
R4577 VDDD.n2526 VDDD.n2525 5.66204
R4578 VDDD.n2525 VDDD.n2505 5.66204
R4579 VDDD.n2521 VDDD.n2505 5.66204
R4580 VDDD.n2521 VDDD.n2520 5.66204
R4581 VDDD.n2520 VDDD.n2519 5.66204
R4582 VDDD.n2287 VDDD.n2286 5.66204
R4583 VDDD.n2286 VDDD.n2285 5.66204
R4584 VDDD.n2282 VDDD.n2281 5.66204
R4585 VDDD.n2281 VDDD.n2280 5.66204
R4586 VDDD.n2280 VDDD.n2233 5.66204
R4587 VDDD.n2276 VDDD.n2233 5.66204
R4588 VDDD.n2276 VDDD.n2275 5.66204
R4589 VDDD.n2275 VDDD.n2274 5.66204
R4590 VDDD.n2267 VDDD.n2266 5.66204
R4591 VDDD.n2266 VDDD.n2265 5.66204
R4592 VDDD.n2262 VDDD.n2261 5.66204
R4593 VDDD.n2261 VDDD.n2260 5.66204
R4594 VDDD.n2260 VDDD.n2240 5.66204
R4595 VDDD.n2256 VDDD.n2240 5.66204
R4596 VDDD.n2256 VDDD.n2255 5.66204
R4597 VDDD.n2255 VDDD.n2254 5.66204
R4598 VDDD.n2945 VDDD.n1247 5.40233
R4599 VDDD.n2885 VDDD.n2884 5.40233
R4600 VDDD.n3511 VDDD.n3510 5.39554
R4601 VDDD.n3241 VDDD.n3240 5.3712
R4602 VDDD.n1215 VDDD.n1157 5.29281
R4603 VDDD.n1202 VDDD.n1163 5.29281
R4604 VDDD.n1195 VDDD.n1164 5.29281
R4605 VDDD.n1182 VDDD.n1170 5.29281
R4606 VDDD.n2552 VDDD.n2494 5.29281
R4607 VDDD.n2539 VDDD.n2500 5.29281
R4608 VDDD.n2532 VDDD.n2501 5.29281
R4609 VDDD.n2519 VDDD.n2507 5.29281
R4610 VDDD.n2287 VDDD.n2229 5.29281
R4611 VDDD.n2274 VDDD.n2235 5.29281
R4612 VDDD.n2267 VDDD.n2236 5.29281
R4613 VDDD.n2254 VDDD.n2242 5.29281
R4614 VDDD.n397 VDDD.n396 5.28746
R4615 VDDD.n684 VDDD.n683 5.27109
R4616 VDDD.n394 VDDD.n393 5.23129
R4617 VDDD.n3811 VDDD.n5 5.18397
R4618 VDDD.n3791 VDDD.n12 5.18397
R4619 VDDD.n3676 VDDD.n3675 5.18397
R4620 VDDD.n3664 VDDD.n220 5.18397
R4621 VDDD.n3654 VDDD.n225 5.18397
R4622 VDDD.n428 VDDD.n427 5.18397
R4623 VDDD.n450 VDDD.n449 5.18397
R4624 VDDD.n3237 VDDD.n3236 5.18397
R4625 VDDD.n3212 VDDD.n3181 5.18397
R4626 VDDD.n3061 VDDD.n759 5.18397
R4627 VDDD.n3051 VDDD.n764 5.18397
R4628 VDDD.n1150 VDDD.n1136 5.18397
R4629 VDDD.n1753 VDDD.n1730 5.18397
R4630 VDDD.n1762 VDDD.n1727 5.18397
R4631 VDDD.n2442 VDDD.n2441 5.18397
R4632 VDDD.n2132 VDDD.n2131 5.18397
R4633 VDDD.n2109 VDDD.n2108 5.18397
R4634 VDDD.n2115 VDDD.n2065 5.18397
R4635 VDDD.n2171 VDDD.n2170 5.18397
R4636 VDDD.n2176 VDDD.n2175 5.18397
R4637 VDDD.n2009 VDDD.n2008 5.18397
R4638 VDDD.n2323 VDDD.n1968 5.18397
R4639 VDDD.n2312 VDDD.n1972 5.18397
R4640 VDDD.n89 VDDD.n74 5.18397
R4641 VDDD.n108 VDDD.n107 5.18397
R4642 VDDD.n192 VDDD.n174 5.18397
R4643 VDDD.n152 VDDD.n123 5.18397
R4644 VDDD.n257 VDDD.n256 5.05557
R4645 VDDD.n505 VDDD.n500 5.03517
R4646 VDDD.n2077 VDDD.n2076 5.03517
R4647 VDDD.n3169 VDDD.n622 4.98336
R4648 VDDD.n724 VDDD.n723 4.9724
R4649 VDDD.n3447 VDDD.n3446 4.91363
R4650 VDDD.n3558 VDDD.n3557 4.89462
R4651 VDDD.n3537 VDDD.n3536 4.89462
R4652 VDDD.n3367 VDDD.n3341 4.89462
R4653 VDDD.n3392 VDDD.n3391 4.89462
R4654 VDDD.n456 VDDD.n376 4.89462
R4655 VDDD.n706 VDDD.n697 4.89462
R4656 VDDD.n1069 VDDD.n1068 4.89462
R4657 VDDD.n1001 VDDD.n907 4.89462
R4658 VDDD.n964 VDDD.n963 4.89462
R4659 VDDD.n2831 VDDD.n2830 4.89462
R4660 VDDD.n2925 VDDD.n2924 4.89462
R4661 VDDD.n2913 VDDD.n2878 4.89462
R4662 VDDD.n2596 VDDD.n2595 4.89462
R4663 VDDD.n2663 VDDD.n2662 4.89462
R4664 VDDD.n2651 VDDD.n2621 4.89462
R4665 VDDD.n2370 VDDD.n2369 4.89462
R4666 VDDD.n1377 VDDD.n1373 4.75479
R4667 VDDD.n1864 VDDD.n1863 4.75479
R4668 VDDD.n553 VDDD.n552 4.67352
R4669 VDDD.n3441 VDDD.n3440 4.67352
R4670 VDDD.n3440 VDDD.n3439 4.67352
R4671 VDDD.n3406 VDDD.n3405 4.67352
R4672 VDDD.n475 VDDD.n472 4.67352
R4673 VDDD.n3152 VDDD.n636 4.67352
R4674 VDDD.n3154 VDDD.n3152 4.67352
R4675 VDDD.n3095 VDDD.n3094 4.67352
R4676 VDDD.n615 VDDD.n581 4.67352
R4677 VDDD.n3255 VDDD.n3254 4.67352
R4678 VDDD.n3249 VDDD.n3248 4.67352
R4679 VDDD.n1038 VDDD.n1037 4.67352
R4680 VDDD.n986 VDDD.n985 4.67352
R4681 VDDD.n1473 VDDD.n1472 4.67352
R4682 VDDD.n1490 VDDD.n1489 4.67352
R4683 VDDD.n3002 VDDD.n3001 4.67352
R4684 VDDD.n2956 VDDD.n1244 4.67352
R4685 VDDD.n2946 VDDD.n1244 4.67352
R4686 VDDD.n2944 VDDD.n2943 4.67352
R4687 VDDD.n2787 VDDD.n1259 4.67352
R4688 VDDD.n2791 VDDD.n1259 4.67352
R4689 VDDD.n2901 VDDD.n2900 4.67352
R4690 VDDD.n2900 VDDD.n2882 4.67352
R4691 VDDD.n1790 VDDD.n1701 4.67352
R4692 VDDD.n2639 VDDD.n2638 4.67352
R4693 VDDD.n2418 VDDD.n2417 4.67352
R4694 VDDD.n2295 VDDD.n1980 4.67352
R4695 VDDD.n3732 VDDD.n3731 4.67352
R4696 VDDD.n3613 VDDD.n3612 4.65505
R4697 VDDD.n539 VDDD.n513 4.65505
R4698 VDDD.n2198 VDDD.n2197 4.65505
R4699 VDDD.n1397 VDDD.n1374 4.62124
R4700 VDDD.n1941 VDDD.n1940 4.62124
R4701 VDDD.n2163 VDDD.n2043 4.62124
R4702 VDDD.n3446 VDDD.n3295 4.62124
R4703 VDDD.n3169 VDDD.n576 4.62124
R4704 VDDD.n809 VDDD.n781 4.62124
R4705 VDDD.n1832 VDDD.n1830 4.62124
R4706 VDDD.n2414 VDDD.n1659 4.62124
R4707 VDDD.n554 VDDD.n553 4.57193
R4708 VDDD.n617 VDDD.n616 4.57193
R4709 VDDD.n1039 VDDD.n1038 4.57193
R4710 VDDD.n1037 VDDD.n877 4.57193
R4711 VDDD.n1488 VDDD.n1487 4.57193
R4712 VDDD.n2792 VDDD.n2791 4.57193
R4713 VDDD.n1601 VDDD.n1600 4.57193
R4714 VDDD.n3814 VDDD.n5 4.54926
R4715 VDDD.n3794 VDDD.n12 4.54926
R4716 VDDD.n3615 VDDD.n3613 4.54926
R4717 VDDD.n3675 VDDD.n3674 4.54926
R4718 VDDD.n3667 VDDD.n220 4.54926
R4719 VDDD.n3651 VDDD.n225 4.54926
R4720 VDDD.n429 VDDD.n428 4.54926
R4721 VDDD.n449 VDDD.n448 4.54926
R4722 VDDD.n723 VDDD.n667 4.54926
R4723 VDDD.n3209 VDDD.n3181 4.54926
R4724 VDDD.n3058 VDDD.n759 4.54926
R4725 VDDD.n764 VDDD.n761 4.54926
R4726 VDDD.n1839 VDDD.n1824 4.54926
R4727 VDDD.n1750 VDDD.n1730 4.54926
R4728 VDDD.n1775 VDDD.n1709 4.54926
R4729 VDDD.n1727 VDDD.n1726 4.54926
R4730 VDDD.n2441 VDDD.n1639 4.54926
R4731 VDDD.n2108 VDDD.n2067 4.54926
R4732 VDDD.n2118 VDDD.n2065 4.54926
R4733 VDDD.n2170 VDDD.n2039 4.54926
R4734 VDDD.n2177 VDDD.n2176 4.54926
R4735 VDDD.n2200 VDDD.n2198 4.54926
R4736 VDDD.n2008 VDDD.n2007 4.54926
R4737 VDDD.n2000 VDDD.n1968 4.54926
R4738 VDDD.n2309 VDDD.n1972 4.54926
R4739 VDDD.n86 VDDD.n74 4.54926
R4740 VDDD.n107 VDDD.n106 4.54926
R4741 VDDD.n189 VDDD.n174 4.54926
R4742 VDDD.n155 VDDD.n123 4.54926
R4743 VDDD.n2751 VDDD.n2750 4.51815
R4744 VDDD.n2728 VDDD.n2727 4.51815
R4745 VDDD.n2350 VDDD.n2349 4.51815
R4746 VDDD.n3697 VDDD.n3696 4.51401
R4747 VDDD.n111 VDDD.n110 4.51401
R4748 VDDD.n3720 VDDD.n43 4.51401
R4749 VDDD.n3725 VDDD.n3724 4.51401
R4750 VDDD.n3762 VDDD.n3760 4.51401
R4751 VDDD.n3766 VDDD.n3765 4.51401
R4752 VDDD.n3572 VDDD.n3473 4.51401
R4753 VDDD.n3577 VDDD.n3576 4.51401
R4754 VDDD.n3518 VDDD.n3514 4.51401
R4755 VDDD.n3523 VDDD.n3496 4.51401
R4756 VDDD.n3686 VDDD.n209 4.51401
R4757 VDDD.n214 VDDD.n213 4.51401
R4758 VDDD.n3622 VDDD.n343 4.51401
R4759 VDDD.n3626 VDDD.n337 4.51401
R4760 VDDD.n3469 VDDD.n364 4.51401
R4761 VDDD.n3460 VDDD.n3459 4.51401
R4762 VDDD.n3285 VDDD.n3284 4.51401
R4763 VDDD.n559 VDDD.n558 4.51401
R4764 VDDD.n436 VDDD.n434 4.51401
R4765 VDDD.n446 VDDD.n445 4.51401
R4766 VDDD.n3318 VDDD.n3310 4.51401
R4767 VDDD.n3411 VDDD.n3410 4.51401
R4768 VDDD.n3162 VDDD.n628 4.51401
R4769 VDDD.n3167 VDDD.n3166 4.51401
R4770 VDDD.n3114 VDDD.n663 4.51401
R4771 VDDD.n3119 VDDD.n655 4.51401
R4772 VDDD.n3078 VDDD.n3077 4.51401
R4773 VDDD.n746 VDDD.n745 4.51401
R4774 VDDD.n3274 VDDD.n566 4.51401
R4775 VDDD.n3265 VDDD.n3264 4.51401
R4776 VDDD.n867 VDDD.n865 4.51401
R4777 VDDD.n1047 VDDD.n1046 4.51401
R4778 VDDD.n3025 VDDD.n3024 4.51401
R4779 VDDD.n1090 VDDD.n1089 4.51401
R4780 VDDD.n3072 VDDD.n751 4.51401
R4781 VDDD.n756 VDDD.n755 4.51401
R4782 VDDD.n900 VDDD.n898 4.51401
R4783 VDDD.n1004 VDDD.n1003 4.51401
R4784 VDDD.n3015 VDDD.n1097 4.51401
R4785 VDDD.n1110 VDDD.n1109 4.51401
R4786 VDDD.n1427 VDDD.n1426 4.51401
R4787 VDDD.n1421 VDDD.n1420 4.51401
R4788 VDDD.n1515 VDDD.n1323 4.51401
R4789 VDDD.n1328 VDDD.n1327 4.51401
R4790 VDDD.n1139 VDDD.n1137 4.51401
R4791 VDDD.n1234 VDDD.n1233 4.51401
R4792 VDDD.n2797 VDDD.n2795 4.51401
R4793 VDDD.n2851 VDDD.n2850 4.51401
R4794 VDDD.n2755 VDDD.n1283 4.51401
R4795 VDDD.n2760 VDDD.n2759 4.51401
R4796 VDDD.n1318 VDDD.n1316 4.51401
R4797 VDDD.n1559 VDDD.n1558 4.51401
R4798 VDDD.n2962 VDDD.n1239 4.51401
R4799 VDDD.n2954 VDDD.n2953 4.51401
R4800 VDDD.n2580 VDDD.n1635 4.51401
R4801 VDDD.n2572 VDDD.n2571 4.51401
R4802 VDDD.n2207 VDDD.n2031 4.51401
R4803 VDDD.n2212 VDDD.n2027 4.51401
R4804 VDDD.n1630 VDDD.n1584 4.51401
R4805 VDDD.n2585 VDDD.n1577 4.51401
R4806 VDDD.n1880 VDDD.n1680 4.51401
R4807 VDDD.n1871 VDDD.n1867 4.51401
R4808 VDDD.n1771 VDDD.n1770 4.51401
R4809 VDDD.n1765 VDDD.n1764 4.51401
R4810 VDDD.n2705 VDDD.n1566 4.51401
R4811 VDDD.n2688 VDDD.n1571 4.51401
R4812 VDDD.n2153 VDDD.n2047 4.51401
R4813 VDDD.n2158 VDDD.n2157 4.51401
R4814 VDDD.n2424 VDDD.n2422 4.51401
R4815 VDDD.n2483 VDDD.n2482 4.51401
R4816 VDDD.n2339 VDDD.n2338 4.51401
R4817 VDDD.n1957 VDDD.n1956 4.51401
R4818 VDDD.n2375 VDDD.n2373 4.51401
R4819 VDDD.n2380 VDDD.n2379 4.51401
R4820 VDDD.n2092 VDDD.n2073 4.51401
R4821 VDDD.n2102 VDDD.n2068 4.51401
R4822 VDDD.n2333 VDDD.n1961 4.51401
R4823 VDDD.n1966 VDDD.n1965 4.51401
R4824 VDDD.n161 VDDD.n160 4.51401
R4825 VDDD.n203 VDDD.n202 4.51401
R4826 VDDD.n3685 VDDD.n3684 4.5005
R4827 VDDD.n3683 VDDD.n3682 4.5005
R4828 VDDD.n3679 VDDD.n3678 4.5005
R4829 VDDD.n3517 VDDD.n3516 4.5005
R4830 VDDD.n3501 VDDD.n3499 4.5005
R4831 VDDD.n3525 VDDD.n3524 4.5005
R4832 VDDD.n3571 VDDD.n3570 4.5005
R4833 VDDD.n3479 VDDD.n3478 4.5005
R4834 VDDD.n3476 VDDD.n359 4.5005
R4835 VDDD.n3621 VDDD.n3620 4.5005
R4836 VDDD.n3618 VDDD.n3617 4.5005
R4837 VDDD.n3628 VDDD.n3627 4.5005
R4838 VDDD.n438 VDDD.n437 4.5005
R4839 VDDD.n441 VDDD.n440 4.5005
R4840 VDDD.n383 VDDD.n382 4.5005
R4841 VDDD.n484 VDDD.n483 4.5005
R4842 VDDD.n492 VDDD.n491 4.5005
R4843 VDDD.n494 VDDD.n487 4.5005
R4844 VDDD.n3468 VDDD.n3467 4.5005
R4845 VDDD.n3455 VDDD.n3454 4.5005
R4846 VDDD.n3458 VDDD.n3294 4.5005
R4847 VDDD.n3317 VDDD.n3316 4.5005
R4848 VDDD.n3416 VDDD.n3415 4.5005
R4849 VDDD.n3321 VDDD.n3315 4.5005
R4850 VDDD.n698 VDDD.n691 4.5005
R4851 VDDD.n702 VDDD.n701 4.5005
R4852 VDDD.n703 VDDD.n694 4.5005
R4853 VDDD.n3113 VDDD.n3112 4.5005
R4854 VDDD.n661 VDDD.n659 4.5005
R4855 VDDD.n3121 VDDD.n3120 4.5005
R4856 VDDD.n3161 VDDD.n3160 4.5005
R4857 VDDD.n632 VDDD.n631 4.5005
R4858 VDDD.n624 VDDD.n623 4.5005
R4859 VDDD.n3273 VDDD.n3272 4.5005
R4860 VDDD.n3260 VDDD.n569 4.5005
R4861 VDDD.n3263 VDDD.n572 4.5005
R4862 VDDD.n3071 VDDD.n3070 4.5005
R4863 VDDD.n3069 VDDD.n3068 4.5005
R4864 VDDD.n3065 VDDD.n3064 4.5005
R4865 VDDD.n822 VDDD.n821 4.5005
R4866 VDDD.n834 VDDD.n833 4.5005
R4867 VDDD.n835 VDDD.n825 4.5005
R4868 VDDD.n866 VDDD.n862 4.5005
R4869 VDDD.n1052 VDDD.n1051 4.5005
R4870 VDDD.n870 VDDD.n864 4.5005
R4871 VDDD.n899 VDDD.n894 4.5005
R4872 VDDD.n1009 VDDD.n1008 4.5005
R4873 VDDD.n897 VDDD.n895 4.5005
R4874 VDDD.n1514 VDDD.n1513 4.5005
R4875 VDDD.n1512 VDDD.n1511 4.5005
R4876 VDDD.n1508 VDDD.n1507 4.5005
R4877 VDDD.n1354 VDDD.n1347 4.5005
R4878 VDDD.n1359 VDDD.n1358 4.5005
R4879 VDDD.n1360 VDDD.n1350 4.5005
R4880 VDDD.n3014 VDDD.n3013 4.5005
R4881 VDDD.n1106 VDDD.n1105 4.5005
R4882 VDDD.n1108 VDDD.n1107 4.5005
R4883 VDDD.n2970 VDDD.n2969 4.5005
R4884 VDDD.n1145 VDDD.n1140 4.5005
R4885 VDDD.n1146 VDDD.n1144 4.5005
R4886 VDDD.n2717 VDDD.n2716 4.5005
R4887 VDDD.n1319 VDDD.n1317 4.5005
R4888 VDDD.n1522 VDDD.n1519 4.5005
R4889 VDDD.n2754 VDDD.n2753 4.5005
R4890 VDDD.n1288 VDDD.n1287 4.5005
R4891 VDDD.n1279 VDDD.n1278 4.5005
R4892 VDDD.n2796 VDDD.n1254 4.5005
R4893 VDDD.n2856 VDDD.n2855 4.5005
R4894 VDDD.n1257 VDDD.n1256 4.5005
R4895 VDDD.n2961 VDDD.n2960 4.5005
R4896 VDDD.n2949 VDDD.n1242 4.5005
R4897 VDDD.n2952 VDDD.n1245 4.5005
R4898 VDDD.n1720 VDDD.n1712 4.5005
R4899 VDDD.n1722 VDDD.n1721 4.5005
R4900 VDDD.n1723 VDDD.n1715 4.5005
R4901 VDDD.n1879 VDDD.n1878 4.5005
R4902 VDDD.n1868 VDDD.n1682 4.5005
R4903 VDDD.n1873 VDDD.n1872 4.5005
R4904 VDDD.n1629 VDDD.n1628 4.5005
R4905 VDDD.n1585 VDDD.n1579 4.5005
R4906 VDDD.n2587 VDDD.n2586 4.5005
R4907 VDDD.n2704 VDDD.n2703 4.5005
R4908 VDDD.n2685 VDDD.n2684 4.5005
R4909 VDDD.n2690 VDDD.n2689 4.5005
R4910 VDDD.n1918 VDDD.n1908 4.5005
R4911 VDDD.n1922 VDDD.n1921 4.5005
R4912 VDDD.n1923 VDDD.n1911 4.5005
R4913 VDDD.n2423 VDDD.n1650 4.5005
R4914 VDDD.n2488 VDDD.n2487 4.5005
R4915 VDDD.n1653 VDDD.n1652 4.5005
R4916 VDDD.n2579 VDDD.n2578 4.5005
R4917 VDDD.n2567 VDDD.n1638 4.5005
R4918 VDDD.n2570 VDDD.n1642 4.5005
R4919 VDDD.n2374 VDDD.n1674 4.5005
R4920 VDDD.n2385 VDDD.n2384 4.5005
R4921 VDDD.n2378 VDDD.n1676 4.5005
R4922 VDDD.n2095 VDDD.n2094 4.5005
R4923 VDDD.n2096 VDDD.n2070 4.5005
R4924 VDDD.n2104 VDDD.n2103 4.5005
R4925 VDDD.n2152 VDDD.n2151 4.5005
R4926 VDDD.n2054 VDDD.n2053 4.5005
R4927 VDDD.n2051 VDDD.n2044 4.5005
R4928 VDDD.n2206 VDDD.n2205 4.5005
R4929 VDDD.n2203 VDDD.n2202 4.5005
R4930 VDDD.n2214 VDDD.n2213 4.5005
R4931 VDDD.n2332 VDDD.n2331 4.5005
R4932 VDDD.n2330 VDDD.n2329 4.5005
R4933 VDDD.n2326 VDDD.n2325 4.5005
R4934 VDDD.n162 VDDD.n121 4.5005
R4935 VDDD.n167 VDDD.n166 4.5005
R4936 VDDD.n168 VDDD.n117 4.5005
R4937 VDDD.n54 VDDD.n53 4.5005
R4938 VDDD.n65 VDDD.n64 4.5005
R4939 VDDD.n58 VDDD.n57 4.5005
R4940 VDDD.n3719 VDDD.n3718 4.5005
R4941 VDDD.n3712 VDDD.n3711 4.5005
R4942 VDDD.n3713 VDDD.n39 4.5005
R4943 VDDD.n3761 VDDD.n21 4.5005
R4944 VDDD.n3771 VDDD.n3770 4.5005
R4945 VDDD.n24 VDDD.n22 4.5005
R4946 VDDD.n798 VDDD.n797 4.47034
R4947 VDDD.n3251 VDDD.n574 4.41955
R4948 VDDD.n950 VDDD.n949 4.41955
R4949 VDDD.n534 VDDD.n518 4.38907
R4950 VDDD.n3831 VDDD.n3830 4.36875
R4951 VDDD.n249 VDDD.n248 4.36875
R4952 VDDD.n248 VDDD.n247 4.36875
R4953 VDDD.n3439 VDDD.n3304 4.36875
R4954 VDDD.n3408 VDDD.n3325 4.36875
R4955 VDDD.n3408 VDDD.n3407 4.36875
R4956 VDDD.n3402 VDDD.n3326 4.36875
R4957 VDDD.n3402 VDDD.n3401 4.36875
R4958 VDDD.n416 VDDD.n413 4.36875
R4959 VDDD.n416 VDDD.n415 4.36875
R4960 VDDD.n582 VDDD.n581 4.36875
R4961 VDDD.n3258 VDDD.n571 4.36875
R4962 VDDD.n3251 VDDD.n3250 4.36875
R4963 VDDD.n799 VDDD.n798 4.36875
R4964 VDDD.n796 VDDD.n788 4.36875
R4965 VDDD.n1040 VDDD.n873 4.36875
R4966 VDDD.n1034 VDDD.n1033 4.36875
R4967 VDDD.n985 VDDD.n984 4.36875
R4968 VDDD.n949 VDDD.n948 4.36875
R4969 VDDD.n1386 VDDD.n1100 4.36875
R4970 VDDD.n1487 VDDD.n1340 4.36875
R4971 VDDD.n2980 VDDD.n2979 4.36875
R4972 VDDD.n2787 VDDD.n2786 4.36875
R4973 VDDD.n2793 VDDD.n1253 4.36875
R4974 VDDD.n2896 VDDD.n2895 4.36875
R4975 VDDD.n1603 VDDD.n1602 4.36875
R4976 VDDD.n2638 VDDD.n2626 4.36875
R4977 VDDD.n2420 VDDD.n1649 4.36875
R4978 VDDD.n3732 VDDD.n36 4.36875
R4979 VDDD.n3702 VDDD.n3701 4.36875
R4980 VDDD.n143 VDDD.n126 4.36875
R4981 VDDD.n134 VDDD.n131 4.36875
R4982 VDDD.n524 VDDD.n367 4.35149
R4983 VDDD.n3236 VDDD.n3235 4.33769
R4984 VDDD.n2296 VDDD.n2295 4.29549
R4985 VDDD.n506 VDDD.n505 4.26717
R4986 VDDD.n2079 VDDD.n2077 4.26717
R4987 VDDD.n511 VDDD.n509 4.16908
R4988 VDDD.n3146 VDDD.n3145 4.14168
R4989 VDDD.n1431 VDDD.n1344 4.14168
R4990 VDDD.n681 VDDD.n680 4.06399
R4991 VDDD.n2817 VDDD.n1243 4.06399
R4992 VDDD.n2881 VDDD.n2880 4.06399
R4993 VDDD.n1703 VDDD.n1702 4.06399
R4994 VDDD.n305 VDDD.n285 4.02033
R4995 VDDD.n266 VDDD.n261 4.02033
R4996 VDDD.n266 VDDD.n265 4.02033
R4997 VDDD.n300 VDDD.n295 4.02033
R4998 VDDD.n300 VDDD.n298 4.02033
R4999 VDDD.n3288 VDDD.n482 4.02033
R5000 VDDD.n404 VDDD.n400 4.02033
R5001 VDDD.n404 VDDD.n403 4.02033
R5002 VDDD.n3360 VDDD.n3355 4.02033
R5003 VDDD.n3360 VDDD.n3358 4.02033
R5004 VDDD.n676 VDDD.n672 4.02033
R5005 VDDD.n676 VDDD.n675 4.02033
R5006 VDDD.n3195 VDDD.n3190 4.02033
R5007 VDDD.n3195 VDDD.n3193 4.02033
R5008 VDDD.n780 VDDD.n776 4.02033
R5009 VDDD.n780 VDDD.n779 4.02033
R5010 VDDD.n944 VDDD.n940 4.02033
R5011 VDDD.n944 VDDD.n943 4.02033
R5012 VDDD.n1445 VDDD.n1441 4.02033
R5013 VDDD.n1445 VDDD.n1444 4.02033
R5014 VDDD.n1178 VDDD.n1173 4.02033
R5015 VDDD.n1178 VDDD.n1176 4.02033
R5016 VDDD.n1303 VDDD.n1299 4.02033
R5017 VDDD.n1303 VDDD.n1302 4.02033
R5018 VDDD.n2893 VDDD.n2888 4.02033
R5019 VDDD.n2893 VDDD.n2891 4.02033
R5020 VDDD.n1832 VDDD.n1829 4.02033
R5021 VDDD.n1697 VDDD.n1693 4.02033
R5022 VDDD.n1697 VDDD.n1696 4.02033
R5023 VDDD.n2634 VDDD.n2629 4.02033
R5024 VDDD.n2634 VDDD.n2632 4.02033
R5025 VDDD.n1896 VDDD.n1892 4.02033
R5026 VDDD.n1896 VDDD.n1895 4.02033
R5027 VDDD.n2515 VDDD.n2510 4.02033
R5028 VDDD.n2515 VDDD.n2513 4.02033
R5029 VDDD.n1993 VDDD.n1989 4.02033
R5030 VDDD.n1993 VDDD.n1992 4.02033
R5031 VDDD.n2163 VDDD.n2162 4.02033
R5032 VDDD.n1986 VDDD.n1985 4.02033
R5033 VDDD.n2250 VDDD.n2245 4.02033
R5034 VDDD.n2250 VDDD.n2248 4.02033
R5035 VDDD.n3448 VDDD.n3296 4.00858
R5036 VDDD.n525 VDDD.n524 3.99734
R5037 VDDD.n506 VDDD.n504 3.8405
R5038 VDDD.n2079 VDDD.n2078 3.8405
R5039 VDDD.n1709 VDDD.n1707 3.80876
R5040 VDDD.n323 VDDD.n322 3.76521
R5041 VDDD.n3538 VDDD.n3491 3.76521
R5042 VDDD.n3379 VDDD.n3377 3.76521
R5043 VDDD.n3383 VDDD.n3336 3.76521
R5044 VDDD.n709 VDDD.n707 3.76521
R5045 VDDD.n829 VDDD.n828 3.76521
R5046 VDDD.n1067 VDDD.n851 3.76521
R5047 VDDD.n1021 VDDD.n1020 3.76521
R5048 VDDD.n1015 VDDD.n889 3.76521
R5049 VDDD.n923 VDDD.n920 3.76521
R5050 VDDD.n973 VDDD.n923 3.76521
R5051 VDDD.n967 VDDD.n926 3.76521
R5052 VDDD.n1460 VDDD.n1458 3.76521
R5053 VDDD.n2989 VDDD.n2988 3.76521
R5054 VDDD.n2834 VDDD.n2808 3.76521
R5055 VDDD.n2840 VDDD.n2804 3.76521
R5056 VDDD.n2804 VDDD.n2801 3.76521
R5057 VDDD.n2771 VDDD.n2770 3.76521
R5058 VDDD.n2769 VDDD.n2768 3.76521
R5059 VDDD.n2719 VDDD.n1315 3.76521
R5060 VDDD.n1526 VDDD.n1524 3.76521
R5061 VDDD.n2927 VDDD.n2869 3.76521
R5062 VDDD.n1619 VDDD.n1591 3.76521
R5063 VDDD.n1624 VDDD.n1588 3.76521
R5064 VDDD.n2665 VDDD.n2612 3.76521
R5065 VDDD.n1926 VDDD.n1925 3.76521
R5066 VDDD.n1917 VDDD.n1916 3.76521
R5067 VDDD.n2399 VDDD.n2398 3.76521
R5068 VDDD.n2393 VDDD.n2392 3.76521
R5069 VDDD.n3755 VDDD.n3754 3.76521
R5070 VDDD.n3243 VDDD.n3242 3.75222
R5071 VDDD.n509 VDDD.n503 3.7277
R5072 VDDD.n1451 VDDD.n1450 3.70844
R5073 VDDD.n2419 VDDD.n2418 3.70844
R5074 VDDD.n3606 VDDD.n345 3.70298
R5075 VDDD.n3637 VDDD.n3636 3.70298
R5076 VDDD.n3512 VDDD.n3511 3.70298
R5077 VDDD.n3202 VDDD.n3186 3.70298
R5078 VDDD.n1230 VDDD.n1229 3.70298
R5079 VDDD.n1781 VDDD.n1780 3.70298
R5080 VDDD.n2135 VDDD.n2058 3.70298
R5081 VDDD.n2191 VDDD.n2032 3.70298
R5082 VDDD.n2943 VDDD.n1248 3.69947
R5083 VDDD.n1833 VDDD.n1568 3.59719
R5084 VDDD.n301 VDDD.n289 3.56582
R5085 VDDD.n3361 VDDD.n3349 3.56582
R5086 VDDD.n621 VDDD.n620 3.56582
R5087 VDDD.n804 VDDD.n803 3.56582
R5088 VDDD.n267 VDDD.n258 3.52514
R5089 VDDD.n3830 VDDD.n3829 3.50526
R5090 VDDD.n3702 VDDD.n51 3.50526
R5091 VDDD.n143 VDDD.n142 3.50526
R5092 VDDD.n134 VDDD.n133 3.50526
R5093 VDDD.n396 VDDD.n394 3.47876
R5094 VDDD.n2562 VDDD.n2561 3.47425
R5095 VDDD.n2147 VDDD.n2146 3.47425
R5096 VDDD.n2223 VDDD.n2026 3.47425
R5097 VDDD.n2224 VDDD.n2223 3.47425
R5098 VDDD.n2300 VDDD.n2299 3.47425
R5099 VDDD.n112 VDDD.n111 3.43925
R5100 VDDD.n3696 VDDD.n3695 3.43925
R5101 VDDD.n3724 VDDD.n3723 3.43925
R5102 VDDD.n3721 VDDD.n3720 3.43925
R5103 VDDD.n3767 VDDD.n3766 3.43925
R5104 VDDD.n3763 VDDD.n3762 3.43925
R5105 VDDD.n3576 VDDD.n3575 3.43925
R5106 VDDD.n3573 VDDD.n3572 3.43925
R5107 VDDD.n3523 VDDD.n3522 3.43925
R5108 VDDD.n3519 VDDD.n3518 3.43925
R5109 VDDD.n213 VDDD.n206 3.43925
R5110 VDDD.n3687 VDDD.n3686 3.43925
R5111 VDDD.n3626 VDDD.n3625 3.43925
R5112 VDDD.n3623 VDDD.n3622 3.43925
R5113 VDDD.n3459 VDDD.n361 3.43925
R5114 VDDD.n3470 VDDD.n3469 3.43925
R5115 VDDD.n560 VDDD.n559 3.43925
R5116 VDDD.n3284 VDDD.n3283 3.43925
R5117 VDDD.n445 VDDD.n444 3.43925
R5118 VDDD.n436 VDDD.n435 3.43925
R5119 VDDD.n3412 VDDD.n3411 3.43925
R5120 VDDD.n3319 VDDD.n3318 3.43925
R5121 VDDD.n3166 VDDD.n3165 3.43925
R5122 VDDD.n3163 VDDD.n3162 3.43925
R5123 VDDD.n3119 VDDD.n3118 3.43925
R5124 VDDD.n3115 VDDD.n3114 3.43925
R5125 VDDD.n747 VDDD.n746 3.43925
R5126 VDDD.n3077 VDDD.n3076 3.43925
R5127 VDDD.n3264 VDDD.n563 3.43925
R5128 VDDD.n3275 VDDD.n3274 3.43925
R5129 VDDD.n1048 VDDD.n1047 3.43925
R5130 VDDD.n868 VDDD.n867 3.43925
R5131 VDDD.n1091 VDDD.n1090 3.43925
R5132 VDDD.n3024 VDDD.n3023 3.43925
R5133 VDDD.n755 VDDD.n748 3.43925
R5134 VDDD.n3073 VDDD.n3072 3.43925
R5135 VDDD.n1005 VDDD.n1004 3.43925
R5136 VDDD.n901 VDDD.n900 3.43925
R5137 VDDD.n1109 VDDD.n1094 3.43925
R5138 VDDD.n3016 VDDD.n3015 3.43925
R5139 VDDD.n1422 VDDD.n1421 3.43925
R5140 VDDD.n1426 VDDD.n1425 3.43925
R5141 VDDD.n1327 VDDD.n1321 3.43925
R5142 VDDD.n1516 VDDD.n1515 3.43925
R5143 VDDD.n1235 VDDD.n1234 3.43925
R5144 VDDD.n2966 VDDD.n1139 3.43925
R5145 VDDD.n2852 VDDD.n2851 3.43925
R5146 VDDD.n2798 VDDD.n2797 3.43925
R5147 VDDD.n2759 VDDD.n2758 3.43925
R5148 VDDD.n2756 VDDD.n2755 3.43925
R5149 VDDD.n1560 VDDD.n1559 3.43925
R5150 VDDD.n2713 VDDD.n1318 3.43925
R5151 VDDD.n2953 VDDD.n1236 3.43925
R5152 VDDD.n2963 VDDD.n2962 3.43925
R5153 VDDD.n2571 VDDD.n1632 3.43925
R5154 VDDD.n2581 VDDD.n2580 3.43925
R5155 VDDD.n2212 VDDD.n2211 3.43925
R5156 VDDD.n2208 VDDD.n2207 3.43925
R5157 VDDD.n1871 VDDD.n1678 3.43925
R5158 VDDD.n1881 VDDD.n1880 3.43925
R5159 VDDD.n1766 VDDD.n1765 3.43925
R5160 VDDD.n1770 VDDD.n1769 3.43925
R5161 VDDD.n2688 VDDD.n1563 3.43925
R5162 VDDD.n2706 VDDD.n2705 3.43925
R5163 VDDD.n2157 VDDD.n2156 3.43925
R5164 VDDD.n2154 VDDD.n2153 3.43925
R5165 VDDD.n1958 VDDD.n1957 3.43925
R5166 VDDD.n2338 VDDD.n2337 3.43925
R5167 VDDD.n2381 VDDD.n2380 3.43925
R5168 VDDD.n2376 VDDD.n2375 3.43925
R5169 VDDD.n1965 VDDD.n1959 3.43925
R5170 VDDD.n2334 VDDD.n2333 3.43925
R5171 VDDD.n62 VDDD.n55 3.4105
R5172 VDDD.n63 VDDD.n56 3.4105
R5173 VDDD.n44 VDDD.n42 3.4105
R5174 VDDD.n3710 VDDD.n40 3.4105
R5175 VDDD.n25 VDDD.n23 3.4105
R5176 VDDD.n3769 VDDD.n3768 3.4105
R5177 VDDD.n3474 VDDD.n3472 3.4105
R5178 VDDD.n3477 VDDD.n360 3.4105
R5179 VDDD.n3520 VDDD.n3502 3.4105
R5180 VDDD.n3521 VDDD.n3500 3.4105
R5181 VDDD.n210 VDDD.n208 3.4105
R5182 VDDD.n3681 VDDD.n3680 3.4105
R5183 VDDD.n344 VDDD.n342 3.4105
R5184 VDDD.n340 VDDD.n339 3.4105
R5185 VDDD.n365 VDDD.n363 3.4105
R5186 VDDD.n3457 VDDD.n3456 3.4105
R5187 VDDD.n489 VDDD.n485 3.4105
R5188 VDDD.n490 VDDD.n486 3.4105
R5189 VDDD.n385 VDDD.n384 3.4105
R5190 VDDD.n443 VDDD.n442 3.4105
R5191 VDDD.n3320 VDDD.n3314 3.4105
R5192 VDDD.n3414 VDDD.n3413 3.4105
R5193 VDDD.n629 VDDD.n627 3.4105
R5194 VDDD.n630 VDDD.n625 3.4105
R5195 VDDD.n3116 VDDD.n662 3.4105
R5196 VDDD.n3117 VDDD.n660 3.4105
R5197 VDDD.n699 VDDD.n692 3.4105
R5198 VDDD.n700 VDDD.n693 3.4105
R5199 VDDD.n567 VDDD.n565 3.4105
R5200 VDDD.n3262 VDDD.n3261 3.4105
R5201 VDDD.n869 VDDD.n863 3.4105
R5202 VDDD.n1050 VDDD.n1049 3.4105
R5203 VDDD.n831 VDDD.n823 3.4105
R5204 VDDD.n832 VDDD.n824 3.4105
R5205 VDDD.n752 VDDD.n750 3.4105
R5206 VDDD.n3067 VDDD.n3066 3.4105
R5207 VDDD.n902 VDDD.n896 3.4105
R5208 VDDD.n1007 VDDD.n1006 3.4105
R5209 VDDD.n1098 VDDD.n1096 3.4105
R5210 VDDD.n1104 VDDD.n1103 3.4105
R5211 VDDD.n1424 VDDD.n1348 3.4105
R5212 VDDD.n1423 VDDD.n1349 3.4105
R5213 VDDD.n1324 VDDD.n1322 3.4105
R5214 VDDD.n1510 VDDD.n1509 3.4105
R5215 VDDD.n2968 VDDD.n2967 3.4105
R5216 VDDD.n1143 VDDD.n1141 3.4105
R5217 VDDD.n2799 VDDD.n1255 3.4105
R5218 VDDD.n2854 VDDD.n2853 3.4105
R5219 VDDD.n1284 VDDD.n1282 3.4105
R5220 VDDD.n1286 VDDD.n1280 3.4105
R5221 VDDD.n2715 VDDD.n2714 3.4105
R5222 VDDD.n1518 VDDD.n1320 3.4105
R5223 VDDD.n1240 VDDD.n1238 3.4105
R5224 VDDD.n2951 VDDD.n2950 3.4105
R5225 VDDD.n1636 VDDD.n1634 3.4105
R5226 VDDD.n2569 VDDD.n2568 3.4105
R5227 VDDD.n2209 VDDD.n2030 3.4105
R5228 VDDD.n2210 VDDD.n2029 3.4105
R5229 VDDD.n2584 VDDD.n2583 3.4105
R5230 VDDD.n2583 VDDD.n1631 3.4105
R5231 VDDD.n2585 VDDD.n2584 3.4105
R5232 VDDD.n1631 VDDD.n1630 3.4105
R5233 VDDD.n1586 VDDD.n1583 3.4105
R5234 VDDD.n1581 VDDD.n1580 3.4105
R5235 VDDD.n1681 VDDD.n1679 3.4105
R5236 VDDD.n1870 VDDD.n1869 3.4105
R5237 VDDD.n1768 VDDD.n1713 3.4105
R5238 VDDD.n1767 VDDD.n1714 3.4105
R5239 VDDD.n1567 VDDD.n1565 3.4105
R5240 VDDD.n2687 VDDD.n2686 3.4105
R5241 VDDD.n2048 VDDD.n2046 3.4105
R5242 VDDD.n2052 VDDD.n2045 3.4105
R5243 VDDD.n2484 VDDD.n1564 3.4105
R5244 VDDD.n2425 VDDD.n1564 3.4105
R5245 VDDD.n2484 VDDD.n2483 3.4105
R5246 VDDD.n2425 VDDD.n2424 3.4105
R5247 VDDD.n2426 VDDD.n1651 3.4105
R5248 VDDD.n2486 VDDD.n2485 3.4105
R5249 VDDD.n1919 VDDD.n1909 3.4105
R5250 VDDD.n1920 VDDD.n1910 3.4105
R5251 VDDD.n1677 VDDD.n1675 3.4105
R5252 VDDD.n2383 VDDD.n2382 3.4105
R5253 VDDD.n2101 VDDD.n1883 3.4105
R5254 VDDD.n2072 VDDD.n1883 3.4105
R5255 VDDD.n2102 VDDD.n2101 3.4105
R5256 VDDD.n2073 VDDD.n2072 3.4105
R5257 VDDD.n2098 VDDD.n2097 3.4105
R5258 VDDD.n2100 VDDD.n2071 3.4105
R5259 VDDD.n1962 VDDD.n1960 3.4105
R5260 VDDD.n2328 VDDD.n2327 3.4105
R5261 VDDD.n205 VDDD.n204 3.4105
R5262 VDDD.n205 VDDD.n115 3.4105
R5263 VDDD.n204 VDDD.n203 3.4105
R5264 VDDD.n161 VDDD.n115 3.4105
R5265 VDDD.n164 VDDD.n163 3.4105
R5266 VDDD.n165 VDDD.n116 3.4105
R5267 VDDD.n3132 VDDD.n651 3.38874
R5268 VDDD.n598 VDDD.n597 3.38874
R5269 VDDD.n889 VDDD.n886 3.38874
R5270 VDDD.n1621 VDDD.n1588 3.38874
R5271 VDDD.n2392 VDDD.n1668 3.38874
R5272 VDDD.t1437 VDDD.t677 3.35739
R5273 VDDD.t1961 VDDD.t185 3.35739
R5274 VDDD.t438 VDDD 3.35739
R5275 VDDD.t1124 VDDD.t774 3.35739
R5276 VDDD.t884 VDDD.t220 3.35739
R5277 VDDD.t259 VDDD.t1896 3.35739
R5278 VDDD.t943 VDDD.t1066 3.35739
R5279 VDDD VDDD.t1502 3.35739
R5280 VDDD.t520 VDDD.t577 3.35739
R5281 VDDD.t1466 VDDD.t401 3.35739
R5282 VDDD.t1670 VDDD.t1432 3.35739
R5283 VDDD.t1088 VDDD.t39 3.35739
R5284 VDDD VDDD.t553 3.35739
R5285 VDDD.t1280 VDDD.t1830 3.35739
R5286 VDDD.n507 VDDD.n506 3.29837
R5287 VDDD.n2080 VDDD.n2079 3.29837
R5288 VDDD.n792 VDDD.n791 3.26444
R5289 VDDD.n579 VDDD.n577 3.25799
R5290 VDDD.n787 VDDD.n784 3.25799
R5291 VDDD.n2563 VDDD.n2562 3.2477
R5292 VDDD.n2561 VDDD.n1644 3.2477
R5293 VDDD.n2148 VDDD.n2147 3.2477
R5294 VDDD.n2219 VDDD.n2217 3.2477
R5295 VDDD.n2225 VDDD.n2224 3.2477
R5296 VDDD.n2302 VDDD.n1977 3.2477
R5297 VDDD.n2299 VDDD.n1978 3.2477
R5298 VDDD.n3221 VDDD.n3220 3.21089
R5299 VDDD.n250 VDDD.n237 3.2005
R5300 VDDD.n257 VDDD.n233 3.2005
R5301 VDDD.n1600 VDDD.n1598 3.2005
R5302 VDDD.n3670 VDDD.n3669 3.17405
R5303 VDDD.n431 VDDD.n430 3.17405
R5304 VDDD.n3214 VDDD.n3213 3.17405
R5305 VDDD.n3057 VDDD.n3056 3.17405
R5306 VDDD.n1151 VDDD.n1150 3.17405
R5307 VDDD.n1824 VDDD.n1822 3.17405
R5308 VDDD.n1719 VDDD.n1710 3.17405
R5309 VDDD.n2121 VDDD.n2120 3.17405
R5310 VDDD.n2181 VDDD.n2036 3.17405
R5311 VDDD.n2003 VDDD.n2002 3.17405
R5312 VDDD.n541 VDDD.n540 3.13726
R5313 VDDD.n395 VDDD.n394 3.13093
R5314 VDDD.n3152 VDDD.n635 3.12116
R5315 VDDD.n2787 VDDD.n1263 3.12116
R5316 VDDD.n241 VDDD.n240 3.06827
R5317 VDDD.n422 VDDD.n421 3.06827
R5318 VDDD.n2015 VDDD.n2014 3.06827
R5319 VDDD.n266 VDDD.n262 3.05586
R5320 VDDD.n405 VDDD.n404 3.05586
R5321 VDDD.n677 VDDD.n676 3.05586
R5322 VDDD.n782 VDDD.n780 3.05586
R5323 VDDD.n1446 VDDD.n1445 3.05586
R5324 VDDD.n1304 VDDD.n1303 3.05586
R5325 VDDD.n1698 VDDD.n1697 3.05586
R5326 VDDD.n1897 VDDD.n1896 3.05586
R5327 VDDD.n1994 VDDD.n1993 3.05586
R5328 VDDD.n2699 VDDD.n1569 3.05371
R5329 VDDD.n300 VDDD.n299 3.04861
R5330 VDDD.n305 VDDD.n304 3.04861
R5331 VDDD.n3360 VDDD.n3359 3.04861
R5332 VDDD.n3195 VDDD.n3194 3.04861
R5333 VDDD.n945 VDDD.n944 3.04861
R5334 VDDD.n1178 VDDD.n1177 3.04861
R5335 VDDD.n2893 VDDD.n2892 3.04861
R5336 VDDD.n2634 VDDD.n2633 3.04861
R5337 VDDD.n2515 VDDD.n2514 3.04861
R5338 VDDD.n2250 VDDD.n2249 3.04861
R5339 VDDD.n2018 VDDD.n1986 3.04861
R5340 VDDD.n3288 VDDD.n3287 3.04861
R5341 VDDD.n546 VDDD.n503 3.04861
R5342 VDDD.n3240 VDDD.n3239 3.04861
R5343 VDDD.n1213 VDDD.n1159 3.01588
R5344 VDDD.n1193 VDDD.n1166 3.01588
R5345 VDDD.n2550 VDDD.n2496 3.01588
R5346 VDDD.n2530 VDDD.n2503 3.01588
R5347 VDDD.n2285 VDDD.n2231 3.01588
R5348 VDDD.n2265 VDDD.n2238 3.01588
R5349 VDDD.n555 VDDD.n498 2.99733
R5350 VDDD.n3441 VDDD.n3303 2.99733
R5351 VDDD.n637 VDDD.n636 2.99733
R5352 VDDD.n1490 VDDD.n1338 2.99733
R5353 VDDD.n2417 VDDD.n1655 2.99733
R5354 VDDD.n542 VDDD.n541 2.98548
R5355 VDDD.n2090 VDDD.n2085 2.96248
R5356 VDDD.n3001 VDDD.n3000 2.94653
R5357 VDDD.n301 VDDD.n292 2.91308
R5358 VDDD.n3361 VDDD.n3352 2.91308
R5359 VDDD.n620 VDDD.n577 2.91308
R5360 VDDD.n803 VDDD.n784 2.91308
R5361 VDDD.n1935 VDDD.n1934 2.91308
R5362 VDDD.n1936 VDDD.n1935 2.91308
R5363 VDDD.n1388 VDDD.n1387 2.89574
R5364 VDDD.n287 VDDD.n282 2.87861
R5365 VDDD.n496 VDDD.n479 2.87861
R5366 VDDD.n3301 VDDD.n3299 2.87861
R5367 VDDD.n3364 VDDD.n3344 2.87861
R5368 VDDD.n642 VDDD.n639 2.87861
R5369 VDDD.n809 VDDD.n807 2.87861
R5370 VDDD.n1493 VDDD.n1335 2.87861
R5371 VDDD.n2414 VDDD.n1657 2.87861
R5372 VDDD.n474 VDDD.n473 2.84494
R5373 VDDD.n3220 VDDD.n3218 2.78608
R5374 VDDD.n1210 VDDD.n1159 2.64665
R5375 VDDD.n1190 VDDD.n1166 2.64665
R5376 VDDD.n2547 VDDD.n2496 2.64665
R5377 VDDD.n2527 VDDD.n2503 2.64665
R5378 VDDD.n2282 VDDD.n2231 2.64665
R5379 VDDD.n2262 VDDD.n2238 2.64665
R5380 VDDD.n1938 VDDD.n1937 2.64481
R5381 VDDD.n3529 VDDD.n3528 2.63579
R5382 VDDD.n688 VDDD.n685 2.63579
R5383 VDDD.n590 VDDD.n586 2.63579
R5384 VDDD.n842 VDDD.n841 2.63579
R5385 VDDD.n846 VDDD.n843 2.63579
R5386 VDDD.n285 VDDD.n283 2.63539
R5387 VDDD.n261 VDDD.n259 2.63539
R5388 VDDD.n265 VDDD.n263 2.63539
R5389 VDDD.n295 VDDD.n293 2.63539
R5390 VDDD.n298 VDDD.n296 2.63539
R5391 VDDD.n482 VDDD.n480 2.63539
R5392 VDDD.n400 VDDD.n398 2.63539
R5393 VDDD.n403 VDDD.n401 2.63539
R5394 VDDD.n3355 VDDD.n3353 2.63539
R5395 VDDD.n3358 VDDD.n3356 2.63539
R5396 VDDD.n635 VDDD.n633 2.63539
R5397 VDDD.n672 VDDD.n670 2.63539
R5398 VDDD.n675 VDDD.n673 2.63539
R5399 VDDD.n3190 VDDD.n3188 2.63539
R5400 VDDD.n3193 VDDD.n3191 2.63539
R5401 VDDD.n776 VDDD.n774 2.63539
R5402 VDDD.n779 VDDD.n777 2.63539
R5403 VDDD.n940 VDDD.n938 2.63539
R5404 VDDD.n943 VDDD.n941 2.63539
R5405 VDDD.n1441 VDDD.n1439 2.63539
R5406 VDDD.n1444 VDDD.n1442 2.63539
R5407 VDDD.n1173 VDDD.n1171 2.63539
R5408 VDDD.n1176 VDDD.n1174 2.63539
R5409 VDDD.n1263 VDDD.n1261 2.63539
R5410 VDDD.n1299 VDDD.n1297 2.63539
R5411 VDDD.n1302 VDDD.n1300 2.63539
R5412 VDDD.n2888 VDDD.n2886 2.63539
R5413 VDDD.n2891 VDDD.n2889 2.63539
R5414 VDDD.n1829 VDDD.n1827 2.63539
R5415 VDDD.n1693 VDDD.n1691 2.63539
R5416 VDDD.n1696 VDDD.n1694 2.63539
R5417 VDDD.n2629 VDDD.n2627 2.63539
R5418 VDDD.n2632 VDDD.n2630 2.63539
R5419 VDDD.n1892 VDDD.n1890 2.63539
R5420 VDDD.n1895 VDDD.n1893 2.63539
R5421 VDDD.n2510 VDDD.n2508 2.63539
R5422 VDDD.n2513 VDDD.n2511 2.63539
R5423 VDDD.n1989 VDDD.n1987 2.63539
R5424 VDDD.n1992 VDDD.n1990 2.63539
R5425 VDDD.n2162 VDDD.n2160 2.63539
R5426 VDDD.n1985 VDDD.n1983 2.63539
R5427 VDDD.n2245 VDDD.n2243 2.63539
R5428 VDDD.n2248 VDDD.n2246 2.63539
R5429 VDDD.n288 VDDD.n286 2.61352
R5430 VDDD.n498 VDDD.n497 2.61352
R5431 VDDD.n3303 VDDD.n3302 2.61352
R5432 VDDD.n3348 VDDD.n3347 2.61352
R5433 VDDD.n638 VDDD.n637 2.61352
R5434 VDDD.n806 VDDD.n805 2.61352
R5435 VDDD.n1338 VDDD.n1337 2.61352
R5436 VDDD.n1656 VDDD.n1655 2.61352
R5437 VDDD.n515 VDDD.n513 2.53014
R5438 VDDD.n1543 VDDD.n1542 2.50603
R5439 VDDD.n1542 VDDD.n1541 2.50603
R5440 VDDD.n1541 VDDD.n1537 2.50603
R5441 VDDD.n2982 VDDD.n2981 2.48939
R5442 VDDD.n2978 VDDD.n1134 2.44862
R5443 VDDD.n3258 VDDD.n3257 2.4386
R5444 VDDD.n2958 VDDD.n2957 2.4386
R5445 VDDD.n3156 VDDD.n622 2.37764
R5446 VDDD.n284 VDDD.n283 2.37495
R5447 VDDD.n264 VDDD.n263 2.37495
R5448 VDDD.n260 VDDD.n259 2.37495
R5449 VDDD.n297 VDDD.n296 2.37495
R5450 VDDD.n294 VDDD.n293 2.37495
R5451 VDDD.n481 VDDD.n480 2.37495
R5452 VDDD.n402 VDDD.n401 2.37495
R5453 VDDD.n399 VDDD.n398 2.37495
R5454 VDDD.n3357 VDDD.n3356 2.37495
R5455 VDDD.n3354 VDDD.n3353 2.37495
R5456 VDDD.n634 VDDD.n633 2.37495
R5457 VDDD.n674 VDDD.n673 2.37495
R5458 VDDD.n671 VDDD.n670 2.37495
R5459 VDDD.n3192 VDDD.n3191 2.37495
R5460 VDDD.n3189 VDDD.n3188 2.37495
R5461 VDDD.n778 VDDD.n777 2.37495
R5462 VDDD.n775 VDDD.n774 2.37495
R5463 VDDD.n942 VDDD.n941 2.37495
R5464 VDDD.n939 VDDD.n938 2.37495
R5465 VDDD.n1443 VDDD.n1442 2.37495
R5466 VDDD.n1440 VDDD.n1439 2.37495
R5467 VDDD.n1175 VDDD.n1174 2.37495
R5468 VDDD.n1172 VDDD.n1171 2.37495
R5469 VDDD.n1262 VDDD.n1261 2.37495
R5470 VDDD.n1301 VDDD.n1300 2.37495
R5471 VDDD.n1298 VDDD.n1297 2.37495
R5472 VDDD.n2890 VDDD.n2889 2.37495
R5473 VDDD.n2887 VDDD.n2886 2.37495
R5474 VDDD.n1828 VDDD.n1827 2.37495
R5475 VDDD.n1695 VDDD.n1694 2.37495
R5476 VDDD.n1692 VDDD.n1691 2.37495
R5477 VDDD.n2631 VDDD.n2630 2.37495
R5478 VDDD.n2628 VDDD.n2627 2.37495
R5479 VDDD.n1894 VDDD.n1893 2.37495
R5480 VDDD.n1891 VDDD.n1890 2.37495
R5481 VDDD.n2512 VDDD.n2511 2.37495
R5482 VDDD.n2509 VDDD.n2508 2.37495
R5483 VDDD.n1991 VDDD.n1990 2.37495
R5484 VDDD.n1988 VDDD.n1987 2.37495
R5485 VDDD.n2161 VDDD.n2160 2.37495
R5486 VDDD.n1984 VDDD.n1983 2.37495
R5487 VDDD.n2247 VDDD.n2246 2.37495
R5488 VDDD.n2244 VDDD.n2243 2.37495
R5489 VDDD.n1543 VDDD.n1535 2.34263
R5490 VDDD.n1537 VDDD.n1536 2.34263
R5491 VDDD.n552 VDDD.n500 2.33701
R5492 VDDD.n412 VDDD.n411 2.33701
R5493 VDDD.n472 VDDD.n471 2.33701
R5494 VDDD.n3095 VDDD.n679 2.33701
R5495 VDDD.n951 VDDD.n937 2.33701
R5496 VDDD.n1474 VDDD.n1473 2.33701
R5497 VDDD.n1389 VDDD.n1388 2.33701
R5498 VDDD.n2982 VDDD.n1132 2.33701
R5499 VDDD.n2946 VDDD.n2945 2.33701
R5500 VDDD.n2945 VDDD.n2944 2.33701
R5501 VDDD.n2885 VDDD.n2882 2.33701
R5502 VDDD.n2896 VDDD.n2885 2.33701
R5503 VDDD.n1791 VDDD.n1790 2.33701
R5504 VDDD.n2076 VDDD.n1980 2.33701
R5505 VDDD.n3731 VDDD.n3730 2.33701
R5506 VDDD.n526 VDDD.n522 2.32777
R5507 VDDD.n3240 VDDD.n3173 2.28432
R5508 VDDD.n253 VDDD.n234 2.28407
R5509 VDDD.n254 VDDD.n253 2.28407
R5510 VDDD.n2695 VDDD.n1570 2.28407
R5511 VDDD.n2696 VDDD.n2695 2.28407
R5512 VDDD.n1833 VDDD.n1832 2.27488
R5513 VDDD.n3557 VDDD.n3556 2.25932
R5514 VDDD.n3528 VDDD.n3527 2.25932
R5515 VDDD.n3085 VDDD.n685 2.25932
R5516 VDDD.n3030 VDDD.n3029 2.25932
R5517 VDDD.n1087 VDDD.n1086 2.25932
R5518 VDDD.n1077 VDDD.n843 2.25932
R5519 VDDD.n997 VDDD.n996 2.25932
R5520 VDDD.n991 VDDD.n990 2.25932
R5521 VDDD.n1362 VDDD.n1353 2.25932
R5522 VDDD.n2738 VDDD.n1296 2.25932
R5523 VDDD.n2742 VDDD.n2741 2.25932
R5524 VDDD.n2906 VDDD.n2879 2.25932
R5525 VDDD.n1856 VDDD.n1855 2.25932
R5526 VDDD.n2598 VDDD.n1572 2.25932
R5527 VDDD.n2644 VDDD.n2622 2.25932
R5528 VDDD.n2359 VDDD.n2358 2.25932
R5529 VDDD.n2453 VDDD.n2452 2.25932
R5530 VDDD.n2479 VDDD.n2478 2.25932
R5531 VDDD.n2364 VDDD.n2363 2.25932
R5532 VDDD.n303 VDDD.n282 2.25312
R5533 VDDD.n3443 VDDD.n3299 2.25312
R5534 VDDD.n3364 VDDD.n3363 2.25312
R5535 VDDD.n3149 VDDD.n642 2.25312
R5536 VDDD.n620 VDDD.n619 2.25312
R5537 VDDD.n803 VDDD.n802 2.25312
R5538 VDDD.n1493 VDDD.n1492 2.25312
R5539 VDDD.n1942 VDDD.n1935 2.25312
R5540 VDDD.n302 VDDD.n301 2.25293
R5541 VDDD.n3362 VDDD.n3361 2.25293
R5542 VDDD.n916 VDDD.n915 2.23542
R5543 VDDD.n2957 VDDD.n2956 2.23542
R5544 VDDD.n956 VDDD.n955 2.23239
R5545 VDDD.n2558 VDDD.n2557 2.20671
R5546 VDDD.n2226 VDDD.n2023 2.20671
R5547 VDDD.n1371 VDDD.n1368 2.19479
R5548 VDDD.n1802 VDDD.n1684 2.19479
R5549 VDDD.n2981 VDDD.n2980 2.18463
R5550 VDDD.n289 VDDD.n288 2.13621
R5551 VDDD.n3349 VDDD.n3348 2.13621
R5552 VDDD.n622 VDDD.n621 2.13621
R5553 VDDD.n805 VDDD.n804 2.13621
R5554 VDDD.n3447 VDDD.n3296 2.13383
R5555 VDDD.n237 VDDD.n236 2.07374
R5556 VDDD.n255 VDDD.n233 2.07374
R5557 VDDD.n1598 VDDD.n1597 2.07374
R5558 VDDD.n2697 VDDD.n1569 2.07374
R5559 VDDD.n501 VDDD.n500 2.03225
R5560 VDDD.n411 VDDD.n410 2.03225
R5561 VDDD.n471 VDDD.n470 2.03225
R5562 VDDD.n679 VDDD.n669 2.03225
R5563 VDDD.n915 VDDD.n914 2.03225
R5564 VDDD.n937 VDDD.n935 2.03225
R5565 VDDD.n1390 VDDD.n1389 2.03225
R5566 VDDD.n1117 VDDD.n1116 2.03225
R5567 VDDD.n1132 VDDD.n1131 2.03225
R5568 VDDD.n1792 VDDD.n1791 2.03225
R5569 VDDD.n2624 VDDD.n2623 2.03225
R5570 VDDD.n2625 VDDD.n2624 2.03225
R5571 VDDD.n2076 VDDD.n2075 2.03225
R5572 VDDD.n3730 VDDD.n3729 2.03225
R5573 VDDD.n522 VDDD.n521 2.02422
R5574 VDDD.n292 VDDD.n290 2.01703
R5575 VDDD.n3352 VDDD.n3350 2.01703
R5576 VDDD.n1934 VDDD.n1932 2.01703
R5577 VDDD.n3657 VDDD.n3656 2.01042
R5578 VDDD.n3229 VDDD.n3228 2.01042
R5579 VDDD.n1842 VDDD.n1822 2.01042
R5580 VDDD.n1755 VDDD.n1754 2.01042
R5581 VDDD.n2445 VDDD.n2440 2.01042
R5582 VDDD.n2109 VDDD.n2107 2.01042
R5583 VDDD.n2168 VDDD.n2041 2.01042
R5584 VDDD.n2315 VDDD.n2314 2.01042
R5585 VDDD.n2975 VDDD.n1134 1.89415
R5586 VDDD.n291 VDDD.n290 1.88416
R5587 VDDD.n3351 VDDD.n3350 1.88416
R5588 VDDD.n1933 VDDD.n1932 1.88416
R5589 VDDD.n1001 VDDD.n1000 1.88285
R5590 VDDD.n2816 VDDD.n2813 1.88285
R5591 VDDD.n2912 VDDD.n2911 1.88285
R5592 VDDD.n2906 VDDD.n2905 1.88285
R5593 VDDD.n2597 VDDD.n2596 1.88285
R5594 VDDD.n2681 VDDD.n1573 1.88285
R5595 VDDD.n2650 VDDD.n2649 1.88285
R5596 VDDD.n2644 VDDD.n2643 1.88285
R5597 VDDD.n2457 VDDD.n2456 1.88285
R5598 VDDD.n516 VDDD.n515 1.82184
R5599 VDDD.n2219 VDDD.n2218 1.81289
R5600 VDDD.n2302 VDDD.n2301 1.81289
R5601 VDDD.n3256 VDDD.n3255 1.77828
R5602 VDDD.n1387 VDDD.n1386 1.77828
R5603 VDDD.n253 VDDD.n252 1.76897
R5604 VDDD.n2695 VDDD.n2694 1.76897
R5605 VDDD.n2146 VDDD.n2055 1.73737
R5606 VDDD.n1735 VDDD.n1733 1.69306
R5607 VDDD.n2211 VDDD.n1633 1.69188
R5608 VDDD.n2208 VDDD.n1633 1.69188
R5609 VDDD.n2582 VDDD.n1632 1.69188
R5610 VDDD.n2582 VDDD.n2581 1.69188
R5611 VDDD.n2964 VDDD.n1236 1.69188
R5612 VDDD.n2964 VDDD.n2963 1.69188
R5613 VDDD.n2965 VDDD.n1235 1.69188
R5614 VDDD.n2966 VDDD.n2965 1.69188
R5615 VDDD.n1005 VDDD.n564 1.69188
R5616 VDDD.n901 VDDD.n564 1.69188
R5617 VDDD.n3276 VDDD.n563 1.69188
R5618 VDDD.n3276 VDDD.n3275 1.69188
R5619 VDDD.n3412 VDDD.n341 1.69188
R5620 VDDD.n3319 VDDD.n341 1.69188
R5621 VDDD.n3625 VDDD.n3624 1.69188
R5622 VDDD.n3624 VDDD.n3623 1.69188
R5623 VDDD.n3767 VDDD.n3764 1.69188
R5624 VDDD.n3764 VDDD.n3763 1.69188
R5625 VDDD.n2583 VDDD.n1582 1.69188
R5626 VDDD.n2156 VDDD.n2155 1.69188
R5627 VDDD.n2155 VDDD.n2154 1.69188
R5628 VDDD.n2707 VDDD.n1563 1.69188
R5629 VDDD.n2707 VDDD.n2706 1.69188
R5630 VDDD.n2852 VDDD.n1095 1.69188
R5631 VDDD.n2798 VDDD.n1095 1.69188
R5632 VDDD.n3017 VDDD.n1094 1.69188
R5633 VDDD.n3017 VDDD.n3016 1.69188
R5634 VDDD.n1048 VDDD.n626 1.69188
R5635 VDDD.n868 VDDD.n626 1.69188
R5636 VDDD.n3165 VDDD.n3164 1.69188
R5637 VDDD.n3164 VDDD.n3163 1.69188
R5638 VDDD.n3471 VDDD.n361 1.69188
R5639 VDDD.n3471 VDDD.n3470 1.69188
R5640 VDDD.n3575 VDDD.n3574 1.69188
R5641 VDDD.n3574 VDDD.n3573 1.69188
R5642 VDDD.n3723 VDDD.n3722 1.69188
R5643 VDDD.n3722 VDDD.n3721 1.69188
R5644 VDDD.n2427 VDDD.n1564 1.69188
R5645 VDDD.n2381 VDDD.n2377 1.69188
R5646 VDDD.n2377 VDDD.n2376 1.69188
R5647 VDDD.n1882 VDDD.n1678 1.69188
R5648 VDDD.n1882 VDDD.n1881 1.69188
R5649 VDDD.n2758 VDDD.n2757 1.69188
R5650 VDDD.n2757 VDDD.n2756 1.69188
R5651 VDDD.n1422 VDDD.n1092 1.69188
R5652 VDDD.n1425 VDDD.n1092 1.69188
R5653 VDDD.n3022 VDDD.n1091 1.69188
R5654 VDDD.n3023 VDDD.n3022 1.69188
R5655 VDDD.n3118 VDDD.n561 1.69188
R5656 VDDD.n3115 VDDD.n561 1.69188
R5657 VDDD.n3282 VDDD.n560 1.69188
R5658 VDDD.n3283 VDDD.n3282 1.69188
R5659 VDDD.n3522 VDDD.n113 1.69188
R5660 VDDD.n3519 VDDD.n113 1.69188
R5661 VDDD.n3694 VDDD.n112 1.69188
R5662 VDDD.n3695 VDDD.n3694 1.69188
R5663 VDDD.n2099 VDDD.n1883 1.69188
R5664 VDDD.n2335 VDDD.n1959 1.69188
R5665 VDDD.n2335 VDDD.n2334 1.69188
R5666 VDDD.n2336 VDDD.n1958 1.69188
R5667 VDDD.n2337 VDDD.n2336 1.69188
R5668 VDDD.n1766 VDDD.n1561 1.69188
R5669 VDDD.n1769 VDDD.n1561 1.69188
R5670 VDDD.n2712 VDDD.n1560 1.69188
R5671 VDDD.n2713 VDDD.n2712 1.69188
R5672 VDDD.n1517 VDDD.n1321 1.69188
R5673 VDDD.n1517 VDDD.n1516 1.69188
R5674 VDDD.n3074 VDDD.n748 1.69188
R5675 VDDD.n3074 VDDD.n3073 1.69188
R5676 VDDD.n3075 VDDD.n747 1.69188
R5677 VDDD.n3076 VDDD.n3075 1.69188
R5678 VDDD.n444 VDDD.n207 1.69188
R5679 VDDD.n435 VDDD.n207 1.69188
R5680 VDDD.n3688 VDDD.n206 1.69188
R5681 VDDD.n3688 VDDD.n3687 1.69188
R5682 VDDD.n205 VDDD.n114 1.69188
R5683 VDDD.t1702 VDDD.t239 1.67895
R5684 VDDD.t656 VDDD.n3292 1.67895
R5685 VDDD.t1201 VDDD.t1207 1.67895
R5686 VDDD VDDD.t1959 1.67895
R5687 VDDD.t931 VDDD.t243 1.67895
R5688 VDDD VDDD.t1678 1.67895
R5689 VDDD.t295 VDDD 1.67895
R5690 VDDD.t381 VDDD.t949 1.67895
R5691 VDDD VDDD.t309 1.67895
R5692 VDDD.t666 VDDD.t267 1.67895
R5693 VDDD.n2218 VDDD.n2026 1.66186
R5694 VDDD.n2301 VDDD.n2300 1.66186
R5695 VDDD.n258 VDDD.n233 1.53093
R5696 VDDD.n475 VDDD.n474 1.52431
R5697 VDDD.n540 VDDD.n539 1.51829
R5698 VDDD.n2142 VDDD.n2055 1.51082
R5699 VDDD.n322 VDDD.n320 1.50638
R5700 VDDD.n329 VDDD.n328 1.50638
R5701 VDDD.n3590 VDDD.n350 1.50638
R5702 VDDD.n3583 VDDD.n355 1.50638
R5703 VDDD.n3428 VDDD.n3427 1.50638
R5704 VDDD.n3420 VDDD.n3419 1.50638
R5705 VDDD.n1083 VDDD.n1082 1.50638
R5706 VDDD.n1458 VDDD.n1456 1.50638
R5707 VDDD.n1464 VDDD.n1454 1.50638
R5708 VDDD.n2746 VDDD.n2745 1.50638
R5709 VDDD.n2733 VDDD.n2732 1.50638
R5710 VDDD.n2353 VDDD.n1902 1.50638
R5711 VDDD.n2475 VDDD.n2474 1.50638
R5712 VDDD.n2369 VDDD.n2368 1.50638
R5713 VDDD.n2362 VDDD.n1887 1.50638
R5714 VDDD.n549 VDDD.n548 1.47352
R5715 VDDD.n409 VDDD.n397 1.47352
R5716 VDDD.n1476 VDDD.n1475 1.47352
R5717 VDDD.n2084 VDDD.n2074 1.47352
R5718 VDDD.n1876 VDDD.n1807 1.46336
R5719 VDDD.n1118 VDDD.n1117 1.42272
R5720 VDDD.n3000 VDDD.n2999 1.42272
R5721 VDDD.n238 VDDD.n216 1.37571
R5722 VDDD.n424 VDDD.n389 1.37571
R5723 VDDD.n721 VDDD.n720 1.37571
R5724 VDDD.n3207 VDDD.n3206 1.37571
R5725 VDDD.n789 VDDD.n758 1.37571
R5726 VDDD.n1152 VDDD.n1151 1.37571
R5727 VDDD.n1778 VDDD.n1707 1.37571
R5728 VDDD.n2130 VDDD.n2129 1.37571
R5729 VDDD.n2012 VDDD.n1998 1.37571
R5730 VDDD.n1938 VDDD.n1936 1.26517
R5731 VDDD.n288 VDDD.n287 1.2502
R5732 VDDD.n498 VDDD.n496 1.2502
R5733 VDDD.n3303 VDDD.n3301 1.2502
R5734 VDDD.n3348 VDDD.n3344 1.2502
R5735 VDDD.n639 VDDD.n637 1.2502
R5736 VDDD.n807 VDDD.n805 1.2502
R5737 VDDD.n1338 VDDD.n1335 1.2502
R5738 VDDD.n1657 VDDD.n1655 1.2502
R5739 VDDD.n3643 VDDD.n3641 1.2395
R5740 VDDD.n3604 VDDD.n3603 1.16678
R5741 VDDD.n2189 VDDD.n2188 1.16678
R5742 VDDD.n793 VDDD.n792 1.15996
R5743 VDDD.n1742 VDDD.n1741 1.1546
R5744 VDDD.n815 VDDD.n812 1.12991
R5745 VDDD.n1429 VDDD.n1346 1.12991
R5746 VDDD.n1939 VDDD.n1938 1.11173
R5747 VDDD.n955 VDDD.n954 1.11123
R5748 VDDD.n237 VDDD.n234 0.992049
R5749 VDDD.n254 VDDD.n233 0.992049
R5750 VDDD.n1598 VDDD.n1570 0.992049
R5751 VDDD.n2696 VDDD.n1569 0.992049
R5752 VDDD.n2420 VDDD.n2419 0.965579
R5753 VDDD.n3002 VDDD.n1118 0.914786
R5754 VDDD.n1986 VDDD.n1982 0.899674
R5755 VDDD.n3829 VDDD.n3828 0.863992
R5756 VDDD.n51 VDDD.n50 0.863992
R5757 VDDD.n142 VDDD.n141 0.863992
R5758 VDDD.n133 VDDD.n132 0.863992
R5759 VDDD.n2131 VDDD.n2058 0.846781
R5760 VDDD.n308 VDDD.n307 0.753441
R5761 VDDD.n326 VDDD.n272 0.753441
R5762 VDDD.n3564 VDDD.n3563 0.753441
R5763 VDDD.n3535 VDDD.n3534 0.753441
R5764 VDDD.n3367 VDDD.n3366 0.753441
R5765 VDDD.n3392 VDDD.n3330 0.753441
R5766 VDDD.n3433 VDDD.n3305 0.753441
R5767 VDDD.n3419 VDDD.n3418 0.753441
R5768 VDDD.n463 VDDD.n462 0.753441
R5769 VDDD.n657 VDDD.n654 0.753441
R5770 VDDD.n3080 VDDD.n689 0.753441
R5771 VDDD.n3044 VDDD.n3043 0.753441
R5772 VDDD.n3039 VDDD.n3038 0.753441
R5773 VDDD.n1072 VDDD.n847 0.753441
R5774 VDDD.n1028 VDDD.n882 0.753441
R5775 VDDD.n906 VDDD.n893 0.753441
R5776 VDDD.n959 VDDD.n931 0.753441
R5777 VDDD.n1497 VDDD.n1334 0.753441
R5778 VDDD.n1462 VDDD.n1461 0.753441
R5779 VDDD.n3007 VDDD.n3006 0.753441
R5780 VDDD.n2994 VDDD.n1125 0.753441
R5781 VDDD.n2820 VDDD.n2816 0.753441
R5782 VDDD.n2826 VDDD.n2812 0.753441
R5783 VDDD.n2750 VDDD.n2749 0.753441
R5784 VDDD.n2729 VDDD.n2728 0.753441
R5785 VDDD.n1850 VDDD.n1817 0.753441
R5786 VDDD.n1610 VDDD.n1609 0.753441
R5787 VDDD.n2594 VDDD.n1576 0.753441
R5788 VDDD.n2351 VDDD.n2350 0.753441
R5789 VDDD.n2409 VDDD.n2408 0.753441
R5790 VDDD.n2371 VDDD.n1673 0.753441
R5791 VDDD.n3742 VDDD.n3741 0.753441
R5792 VDDD.n1412 VDDD.n1367 0.731929
R5793 VDDD.n1875 VDDD.n1809 0.731929
R5794 VDDD.n1472 VDDD.n1450 0.660817
R5795 VDDD.n526 VDDD.n525 0.658208
R5796 VDDD.n579 VDDD.n578 0.651997
R5797 VDDD.n787 VDDD.n786 0.651997
R5798 VDDD.n3806 VDDD.n7 0.635211
R5799 VDDD.n3822 VDDD.n1 0.635211
R5800 VDDD.n3786 VDDD.n14 0.635211
R5801 VDDD.n3805 VDDD.n8 0.635211
R5802 VDDD.n3605 VDDD.n3604 0.635211
R5803 VDDD.n3614 VDDD.n338 0.635211
R5804 VDDD.n3631 VDDD.n3630 0.635211
R5805 VDDD.n3641 VDDD.n334 0.635211
R5806 VDDD.n242 VDDD.n241 0.635211
R5807 VDDD.n3662 VDDD.n3661 0.635211
R5808 VDDD.n224 VDDD.n222 0.635211
R5809 VDDD.n3504 VDDD.n229 0.635211
R5810 VDDD.n3510 VDDD.n3498 0.635211
R5811 VDDD.n421 VDDD.n420 0.635211
R5812 VDDD.n454 VDDD.n378 0.635211
R5813 VDDD.n720 VDDD.n718 0.635211
R5814 VDDD.n3123 VDDD.n658 0.635211
R5815 VDDD.n3222 VDDD.n3221 0.635211
R5816 VDDD.n3218 VDDD.n3179 0.635211
R5817 VDDD.n3196 VDDD.n3187 0.635211
R5818 VDDD.n791 VDDD.n790 0.635211
R5819 VDDD.n3046 VDDD.n765 0.635211
R5820 VDDD.n2975 VDDD.n2974 0.635211
R5821 VDDD.n1224 VDDD.n1223 0.635211
R5822 VDDD.n1219 VDDD.n1156 0.635211
R5823 VDDD.n1821 VDDD.n1819 0.635211
R5824 VDDD.n1759 VDDD.n1728 0.635211
R5825 VDDD.n1784 VDDD.n1704 0.635211
R5826 VDDD.n1761 VDDD.n1760 0.635211
R5827 VDDD.n2448 VDDD.n2447 0.635211
R5828 VDDD.n2125 VDDD.n2061 0.635211
R5829 VDDD.n2141 VDDD.n2056 0.635211
R5830 VDDD.n2124 VDDD.n2062 0.635211
R5831 VDDD.n2165 VDDD.n2164 0.635211
R5832 VDDD.n2186 VDDD.n2034 0.635211
R5833 VDDD.n2190 VDDD.n2189 0.635211
R5834 VDDD.n2199 VDDD.n2028 0.635211
R5835 VDDD.n2016 VDDD.n2015 0.635211
R5836 VDDD.n2319 VDDD.n1969 0.635211
R5837 VDDD.n2318 VDDD.n1970 0.635211
R5838 VDDD.n94 VDDD.n72 0.635211
R5839 VDDD.n3716 VDDD.n46 0.635211
R5840 VDDD.n3699 VDDD.n52 0.635211
R5841 VDDD.n95 VDDD.n71 0.635211
R5842 VDDD.n197 VDDD.n172 0.635211
R5843 VDDD.n178 VDDD.n48 0.635211
R5844 VDDD.n147 VDDD.n125 0.635211
R5845 VDDD.n199 VDDD.n198 0.635211
R5846 VDDD.n1737 VDDD.n1689 0.630008
R5847 VDDD.n2414 VDDD.n1662 0.629194
R5848 VDDD.n3299 VDDD.n3298 0.597579
R5849 VDDD.n511 VDDD.n510 0.568305
R5850 VDDD.n1475 VDDD.n1474 0.55923
R5851 VDDD.n3269 VDDD.n3267 0.5532
R5852 VDDD.n1391 VDDD.n1385 0.5532
R5853 VDDD.n3692 VDDD.n3689 0.551088
R5854 VDDD.n2711 VDDD.n2710 0.551088
R5855 VDDD.n3020 VDDD.n749 0.551088
R5856 VDDD.n3280 VDDD.n562 0.551088
R5857 VDDD.n3612 VDDD.n3611 0.529426
R5858 VDDD.n3201 VDDD.n3200 0.529426
R5859 VDDD.n1228 VDDD.n1153 0.529426
R5860 VDDD.n2137 VDDD.n2136 0.529426
R5861 VDDD.n2197 VDDD.n2196 0.529426
R5862 VDDD.n3257 VDDD.n3256 0.457643
R5863 VDDD.n3635 VDDD.n336 0.42364
R5864 VDDD.n3509 VDDD.n3508 0.42364
R5865 VDDD.n2089 VDDD.n2086 0.42364
R5866 VDDD.n3278 VDDD.n3277 0.3805
R5867 VDDD.n1142 VDDD.n1093 0.3805
R5868 VDDD.n1562 VDDD.n1237 0.3805
R5869 VDDD.n3690 VDDD.n26 0.3805
R5870 VDDD.n3279 VDDD.n362 0.3805
R5871 VDDD.n3019 VDDD.n3018 0.3805
R5872 VDDD.n2709 VDDD.n2708 0.3805
R5873 VDDD.n3691 VDDD.n41 0.3805
R5874 VDDD.n3281 VDDD.n3280 0.3805
R5875 VDDD.n3021 VDDD.n3020 0.3805
R5876 VDDD.n2710 VDDD.n1281 0.3805
R5877 VDDD.n3693 VDDD.n3692 0.3805
R5878 VDDD.n1218 VDDD.n1157 0.369731
R5879 VDDD.n1199 VDDD.n1163 0.369731
R5880 VDDD.n1198 VDDD.n1164 0.369731
R5881 VDDD.n1179 VDDD.n1170 0.369731
R5882 VDDD.n2555 VDDD.n2494 0.369731
R5883 VDDD.n2536 VDDD.n2500 0.369731
R5884 VDDD.n2535 VDDD.n2501 0.369731
R5885 VDDD.n2516 VDDD.n2507 0.369731
R5886 VDDD.n2290 VDDD.n2229 0.369731
R5887 VDDD.n2271 VDDD.n2235 0.369731
R5888 VDDD.n2270 VDDD.n2236 0.369731
R5889 VDDD.n2251 VDDD.n2242 0.369731
R5890 VDDD.n1785 VDDD.n1784 0.32333
R5891 VDDD.n3364 VDDD.n3346 0.317568
R5892 VDDD.n642 VDDD.n641 0.317568
R5893 VDDD.n3346 VDDD.n3345 0.316929
R5894 VDDD.n641 VDDD.n640 0.316929
R5895 VDDD.n3828 VDDD.n3827 0.305262
R5896 VDDD.n250 VDDD.n249 0.305262
R5897 VDDD.n549 VDDD.n501 0.305262
R5898 VDDD.n3436 VDDD.n3304 0.305262
R5899 VDDD.n3407 VDDD.n3406 0.305262
R5900 VDDD.n3405 VDDD.n3326 0.305262
R5901 VDDD.n410 VDDD.n409 0.305262
R5902 VDDD.n413 VDDD.n412 0.305262
R5903 VDDD.n470 VDDD.n469 0.305262
R5904 VDDD.n473 VDDD.n371 0.305262
R5905 VDDD.n3098 VDDD.n669 0.305262
R5906 VDDD.n3094 VDDD.n680 0.305262
R5907 VDDD.n3091 VDDD.n681 0.305262
R5908 VDDD.n611 VDDD.n582 0.305262
R5909 VDDD.n3267 VDDD.n571 0.305262
R5910 VDDD.n3250 VDDD.n3249 0.305262
R5911 VDDD.n800 VDDD.n799 0.305262
R5912 VDDD.n793 VDDD.n788 0.305262
R5913 VDDD.n1043 VDDD.n873 0.305262
R5914 VDDD.n1033 VDDD.n1032 0.305262
R5915 VDDD.n914 VDDD.n911 0.305262
R5916 VDDD.n984 VDDD.n983 0.305262
R5917 VDDD.n954 VDDD.n935 0.305262
R5918 VDDD.n948 VDDD.n947 0.305262
R5919 VDDD.n1477 VDDD.n1476 0.305262
R5920 VDDD.n1469 VDDD.n1451 0.305262
R5921 VDDD.n1391 VDDD.n1390 0.305262
R5922 VDDD.n3011 VDDD.n1100 0.305262
R5923 VDDD.n1484 VDDD.n1340 0.305262
R5924 VDDD.n1116 VDDD.n1113 0.305262
R5925 VDDD.n2999 VDDD.n2998 0.305262
R5926 VDDD.n1131 VDDD.n1129 0.305262
R5927 VDDD.n2979 VDDD.n2978 0.305262
R5928 VDDD.n2818 VDDD.n2817 0.305262
R5929 VDDD.n2958 VDDD.n1243 0.305262
R5930 VDDD.n2786 VDDD.n2785 0.305262
R5931 VDDD.n2858 VDDD.n1253 0.305262
R5932 VDDD.n2904 VDDD.n2880 0.305262
R5933 VDDD.n2901 VDDD.n2881 0.305262
R5934 VDDD.n2895 VDDD.n2894 0.305262
R5935 VDDD.n1793 VDDD.n1792 0.305262
R5936 VDDD.n1702 VDDD.n1701 0.305262
R5937 VDDD.n1786 VDDD.n1703 0.305262
R5938 VDDD.n1602 VDDD.n1595 0.305262
R5939 VDDD.n2642 VDDD.n2623 0.305262
R5940 VDDD.n2639 VDDD.n2625 0.305262
R5941 VDDD.n2635 VDDD.n2626 0.305262
R5942 VDDD.n2490 VDDD.n1649 0.305262
R5943 VDDD.n2075 VDDD.n2074 0.305262
R5944 VDDD.n3729 VDDD.n3728 0.305262
R5945 VDDD.n3735 VDDD.n36 0.305262
R5946 VDDD.n50 VDDD.n47 0.305262
R5947 VDDD.n3701 VDDD.n3700 0.305262
R5948 VDDD.n141 VDDD.n140 0.305262
R5949 VDDD.n146 VDDD.n126 0.305262
R5950 VDDD.n132 VDDD.n130 0.305262
R5951 VDDD.n535 VDDD.n516 0.304057
R5952 VDDD.n529 VDDD.n521 0.304057
R5953 VDDD.n3465 VDDD.n367 0.304057
R5954 VDDD.n3443 VDDD.n3442 0.297291
R5955 VDDD.n1492 VDDD.n1491 0.297291
R5956 VDDD.n252 VDDD 0.2951
R5957 VDDD.n2694 VDDD 0.2951
R5958 VDDD.n3690 VDDD 0.282994
R5959 VDDD.n1562 VDDD 0.282994
R5960 VDDD.n1093 VDDD 0.282994
R5961 VDDD.n3278 VDDD 0.282994
R5962 VDDD.n252 VDDD 0.256072
R5963 VDDD.n2694 VDDD 0.256072
R5964 VDDD.n3324 VDDD.n3313 0.254468
R5965 VDDD.n3254 VDDD.n574 0.254468
R5966 VDDD.n951 VDDD.n950 0.254468
R5967 VDDD.n546 VDDD.n545 0.239381
R5968 VDDD VDDD.n303 0.238178
R5969 VDDD VDDD.n3443 0.238178
R5970 VDDD.n3363 VDDD 0.238178
R5971 VDDD.n3149 VDDD 0.238178
R5972 VDDD.n619 VDDD 0.238178
R5973 VDDD.n802 VDDD 0.238178
R5974 VDDD.n1492 VDDD 0.238178
R5975 VDDD VDDD.n1942 0.238178
R5976 VDDD VDDD.n302 0.237784
R5977 VDDD VDDD.n3362 0.237784
R5978 VDDD.n3363 VDDD 0.237395
R5979 VDDD VDDD.n3149 0.237395
R5980 VDDD.n2564 VDDD.n2563 0.227049
R5981 VDDD.n2558 VDDD.n1644 0.227049
R5982 VDDD.n2143 VDDD.n2142 0.227049
R5983 VDDD.n2149 VDDD.n2148 0.227049
R5984 VDDD.n2217 VDDD.n2216 0.227049
R5985 VDDD.n2226 VDDD.n2225 0.227049
R5986 VDDD.n1977 VDDD.n1975 0.227049
R5987 VDDD.n2296 VDDD.n1978 0.227049
R5988 VDDD.n3463 VDDD.n3462 0.22119
R5989 VDDD.n1177 VDDD 0.217591
R5990 VDDD.n2514 VDDD 0.217591
R5991 VDDD.n2249 VDDD 0.217591
R5992 VDDD.n3651 VDDD.n3650 0.21207
R5993 VDDD.n727 VDDD.n724 0.21207
R5994 VDDD.n3109 VDDD.n665 0.21207
R5995 VDDD.n3235 VDDD.n3234 0.21207
R5996 VDDD.n1837 VDDD.n1826 0.21207
R5997 VDDD.n1749 VDDD.n1748 0.21207
R5998 VDDD.n2576 VDDD.n2575 0.21207
R5999 VDDD.n2090 VDDD.n2089 0.21207
R6000 VDDD.n2309 VDDD.n2308 0.21207
R6001 VDDD.n246 VDDD.n245 0.203675
R6002 VDDD.n3400 VDDD.n3399 0.203675
R6003 VDDD.n414 VDDD.n391 0.203675
R6004 VDDD.n797 VDDD.n796 0.203675
R6005 VDDD.n302 VDDD 0.200023
R6006 VDDD.n3362 VDDD 0.200023
R6007 VDDD.n303 VDDD 0.199635
R6008 VDDD.n619 VDDD 0.199635
R6009 VDDD.n802 VDDD 0.199635
R6010 VDDD.n1942 VDDD 0.199635
R6011 VDDD.n3011 VDDD.n3010 0.192069
R6012 VDDD.n1399 VDDD.n1374 0.180304
R6013 VDDD.n1381 VDDD.n1374 0.180304
R6014 VDDD.n3453 VDDD.n3295 0.180304
R6015 VDDD.n299 VDDD 0.17983
R6016 VDDD.n3359 VDDD 0.17983
R6017 VDDD.n3194 VDDD 0.17983
R6018 VDDD VDDD.n945 0.17983
R6019 VDDD.n2892 VDDD 0.17983
R6020 VDDD.n2633 VDDD 0.17983
R6021 VDDD.n3287 VDDD 0.17983
R6022 VDDD VDDD.n546 0.17983
R6023 VDDD.n3239 VDDD 0.17983
R6024 VDDD.n304 VDDD 0.179485
R6025 VDDD VDDD.n2018 0.179485
R6026 VDDD.n262 VDDD 0.172576
R6027 VDDD VDDD.n405 0.172576
R6028 VDDD VDDD.n677 0.172576
R6029 VDDD VDDD.n782 0.172576
R6030 VDDD VDDD.n1446 0.172576
R6031 VDDD VDDD.n1304 0.172576
R6032 VDDD VDDD.n1698 0.172576
R6033 VDDD VDDD.n1897 0.172576
R6034 VDDD VDDD.n1994 0.172576
R6035 VDDD.n3692 VDDD.n3691 0.171088
R6036 VDDD.n3691 VDDD.n3690 0.171088
R6037 VDDD.n2710 VDDD.n2709 0.171088
R6038 VDDD.n2709 VDDD.n1562 0.171088
R6039 VDDD.n3020 VDDD.n3019 0.171088
R6040 VDDD.n3019 VDDD.n1093 0.171088
R6041 VDDD.n3280 VDDD.n3279 0.171088
R6042 VDDD.n3279 VDDD.n3278 0.171088
R6043 VDDD.n1830 VDDD.n1566 0.167283
R6044 VDDD.n1535 VDDD.n1533 0.163904
R6045 VDDD.n1536 VDDD.n1293 0.163904
R6046 VDDD VDDD.n2043 0.158169
R6047 VDDD.n3624 VDDD.n341 0.1509
R6048 VDDD.n3276 VDDD.n564 0.1509
R6049 VDDD.n2965 VDDD.n2964 0.1509
R6050 VDDD.n2583 VDDD.n2582 0.1509
R6051 VDDD.n2582 VDDD.n1633 0.1509
R6052 VDDD.n3574 VDDD.n3471 0.1509
R6053 VDDD.n3164 VDDD.n626 0.1509
R6054 VDDD.n3017 VDDD.n1095 0.1509
R6055 VDDD.n2707 VDDD.n1564 0.1509
R6056 VDDD.n2155 VDDD.n1564 0.1509
R6057 VDDD.n3282 VDDD.n113 0.1509
R6058 VDDD.n3022 VDDD.n561 0.1509
R6059 VDDD.n2757 VDDD.n1092 0.1509
R6060 VDDD.n2377 VDDD.n1882 0.1509
R6061 VDDD.n2377 VDDD.n1883 0.1509
R6062 VDDD.n3688 VDDD.n207 0.1509
R6063 VDDD.n3075 VDDD.n3074 0.1509
R6064 VDDD.n2712 VDDD.n1517 0.1509
R6065 VDDD.n2336 VDDD.n1561 0.1509
R6066 VDDD.n2336 VDDD.n2335 0.1509
R6067 VDDD.n304 VDDD 0.14207
R6068 VDDD.n2018 VDDD 0.14207
R6069 VDDD.n299 VDDD 0.141725
R6070 VDDD.n3287 VDDD 0.141725
R6071 VDDD.n3359 VDDD 0.141725
R6072 VDDD.n3239 VDDD 0.141725
R6073 VDDD.n3194 VDDD 0.141725
R6074 VDDD.n945 VDDD 0.141725
R6075 VDDD.n1177 VDDD 0.141725
R6076 VDDD.n2892 VDDD 0.141725
R6077 VDDD.n2633 VDDD 0.141725
R6078 VDDD.n2514 VDDD 0.141725
R6079 VDDD.n2249 VDDD 0.141725
R6080 VDDD.n3764 VDDD.n26 0.139565
R6081 VDDD.n3722 VDDD.n41 0.139565
R6082 VDDD.n3694 VDDD.n3693 0.139565
R6083 VDDD.n3689 VDDD.n205 0.139565
R6084 VDDD VDDD.n1941 0.120408
R6085 VDDD VDDD.n781 0.120408
R6086 VDDD.n1830 VDDD 0.120408
R6087 VDDD VDDD.n1659 0.120408
R6088 VDDD.n251 VDDD.n235 0.120292
R6089 VDDD.n244 VDDD.n235 0.120292
R6090 VDDD.n3673 VDDD.n3672 0.120292
R6091 VDDD.n3672 VDDD.n3671 0.120292
R6092 VDDD.n3671 VDDD.n218 0.120292
R6093 VDDD.n3666 VDDD.n218 0.120292
R6094 VDDD.n3666 VDDD.n3665 0.120292
R6095 VDDD.n3665 VDDD.n221 0.120292
R6096 VDDD.n3660 VDDD.n221 0.120292
R6097 VDDD.n3659 VDDD.n3658 0.120292
R6098 VDDD.n3658 VDDD.n223 0.120292
R6099 VDDD.n3653 VDDD.n223 0.120292
R6100 VDDD.n3653 VDDD.n3652 0.120292
R6101 VDDD.n3652 VDDD.n226 0.120292
R6102 VDDD.n3506 VDDD.n3505 0.120292
R6103 VDDD.n3506 VDDD.n3503 0.120292
R6104 VDDD.n3513 VDDD.n3503 0.120292
R6105 VDDD.n3532 VDDD.n3531 0.120292
R6106 VDDD.n3533 VDDD.n3532 0.120292
R6107 VDDD.n3533 VDDD.n3494 0.120292
R6108 VDDD.n3494 VDDD.n3492 0.120292
R6109 VDDD.n3539 VDDD.n3492 0.120292
R6110 VDDD.n3540 VDDD.n3539 0.120292
R6111 VDDD.n3540 VDDD.n3489 0.120292
R6112 VDDD.n3544 VDDD.n3489 0.120292
R6113 VDDD.n3545 VDDD.n3544 0.120292
R6114 VDDD.n3546 VDDD.n3545 0.120292
R6115 VDDD.n3546 VDDD.n3486 0.120292
R6116 VDDD.n3552 VDDD.n3486 0.120292
R6117 VDDD.n3553 VDDD.n3552 0.120292
R6118 VDDD.n3554 VDDD.n3553 0.120292
R6119 VDDD.n3560 VDDD.n3483 0.120292
R6120 VDDD.n3561 VDDD.n3560 0.120292
R6121 VDDD.n3562 VDDD.n3561 0.120292
R6122 VDDD.n358 VDDD.n356 0.120292
R6123 VDDD.n356 VDDD.n353 0.120292
R6124 VDDD.n3584 VDDD.n353 0.120292
R6125 VDDD.n3585 VDDD.n3584 0.120292
R6126 VDDD.n3586 VDDD.n3585 0.120292
R6127 VDDD.n3586 VDDD.n351 0.120292
R6128 VDDD.n3592 VDDD.n351 0.120292
R6129 VDDD.n3593 VDDD.n3592 0.120292
R6130 VDDD.n3594 VDDD.n3593 0.120292
R6131 VDDD.n3594 VDDD.n348 0.120292
R6132 VDDD.n3598 VDDD.n348 0.120292
R6133 VDDD.n3599 VDDD.n3598 0.120292
R6134 VDDD.n3608 VDDD.n346 0.120292
R6135 VDDD.n3609 VDDD.n3608 0.120292
R6136 VDDD.n3610 VDDD.n3609 0.120292
R6137 VDDD.n3634 VDDD.n3633 0.120292
R6138 VDDD.n3634 VDDD.n335 0.120292
R6139 VDDD.n3639 VDDD.n335 0.120292
R6140 VDDD.n3640 VDDD.n3639 0.120292
R6141 VDDD.n332 VDDD.n331 0.120292
R6142 VDDD.n331 VDDD.n271 0.120292
R6143 VDDD.n325 VDDD.n271 0.120292
R6144 VDDD.n325 VDDD.n324 0.120292
R6145 VDDD.n324 VDDD.n273 0.120292
R6146 VDDD.n317 VDDD.n273 0.120292
R6147 VDDD.n317 VDDD.n316 0.120292
R6148 VDDD.n316 VDDD.n315 0.120292
R6149 VDDD.n315 VDDD.n275 0.120292
R6150 VDDD.n311 VDDD.n275 0.120292
R6151 VDDD.n311 VDDD.n310 0.120292
R6152 VDDD.n310 VDDD.n309 0.120292
R6153 VDDD.n309 VDDD.n277 0.120292
R6154 VDDD.n417 VDDD.n392 0.120292
R6155 VDDD.n418 VDDD.n417 0.120292
R6156 VDDD.n419 VDDD.n390 0.120292
R6157 VDDD.n425 VDDD.n390 0.120292
R6158 VDDD.n426 VDDD.n425 0.120292
R6159 VDDD.n426 VDDD.n387 0.120292
R6160 VDDD.n433 VDDD.n387 0.120292
R6161 VDDD.n452 VDDD.n379 0.120292
R6162 VDDD.n453 VDDD.n452 0.120292
R6163 VDDD.n457 VDDD.n377 0.120292
R6164 VDDD.n458 VDDD.n457 0.120292
R6165 VDDD.n459 VDDD.n458 0.120292
R6166 VDDD.n459 VDDD.n374 0.120292
R6167 VDDD.n466 VDDD.n374 0.120292
R6168 VDDD.n468 VDDD.n372 0.120292
R6169 VDDD.n476 VDDD.n372 0.120292
R6170 VDDD.n477 VDDD.n476 0.120292
R6171 VDDD.n557 VDDD.n556 0.120292
R6172 VDDD.n556 VDDD.n495 0.120292
R6173 VDDD.n551 VDDD.n550 0.120292
R6174 VDDD.n545 VDDD.n508 0.120292
R6175 VDDD.n538 VDDD.n508 0.120292
R6176 VDDD.n538 VDDD.n537 0.120292
R6177 VDDD.n537 VDDD.n536 0.120292
R6178 VDDD.n532 VDDD.n519 0.120292
R6179 VDDD.n528 VDDD.n527 0.120292
R6180 VDDD.n3442 VDDD.n3300 0.120292
R6181 VDDD.n3438 VDDD.n3300 0.120292
R6182 VDDD.n3438 VDDD.n3437 0.120292
R6183 VDDD.n3431 VDDD.n3306 0.120292
R6184 VDDD.n3424 VDDD.n3307 0.120292
R6185 VDDD.n3424 VDDD.n3423 0.120292
R6186 VDDD.n3423 VDDD.n3422 0.120292
R6187 VDDD.n3409 VDDD.n3323 0.120292
R6188 VDDD.n3404 VDDD.n3403 0.120292
R6189 VDDD.n3403 VDDD.n3327 0.120292
R6190 VDDD.n3393 VDDD.n3331 0.120292
R6191 VDDD.n3388 VDDD.n3331 0.120292
R6192 VDDD.n3388 VDDD.n3387 0.120292
R6193 VDDD.n3387 VDDD.n3386 0.120292
R6194 VDDD.n3386 VDDD.n3334 0.120292
R6195 VDDD.n3382 VDDD.n3334 0.120292
R6196 VDDD.n3382 VDDD.n3381 0.120292
R6197 VDDD.n3381 VDDD.n3337 0.120292
R6198 VDDD.n3375 VDDD.n3337 0.120292
R6199 VDDD.n3375 VDDD.n3374 0.120292
R6200 VDDD.n3374 VDDD.n3373 0.120292
R6201 VDDD.n3373 VDDD.n3339 0.120292
R6202 VDDD.n3369 VDDD.n3339 0.120292
R6203 VDDD.n3369 VDDD.n3368 0.120292
R6204 VDDD.n3368 VDDD.n3342 0.120292
R6205 VDDD.n3093 VDDD.n3092 0.120292
R6206 VDDD.n3088 VDDD.n682 0.120292
R6207 VDDD.n3088 VDDD.n3087 0.120292
R6208 VDDD.n3084 VDDD.n3083 0.120292
R6209 VDDD.n3083 VDDD.n686 0.120292
R6210 VDDD.n3079 VDDD.n686 0.120292
R6211 VDDD.n744 VDDD.n696 0.120292
R6212 VDDD.n710 VDDD.n696 0.120292
R6213 VDDD.n739 VDDD.n710 0.120292
R6214 VDDD.n739 VDDD.n738 0.120292
R6215 VDDD.n738 VDDD.n737 0.120292
R6216 VDDD.n737 VDDD.n712 0.120292
R6217 VDDD.n717 VDDD.n712 0.120292
R6218 VDDD.n732 VDDD.n717 0.120292
R6219 VDDD.n731 VDDD.n730 0.120292
R6220 VDDD.n730 VDDD.n719 0.120292
R6221 VDDD.n726 VDDD.n719 0.120292
R6222 VDDD.n726 VDDD.n725 0.120292
R6223 VDDD.n3104 VDDD.n3103 0.120292
R6224 VDDD.n3127 VDDD.n3126 0.120292
R6225 VDDD.n3127 VDDD.n652 0.120292
R6226 VDDD.n3134 VDDD.n652 0.120292
R6227 VDDD.n3135 VDDD.n3134 0.120292
R6228 VDDD.n3135 VDDD.n648 0.120292
R6229 VDDD.n3141 VDDD.n648 0.120292
R6230 VDDD.n3142 VDDD.n3141 0.120292
R6231 VDDD.n3143 VDDD.n3142 0.120292
R6232 VDDD.n3143 VDDD.n645 0.120292
R6233 VDDD.n645 VDDD.n643 0.120292
R6234 VDDD.n3151 VDDD.n3150 0.120292
R6235 VDDD.n614 VDDD.n613 0.120292
R6236 VDDD.n613 VDDD.n612 0.120292
R6237 VDDD.n607 VDDD.n584 0.120292
R6238 VDDD.n602 VDDD.n584 0.120292
R6239 VDDD.n602 VDDD.n601 0.120292
R6240 VDDD.n601 VDDD.n600 0.120292
R6241 VDDD.n600 VDDD.n587 0.120292
R6242 VDDD.n593 VDDD.n587 0.120292
R6243 VDDD.n594 VDDD.n593 0.120292
R6244 VDDD.n3259 VDDD.n573 0.120292
R6245 VDDD.n3253 VDDD.n573 0.120292
R6246 VDDD.n3253 VDDD.n3252 0.120292
R6247 VDDD.n3252 VDDD.n575 0.120292
R6248 VDDD.n3233 VDDD.n3232 0.120292
R6249 VDDD.n3232 VDDD.n3231 0.120292
R6250 VDDD.n3231 VDDD.n3176 0.120292
R6251 VDDD.n3226 VDDD.n3176 0.120292
R6252 VDDD.n3226 VDDD.n3225 0.120292
R6253 VDDD.n3225 VDDD.n3224 0.120292
R6254 VDDD.n3224 VDDD.n3178 0.120292
R6255 VDDD.n3217 VDDD.n3216 0.120292
R6256 VDDD.n3216 VDDD.n3180 0.120292
R6257 VDDD.n3211 VDDD.n3180 0.120292
R6258 VDDD.n3211 VDDD.n3210 0.120292
R6259 VDDD.n3210 VDDD.n3182 0.120292
R6260 VDDD.n3205 VDDD.n3182 0.120292
R6261 VDDD.n3205 VDDD.n3204 0.120292
R6262 VDDD.n3204 VDDD.n3203 0.120292
R6263 VDDD.n3203 VDDD.n3185 0.120292
R6264 VDDD.n3198 VDDD.n3185 0.120292
R6265 VDDD.n3198 VDDD.n3197 0.120292
R6266 VDDD.n801 VDDD.n785 0.120292
R6267 VDDD.n795 VDDD.n785 0.120292
R6268 VDDD.n795 VDDD.n794 0.120292
R6269 VDDD.n3060 VDDD.n3059 0.120292
R6270 VDDD.n3059 VDDD.n760 0.120292
R6271 VDDD.n3054 VDDD.n760 0.120292
R6272 VDDD.n3054 VDDD.n3053 0.120292
R6273 VDDD.n3053 VDDD.n3052 0.120292
R6274 VDDD.n3052 VDDD.n762 0.120292
R6275 VDDD.n3048 VDDD.n762 0.120292
R6276 VDDD.n3048 VDDD.n3047 0.120292
R6277 VDDD.n3042 VDDD.n3041 0.120292
R6278 VDDD.n3041 VDDD.n3040 0.120292
R6279 VDDD.n3040 VDDD.n769 0.120292
R6280 VDDD.n3032 VDDD.n813 0.120292
R6281 VDDD.n3026 VDDD.n813 0.120292
R6282 VDDD.n1088 VDDD.n826 0.120292
R6283 VDDD.n1081 VDDD.n826 0.120292
R6284 VDDD.n1081 VDDD.n1080 0.120292
R6285 VDDD.n1080 VDDD.n1079 0.120292
R6286 VDDD.n1076 VDDD.n1075 0.120292
R6287 VDDD.n1075 VDDD.n844 0.120292
R6288 VDDD.n1071 VDDD.n844 0.120292
R6289 VDDD.n1071 VDDD.n1070 0.120292
R6290 VDDD.n1070 VDDD.n848 0.120292
R6291 VDDD.n1066 VDDD.n848 0.120292
R6292 VDDD.n1066 VDDD.n1065 0.120292
R6293 VDDD.n1065 VDDD.n852 0.120292
R6294 VDDD.n853 VDDD.n852 0.120292
R6295 VDDD.n1060 VDDD.n853 0.120292
R6296 VDDD.n1060 VDDD.n1059 0.120292
R6297 VDDD.n1059 VDDD.n1058 0.120292
R6298 VDDD.n1058 VDDD.n855 0.120292
R6299 VDDD.n1042 VDDD.n1041 0.120292
R6300 VDDD.n1041 VDDD.n874 0.120292
R6301 VDDD.n1035 VDDD.n878 0.120292
R6302 VDDD.n1029 VDDD.n880 0.120292
R6303 VDDD.n1025 VDDD.n880 0.120292
R6304 VDDD.n1025 VDDD.n1024 0.120292
R6305 VDDD.n1024 VDDD.n1023 0.120292
R6306 VDDD.n1023 VDDD.n884 0.120292
R6307 VDDD.n1018 VDDD.n884 0.120292
R6308 VDDD.n1018 VDDD.n1017 0.120292
R6309 VDDD.n1017 VDDD.n1016 0.120292
R6310 VDDD.n1016 VDDD.n887 0.120292
R6311 VDDD.n890 VDDD.n887 0.120292
R6312 VDDD.n1002 VDDD.n904 0.120292
R6313 VDDD.n995 VDDD.n904 0.120292
R6314 VDDD.n994 VDDD.n993 0.120292
R6315 VDDD.n987 VDDD.n912 0.120292
R6316 VDDD.n982 VDDD.n912 0.120292
R6317 VDDD.n980 VDDD.n918 0.120292
R6318 VDDD.n976 VDDD.n918 0.120292
R6319 VDDD.n976 VDDD.n975 0.120292
R6320 VDDD.n975 VDDD.n974 0.120292
R6321 VDDD.n974 VDDD.n921 0.120292
R6322 VDDD.n924 VDDD.n921 0.120292
R6323 VDDD.n969 VDDD.n924 0.120292
R6324 VDDD.n969 VDDD.n968 0.120292
R6325 VDDD.n968 VDDD.n927 0.120292
R6326 VDDD.n962 VDDD.n927 0.120292
R6327 VDDD.n962 VDDD.n961 0.120292
R6328 VDDD.n961 VDDD.n960 0.120292
R6329 VDDD.n960 VDDD.n930 0.120292
R6330 VDDD.n933 VDDD.n930 0.120292
R6331 VDDD.n934 VDDD.n933 0.120292
R6332 VDDD.n953 VDDD.n952 0.120292
R6333 VDDD.n952 VDDD.n936 0.120292
R6334 VDDD.n946 VDDD.n936 0.120292
R6335 VDDD.n1478 VDDD.n1448 0.120292
R6336 VDDD.n1471 VDDD.n1448 0.120292
R6337 VDDD.n1471 VDDD.n1470 0.120292
R6338 VDDD.n1467 VDDD.n1466 0.120292
R6339 VDDD.n1466 VDDD.n1465 0.120292
R6340 VDDD.n1465 VDDD.n1453 0.120292
R6341 VDDD.n1459 VDDD.n1453 0.120292
R6342 VDDD.n1503 VDDD.n1502 0.120292
R6343 VDDD.n1502 VDDD.n1501 0.120292
R6344 VDDD.n1501 VDDD.n1331 0.120292
R6345 VDDD.n1496 VDDD.n1331 0.120292
R6346 VDDD.n1496 VDDD.n1495 0.120292
R6347 VDDD.n1491 VDDD.n1336 0.120292
R6348 VDDD.n1486 VDDD.n1336 0.120292
R6349 VDDD.n1433 VDDD.n1432 0.120292
R6350 VDDD.n1419 VDDD.n1351 0.120292
R6351 VDDD.n1413 VDDD.n1365 0.120292
R6352 VDDD.n1407 VDDD.n1365 0.120292
R6353 VDDD.n1407 VDDD.n1406 0.120292
R6354 VDDD.n1406 VDDD.n1405 0.120292
R6355 VDDD.n1405 VDDD.n1369 0.120292
R6356 VDDD.n1401 VDDD.n1369 0.120292
R6357 VDDD.n1401 VDDD.n1400 0.120292
R6358 VDDD.n1400 VDDD.n1399 0.120292
R6359 VDDD.n1394 VDDD.n1381 0.120292
R6360 VDDD.n1394 VDDD.n1393 0.120292
R6361 VDDD.n1392 VDDD.n1383 0.120292
R6362 VDDD.n3004 VDDD.n3003 0.120292
R6363 VDDD.n3003 VDDD.n1114 0.120292
R6364 VDDD.n2997 VDDD.n1114 0.120292
R6365 VDDD.n2995 VDDD.n1121 0.120292
R6366 VDDD.n2991 VDDD.n1121 0.120292
R6367 VDDD.n2991 VDDD.n2990 0.120292
R6368 VDDD.n2990 VDDD.n1128 0.120292
R6369 VDDD.n2984 VDDD.n2983 0.120292
R6370 VDDD.n2983 VDDD.n1130 0.120292
R6371 VDDD.n2977 VDDD.n1130 0.120292
R6372 VDDD.n2976 VDDD.n1135 0.120292
R6373 VDDD.n1232 VDDD.n1148 0.120292
R6374 VDDD.n1227 VDDD.n1148 0.120292
R6375 VDDD.n1227 VDDD.n1226 0.120292
R6376 VDDD.n1226 VDDD.n1154 0.120292
R6377 VDDD.n1217 VDDD.n1216 0.120292
R6378 VDDD.n1216 VDDD.n1158 0.120292
R6379 VDDD.n1212 VDDD.n1158 0.120292
R6380 VDDD.n1212 VDDD.n1211 0.120292
R6381 VDDD.n1211 VDDD.n1160 0.120292
R6382 VDDD.n1207 VDDD.n1160 0.120292
R6383 VDDD.n1207 VDDD.n1206 0.120292
R6384 VDDD.n1206 VDDD.n1205 0.120292
R6385 VDDD.n1205 VDDD.n1162 0.120292
R6386 VDDD.n1201 VDDD.n1162 0.120292
R6387 VDDD.n1201 VDDD.n1200 0.120292
R6388 VDDD.n1197 VDDD.n1196 0.120292
R6389 VDDD.n1196 VDDD.n1165 0.120292
R6390 VDDD.n1192 VDDD.n1165 0.120292
R6391 VDDD.n1192 VDDD.n1191 0.120292
R6392 VDDD.n1191 VDDD.n1167 0.120292
R6393 VDDD.n1187 VDDD.n1167 0.120292
R6394 VDDD.n1187 VDDD.n1186 0.120292
R6395 VDDD.n1186 VDDD.n1185 0.120292
R6396 VDDD.n1185 VDDD.n1169 0.120292
R6397 VDDD.n1181 VDDD.n1169 0.120292
R6398 VDDD.n1181 VDDD.n1180 0.120292
R6399 VDDD.n2736 VDDD.n1306 0.120292
R6400 VDDD.n2731 VDDD.n1306 0.120292
R6401 VDDD.n2731 VDDD.n2730 0.120292
R6402 VDDD.n2730 VDDD.n1308 0.120292
R6403 VDDD.n1311 VDDD.n1308 0.120292
R6404 VDDD.n2724 VDDD.n1311 0.120292
R6405 VDDD.n2724 VDDD.n2723 0.120292
R6406 VDDD.n2723 VDDD.n2722 0.120292
R6407 VDDD.n2722 VDDD.n1313 0.120292
R6408 VDDD.n1557 VDDD.n1521 0.120292
R6409 VDDD.n1528 VDDD.n1521 0.120292
R6410 VDDD.n1529 VDDD.n1528 0.120292
R6411 VDDD.n1551 VDDD.n1529 0.120292
R6412 VDDD.n1551 VDDD.n1550 0.120292
R6413 VDDD.n1550 VDDD.n1549 0.120292
R6414 VDDD.n1545 VDDD.n1544 0.120292
R6415 VDDD.n1544 VDDD.n1534 0.120292
R6416 VDDD.n1540 VDDD.n1534 0.120292
R6417 VDDD.n1540 VDDD.n1539 0.120292
R6418 VDDD.n1539 VDDD.n1538 0.120292
R6419 VDDD.n1292 VDDD.n1291 0.120292
R6420 VDDD.n2747 VDDD.n1291 0.120292
R6421 VDDD.n2748 VDDD.n2747 0.120292
R6422 VDDD.n2761 VDDD.n1275 0.120292
R6423 VDDD.n2765 VDDD.n1275 0.120292
R6424 VDDD.n2766 VDDD.n2765 0.120292
R6425 VDDD.n2767 VDDD.n2766 0.120292
R6426 VDDD.n2767 VDDD.n1271 0.120292
R6427 VDDD.n2773 VDDD.n1271 0.120292
R6428 VDDD.n2774 VDDD.n2773 0.120292
R6429 VDDD.n2775 VDDD.n2774 0.120292
R6430 VDDD.n2775 VDDD.n1269 0.120292
R6431 VDDD.n1269 VDDD.n1268 0.120292
R6432 VDDD.n1268 VDDD.n1266 0.120292
R6433 VDDD.n2781 VDDD.n1266 0.120292
R6434 VDDD.n2782 VDDD.n2781 0.120292
R6435 VDDD.n2788 VDDD.n1260 0.120292
R6436 VDDD.n2789 VDDD.n2788 0.120292
R6437 VDDD.n2848 VDDD.n2800 0.120292
R6438 VDDD.n2843 VDDD.n2800 0.120292
R6439 VDDD.n2843 VDDD.n2842 0.120292
R6440 VDDD.n2842 VDDD.n2841 0.120292
R6441 VDDD.n2841 VDDD.n2802 0.120292
R6442 VDDD.n2837 VDDD.n2802 0.120292
R6443 VDDD.n2837 VDDD.n2836 0.120292
R6444 VDDD.n2836 VDDD.n2835 0.120292
R6445 VDDD.n2835 VDDD.n2806 0.120292
R6446 VDDD.n2829 VDDD.n2806 0.120292
R6447 VDDD.n2829 VDDD.n2828 0.120292
R6448 VDDD.n2828 VDDD.n2827 0.120292
R6449 VDDD.n2827 VDDD.n2811 0.120292
R6450 VDDD.n2823 VDDD.n2811 0.120292
R6451 VDDD.n2823 VDDD.n2822 0.120292
R6452 VDDD.n2821 VDDD.n2815 0.120292
R6453 VDDD.n2948 VDDD.n2947 0.120292
R6454 VDDD.n2947 VDDD.n1246 0.120292
R6455 VDDD.n2942 VDDD.n1246 0.120292
R6456 VDDD.n2936 VDDD.n2935 0.120292
R6457 VDDD.n2935 VDDD.n2864 0.120292
R6458 VDDD.n2865 VDDD.n2864 0.120292
R6459 VDDD.n2930 VDDD.n2865 0.120292
R6460 VDDD.n2930 VDDD.n2929 0.120292
R6461 VDDD.n2929 VDDD.n2928 0.120292
R6462 VDDD.n2928 VDDD.n2867 0.120292
R6463 VDDD.n2922 VDDD.n2867 0.120292
R6464 VDDD.n2922 VDDD.n2921 0.120292
R6465 VDDD.n2921 VDDD.n2920 0.120292
R6466 VDDD.n2920 VDDD.n2872 0.120292
R6467 VDDD.n2874 VDDD.n2872 0.120292
R6468 VDDD.n2915 VDDD.n2874 0.120292
R6469 VDDD.n2915 VDDD.n2914 0.120292
R6470 VDDD.n2914 VDDD.n2876 0.120292
R6471 VDDD.n2908 VDDD.n2876 0.120292
R6472 VDDD.n2908 VDDD.n2907 0.120292
R6473 VDDD.n2903 VDDD.n2902 0.120292
R6474 VDDD.n2899 VDDD.n2898 0.120292
R6475 VDDD.n2898 VDDD.n2897 0.120292
R6476 VDDD.n2897 VDDD.n2883 0.120292
R6477 VDDD.n1788 VDDD.n1787 0.120292
R6478 VDDD.n1783 VDDD.n1782 0.120292
R6479 VDDD.n1782 VDDD.n1705 0.120292
R6480 VDDD.n1777 VDDD.n1705 0.120292
R6481 VDDD.n1777 VDDD.n1776 0.120292
R6482 VDDD.n1776 VDDD.n1708 0.120292
R6483 VDDD.n1772 VDDD.n1708 0.120292
R6484 VDDD.n1763 VDDD.n1717 0.120292
R6485 VDDD.n1758 VDDD.n1757 0.120292
R6486 VDDD.n1757 VDDD.n1729 0.120292
R6487 VDDD.n1752 VDDD.n1729 0.120292
R6488 VDDD.n1752 VDDD.n1751 0.120292
R6489 VDDD.n1751 VDDD.n1731 0.120292
R6490 VDDD.n1746 VDDD.n1731 0.120292
R6491 VDDD.n1745 VDDD.n1744 0.120292
R6492 VDDD.n1744 VDDD.n1734 0.120292
R6493 VDDD.n1739 VDDD.n1734 0.120292
R6494 VDDD.n1739 VDDD.n1738 0.120292
R6495 VDDD.n1799 VDDD.n1798 0.120292
R6496 VDDD.n1804 VDDD.n1803 0.120292
R6497 VDDD.n1866 VDDD.n1810 0.120292
R6498 VDDD.n1860 VDDD.n1810 0.120292
R6499 VDDD.n1860 VDDD.n1859 0.120292
R6500 VDDD.n1859 VDDD.n1858 0.120292
R6501 VDDD.n1858 VDDD.n1815 0.120292
R6502 VDDD.n1852 VDDD.n1815 0.120292
R6503 VDDD.n1852 VDDD.n1851 0.120292
R6504 VDDD.n1846 VDDD.n1845 0.120292
R6505 VDDD.n1845 VDDD.n1820 0.120292
R6506 VDDD.n1841 VDDD.n1820 0.120292
R6507 VDDD.n1841 VDDD.n1840 0.120292
R6508 VDDD.n1840 VDDD.n1823 0.120292
R6509 VDDD.n1836 VDDD.n1823 0.120292
R6510 VDDD.n1836 VDDD.n1835 0.120292
R6511 VDDD.n1605 VDDD.n1604 0.120292
R6512 VDDD.n1612 VDDD.n1611 0.120292
R6513 VDDD.n1613 VDDD.n1612 0.120292
R6514 VDDD.n1613 VDDD.n1592 0.120292
R6515 VDDD.n1617 VDDD.n1592 0.120292
R6516 VDDD.n1618 VDDD.n1617 0.120292
R6517 VDDD.n1618 VDDD.n1589 0.120292
R6518 VDDD.n1622 VDDD.n1589 0.120292
R6519 VDDD.n1623 VDDD.n1622 0.120292
R6520 VDDD.n2593 VDDD.n2592 0.120292
R6521 VDDD.n2593 VDDD.n1574 0.120292
R6522 VDDD.n2601 VDDD.n1574 0.120292
R6523 VDDD.n2602 VDDD.n2601 0.120292
R6524 VDDD.n2674 VDDD.n2673 0.120292
R6525 VDDD.n2673 VDDD.n2607 0.120292
R6526 VDDD.n2608 VDDD.n2607 0.120292
R6527 VDDD.n2668 VDDD.n2608 0.120292
R6528 VDDD.n2668 VDDD.n2667 0.120292
R6529 VDDD.n2667 VDDD.n2666 0.120292
R6530 VDDD.n2666 VDDD.n2610 0.120292
R6531 VDDD.n2660 VDDD.n2610 0.120292
R6532 VDDD.n2660 VDDD.n2659 0.120292
R6533 VDDD.n2659 VDDD.n2658 0.120292
R6534 VDDD.n2658 VDDD.n2615 0.120292
R6535 VDDD.n2616 VDDD.n2615 0.120292
R6536 VDDD.n2653 VDDD.n2616 0.120292
R6537 VDDD.n2653 VDDD.n2652 0.120292
R6538 VDDD.n2652 VDDD.n2619 0.120292
R6539 VDDD.n2646 VDDD.n2619 0.120292
R6540 VDDD.n2646 VDDD.n2645 0.120292
R6541 VDDD.n2641 VDDD.n2640 0.120292
R6542 VDDD.n2637 VDDD.n2636 0.120292
R6543 VDDD.n2356 VDDD.n2355 0.120292
R6544 VDDD.n2355 VDDD.n2354 0.120292
R6545 VDDD.n2354 VDDD.n1901 0.120292
R6546 VDDD.n2347 VDDD.n1901 0.120292
R6547 VDDD.n2347 VDDD.n2346 0.120292
R6548 VDDD.n2346 VDDD.n2345 0.120292
R6549 VDDD.n2345 VDDD.n1905 0.120292
R6550 VDDD.n2341 VDDD.n1905 0.120292
R6551 VDDD.n2341 VDDD.n2340 0.120292
R6552 VDDD.n1955 VDDD.n1913 0.120292
R6553 VDDD.n1951 VDDD.n1913 0.120292
R6554 VDDD.n1951 VDDD.n1950 0.120292
R6555 VDDD.n1950 VDDD.n1949 0.120292
R6556 VDDD.n1949 VDDD.n1929 0.120292
R6557 VDDD.n1944 VDDD.n1929 0.120292
R6558 VDDD.n2366 VDDD.n2365 0.120292
R6559 VDDD.n2366 VDDD.n1884 0.120292
R6560 VDDD.n2372 VDDD.n1884 0.120292
R6561 VDDD.n1670 VDDD.n1669 0.120292
R6562 VDDD.n2394 VDDD.n1669 0.120292
R6563 VDDD.n2395 VDDD.n2394 0.120292
R6564 VDDD.n2396 VDDD.n2395 0.120292
R6565 VDDD.n2396 VDDD.n1666 0.120292
R6566 VDDD.n2401 VDDD.n1666 0.120292
R6567 VDDD.n2402 VDDD.n2401 0.120292
R6568 VDDD.n2403 VDDD.n2402 0.120292
R6569 VDDD.n2403 VDDD.n1664 0.120292
R6570 VDDD.n2410 VDDD.n1664 0.120292
R6571 VDDD.n2411 VDDD.n2410 0.120292
R6572 VDDD.n2416 VDDD.n2415 0.120292
R6573 VDDD.n2416 VDDD.n1654 0.120292
R6574 VDDD.n2480 VDDD.n2428 0.120292
R6575 VDDD.n2473 VDDD.n2428 0.120292
R6576 VDDD.n2473 VDDD.n2472 0.120292
R6577 VDDD.n2472 VDDD.n2431 0.120292
R6578 VDDD.n2467 VDDD.n2431 0.120292
R6579 VDDD.n2467 VDDD.n2466 0.120292
R6580 VDDD.n2466 VDDD.n2465 0.120292
R6581 VDDD.n2465 VDDD.n2434 0.120292
R6582 VDDD.n2459 VDDD.n2434 0.120292
R6583 VDDD.n2459 VDDD.n2458 0.120292
R6584 VDDD.n2458 VDDD.n2436 0.120292
R6585 VDDD.n2451 VDDD.n2436 0.120292
R6586 VDDD.n2449 VDDD.n2439 0.120292
R6587 VDDD.n2444 VDDD.n2439 0.120292
R6588 VDDD.n2444 VDDD.n2443 0.120292
R6589 VDDD.n2565 VDDD.n1643 0.120292
R6590 VDDD.n2560 VDDD.n1643 0.120292
R6591 VDDD.n2560 VDDD.n2559 0.120292
R6592 VDDD.n2554 VDDD.n2553 0.120292
R6593 VDDD.n2553 VDDD.n2495 0.120292
R6594 VDDD.n2549 VDDD.n2495 0.120292
R6595 VDDD.n2549 VDDD.n2548 0.120292
R6596 VDDD.n2548 VDDD.n2497 0.120292
R6597 VDDD.n2544 VDDD.n2497 0.120292
R6598 VDDD.n2544 VDDD.n2543 0.120292
R6599 VDDD.n2543 VDDD.n2542 0.120292
R6600 VDDD.n2542 VDDD.n2499 0.120292
R6601 VDDD.n2538 VDDD.n2499 0.120292
R6602 VDDD.n2538 VDDD.n2537 0.120292
R6603 VDDD.n2534 VDDD.n2533 0.120292
R6604 VDDD.n2533 VDDD.n2502 0.120292
R6605 VDDD.n2529 VDDD.n2502 0.120292
R6606 VDDD.n2529 VDDD.n2528 0.120292
R6607 VDDD.n2528 VDDD.n2504 0.120292
R6608 VDDD.n2524 VDDD.n2504 0.120292
R6609 VDDD.n2524 VDDD.n2523 0.120292
R6610 VDDD.n2523 VDDD.n2522 0.120292
R6611 VDDD.n2522 VDDD.n2506 0.120292
R6612 VDDD.n2518 VDDD.n2506 0.120292
R6613 VDDD.n2518 VDDD.n2517 0.120292
R6614 VDDD.n2017 VDDD.n1996 0.120292
R6615 VDDD.n2011 VDDD.n1996 0.120292
R6616 VDDD.n2011 VDDD.n2010 0.120292
R6617 VDDD.n2010 VDDD.n1999 0.120292
R6618 VDDD.n2005 VDDD.n1999 0.120292
R6619 VDDD.n2005 VDDD.n2004 0.120292
R6620 VDDD.n2321 VDDD.n2320 0.120292
R6621 VDDD.n2317 VDDD.n2316 0.120292
R6622 VDDD.n2316 VDDD.n1971 0.120292
R6623 VDDD.n2311 VDDD.n1971 0.120292
R6624 VDDD.n2311 VDDD.n2310 0.120292
R6625 VDDD.n2310 VDDD.n1973 0.120292
R6626 VDDD.n2304 VDDD.n2303 0.120292
R6627 VDDD.n2303 VDDD.n1976 0.120292
R6628 VDDD.n2298 VDDD.n1976 0.120292
R6629 VDDD.n2298 VDDD.n2297 0.120292
R6630 VDDD.n2082 VDDD.n2081 0.120292
R6631 VDDD.n2111 VDDD.n2110 0.120292
R6632 VDDD.n2112 VDDD.n2111 0.120292
R6633 VDDD.n2112 VDDD.n2066 0.120292
R6634 VDDD.n2116 VDDD.n2066 0.120292
R6635 VDDD.n2117 VDDD.n2116 0.120292
R6636 VDDD.n2117 VDDD.n2063 0.120292
R6637 VDDD.n2122 VDDD.n2063 0.120292
R6638 VDDD.n2123 VDDD.n2122 0.120292
R6639 VDDD.n2127 VDDD.n2126 0.120292
R6640 VDDD.n2127 VDDD.n2059 0.120292
R6641 VDDD.n2133 VDDD.n2059 0.120292
R6642 VDDD.n2134 VDDD.n2133 0.120292
R6643 VDDD.n2134 VDDD.n2057 0.120292
R6644 VDDD.n2139 VDDD.n2057 0.120292
R6645 VDDD.n2140 VDDD.n2139 0.120292
R6646 VDDD.n2145 VDDD.n2144 0.120292
R6647 VDDD.n2167 VDDD.n2166 0.120292
R6648 VDDD.n2167 VDDD.n2040 0.120292
R6649 VDDD.n2172 VDDD.n2040 0.120292
R6650 VDDD.n2173 VDDD.n2172 0.120292
R6651 VDDD.n2174 VDDD.n2173 0.120292
R6652 VDDD.n2174 VDDD.n2037 0.120292
R6653 VDDD.n2179 VDDD.n2037 0.120292
R6654 VDDD.n2180 VDDD.n2179 0.120292
R6655 VDDD.n2180 VDDD.n2035 0.120292
R6656 VDDD.n2184 VDDD.n2035 0.120292
R6657 VDDD.n2185 VDDD.n2184 0.120292
R6658 VDDD.n2193 VDDD.n2033 0.120292
R6659 VDDD.n2194 VDDD.n2193 0.120292
R6660 VDDD.n2195 VDDD.n2194 0.120292
R6661 VDDD.n2221 VDDD.n2220 0.120292
R6662 VDDD.n2222 VDDD.n2221 0.120292
R6663 VDDD.n2222 VDDD.n2025 0.120292
R6664 VDDD.n2227 VDDD.n2025 0.120292
R6665 VDDD.n2289 VDDD.n2288 0.120292
R6666 VDDD.n2288 VDDD.n2230 0.120292
R6667 VDDD.n2284 VDDD.n2230 0.120292
R6668 VDDD.n2284 VDDD.n2283 0.120292
R6669 VDDD.n2283 VDDD.n2232 0.120292
R6670 VDDD.n2279 VDDD.n2232 0.120292
R6671 VDDD.n2279 VDDD.n2278 0.120292
R6672 VDDD.n2278 VDDD.n2277 0.120292
R6673 VDDD.n2277 VDDD.n2234 0.120292
R6674 VDDD.n2273 VDDD.n2234 0.120292
R6675 VDDD.n2273 VDDD.n2272 0.120292
R6676 VDDD.n2269 VDDD.n2268 0.120292
R6677 VDDD.n2268 VDDD.n2237 0.120292
R6678 VDDD.n2264 VDDD.n2237 0.120292
R6679 VDDD.n2264 VDDD.n2263 0.120292
R6680 VDDD.n2263 VDDD.n2239 0.120292
R6681 VDDD.n2259 VDDD.n2239 0.120292
R6682 VDDD.n2259 VDDD.n2258 0.120292
R6683 VDDD.n2258 VDDD.n2257 0.120292
R6684 VDDD.n2257 VDDD.n2241 0.120292
R6685 VDDD.n2253 VDDD.n2241 0.120292
R6686 VDDD.n2253 VDDD.n2252 0.120292
R6687 VDDD.n136 VDDD.n135 0.120292
R6688 VDDD.n144 VDDD.n127 0.120292
R6689 VDDD.n145 VDDD.n144 0.120292
R6690 VDDD.n149 VDDD.n148 0.120292
R6691 VDDD.n149 VDDD.n124 0.120292
R6692 VDDD.n153 VDDD.n124 0.120292
R6693 VDDD.n154 VDDD.n153 0.120292
R6694 VDDD.n154 VDDD.n122 0.120292
R6695 VDDD.n158 VDDD.n122 0.120292
R6696 VDDD.n201 VDDD.n119 0.120292
R6697 VDDD.n196 VDDD.n195 0.120292
R6698 VDDD.n195 VDDD.n173 0.120292
R6699 VDDD.n191 VDDD.n173 0.120292
R6700 VDDD.n191 VDDD.n190 0.120292
R6701 VDDD.n190 VDDD.n175 0.120292
R6702 VDDD.n186 VDDD.n175 0.120292
R6703 VDDD.n186 VDDD.n185 0.120292
R6704 VDDD.n185 VDDD.n184 0.120292
R6705 VDDD.n184 VDDD.n177 0.120292
R6706 VDDD.n180 VDDD.n177 0.120292
R6707 VDDD.n180 VDDD.n179 0.120292
R6708 VDDD.n3704 VDDD.n3703 0.120292
R6709 VDDD.n3703 VDDD.n49 0.120292
R6710 VDDD.n109 VDDD.n59 0.120292
R6711 VDDD.n104 VDDD.n59 0.120292
R6712 VDDD.n104 VDDD.n103 0.120292
R6713 VDDD.n103 VDDD.n102 0.120292
R6714 VDDD.n102 VDDD.n69 0.120292
R6715 VDDD.n98 VDDD.n69 0.120292
R6716 VDDD.n98 VDDD.n97 0.120292
R6717 VDDD.n97 VDDD.n96 0.120292
R6718 VDDD.n93 VDDD.n92 0.120292
R6719 VDDD.n92 VDDD.n73 0.120292
R6720 VDDD.n88 VDDD.n73 0.120292
R6721 VDDD.n88 VDDD.n87 0.120292
R6722 VDDD.n87 VDDD.n75 0.120292
R6723 VDDD.n83 VDDD.n75 0.120292
R6724 VDDD.n83 VDDD.n82 0.120292
R6725 VDDD.n82 VDDD.n81 0.120292
R6726 VDDD.n81 VDDD.n77 0.120292
R6727 VDDD.n3727 VDDD.n37 0.120292
R6728 VDDD.n3733 VDDD.n37 0.120292
R6729 VDDD.n3734 VDDD.n3733 0.120292
R6730 VDDD.n3738 VDDD.n35 0.120292
R6731 VDDD.n3739 VDDD.n3738 0.120292
R6732 VDDD.n3740 VDDD.n3739 0.120292
R6733 VDDD.n3740 VDDD.n32 0.120292
R6734 VDDD.n3745 VDDD.n32 0.120292
R6735 VDDD.n3746 VDDD.n3745 0.120292
R6736 VDDD.n3747 VDDD.n3746 0.120292
R6737 VDDD.n3747 VDDD.n30 0.120292
R6738 VDDD.n3751 VDDD.n30 0.120292
R6739 VDDD.n3752 VDDD.n3751 0.120292
R6740 VDDD.n3753 VDDD.n3752 0.120292
R6741 VDDD.n3753 VDDD.n27 0.120292
R6742 VDDD.n3758 VDDD.n27 0.120292
R6743 VDDD.n3777 VDDD.n18 0.120292
R6744 VDDD.n3778 VDDD.n3777 0.120292
R6745 VDDD.n3779 VDDD.n3778 0.120292
R6746 VDDD.n3788 VDDD.n3787 0.120292
R6747 VDDD.n3788 VDDD.n13 0.120292
R6748 VDDD.n3792 VDDD.n13 0.120292
R6749 VDDD.n3793 VDDD.n3792 0.120292
R6750 VDDD.n3793 VDDD.n11 0.120292
R6751 VDDD.n3797 VDDD.n11 0.120292
R6752 VDDD.n3798 VDDD.n3797 0.120292
R6753 VDDD.n3799 VDDD.n3798 0.120292
R6754 VDDD.n3799 VDDD.n9 0.120292
R6755 VDDD.n3803 VDDD.n9 0.120292
R6756 VDDD.n3804 VDDD.n3803 0.120292
R6757 VDDD.n3808 VDDD.n3807 0.120292
R6758 VDDD.n3808 VDDD.n6 0.120292
R6759 VDDD.n3812 VDDD.n6 0.120292
R6760 VDDD.n3813 VDDD.n3812 0.120292
R6761 VDDD.n3813 VDDD.n4 0.120292
R6762 VDDD.n3817 VDDD.n4 0.120292
R6763 VDDD.n3818 VDDD.n3817 0.120292
R6764 VDDD.n3819 VDDD.n3818 0.120292
R6765 VDDD.n3819 VDDD.n2 0.120292
R6766 VDDD.n3824 VDDD.n2 0.120292
R6767 VDDD.n3825 VDDD.n3824 0.120292
R6768 VDDD.n3826 VDDD.n0 0.120292
R6769 VDDD.n3832 VDDD.n0 0.120292
R6770 VDDD.n3277 VDDD.n341 0.115235
R6771 VDDD.n3471 VDDD.n362 0.115235
R6772 VDDD.n3282 VDDD.n3281 0.115235
R6773 VDDD.n562 VDDD.n207 0.115235
R6774 VDDD.n3562 VDDD.n3473 0.107271
R6775 VDDD.n527 VDDD.n364 0.107271
R6776 VDDD.n3151 VDDD.n628 0.107271
R6777 VDDD.n865 VDDD.n855 0.107271
R6778 VDDD.n1383 VDDD.n1097 0.107271
R6779 VDDD.n2422 VDDD.n1654 0.107271
R6780 VDDD.n2145 VDDD.n2047 0.107271
R6781 VDDD.n77 VDDD.n43 0.107271
R6782 VDDD.n262 VDDD 0.105238
R6783 VDDD.n405 VDDD 0.105238
R6784 VDDD.n677 VDDD 0.105238
R6785 VDDD.n782 VDDD 0.105238
R6786 VDDD.n1446 VDDD 0.105238
R6787 VDDD.n1304 VDDD 0.105238
R6788 VDDD.n1698 VDDD 0.105238
R6789 VDDD.n1897 VDDD 0.105238
R6790 VDDD.n1994 VDDD 0.105238
R6791 VDDD.n247 VDDD.n246 0.102087
R6792 VDDD.n555 VDDD.n554 0.102087
R6793 VDDD.n3401 VDDD.n3400 0.102087
R6794 VDDD.n415 VDDD.n414 0.102087
R6795 VDDD.n616 VDDD.n615 0.102087
R6796 VDDD.n1040 VDDD.n1039 0.102087
R6797 VDDD.n1034 VDDD.n877 0.102087
R6798 VDDD.n986 VDDD.n916 0.102087
R6799 VDDD.n1489 VDDD.n1488 0.102087
R6800 VDDD.n2793 VDDD.n2792 0.102087
R6801 VDDD.n1603 VDDD.n1601 0.102087
R6802 VDDD.n3167 VDDD.n576 0.099575
R6803 VDDD VDDD.n3659 0.0981562
R6804 VDDD VDDD.n358 0.0981562
R6805 VDDD VDDD.n333 0.0981562
R6806 VDDD VDDD.n377 0.0981562
R6807 VDDD VDDD.n532 0.0981562
R6808 VDDD VDDD.n3431 0.0981562
R6809 VDDD VDDD.n3393 0.0981562
R6810 VDDD.n3108 VDDD 0.0981562
R6811 VDDD.n614 VDDD 0.0981562
R6812 VDDD VDDD.n607 0.0981562
R6813 VDDD.n3233 VDDD 0.0981562
R6814 VDDD.n3217 VDDD 0.0981562
R6815 VDDD.n766 VDDD 0.0981562
R6816 VDDD VDDD.n3032 0.0981562
R6817 VDDD VDDD.n1035 0.0981562
R6818 VDDD VDDD.n1029 0.0981562
R6819 VDDD VDDD.n987 0.0981562
R6820 VDDD VDDD.n980 0.0981562
R6821 VDDD VDDD.n1413 0.0981562
R6822 VDDD VDDD.n2995 0.0981562
R6823 VDDD.n1197 VDDD 0.0981562
R6824 VDDD VDDD.n2848 0.0981562
R6825 VDDD VDDD.n2936 0.0981562
R6826 VDDD.n1758 VDDD 0.0981562
R6827 VDDD.n1797 VDDD 0.0981562
R6828 VDDD.n1604 VDDD 0.0981562
R6829 VDDD.n1611 VDDD 0.0981562
R6830 VDDD.n2603 VDDD 0.0981562
R6831 VDDD VDDD.n2674 0.0981562
R6832 VDDD.n2415 VDDD 0.0981562
R6833 VDDD.n1646 VDDD 0.0981562
R6834 VDDD.n2534 VDDD 0.0981562
R6835 VDDD.n2317 VDDD 0.0981562
R6836 VDDD.n1979 VDDD 0.0981562
R6837 VDDD.n2126 VDDD 0.0981562
R6838 VDDD VDDD.n2033 0.0981562
R6839 VDDD.n2228 VDDD 0.0981562
R6840 VDDD.n2269 VDDD 0.0981562
R6841 VDDD.n135 VDDD 0.0981562
R6842 VDDD.n196 VDDD 0.0981562
R6843 VDDD.n3705 VDDD 0.0981562
R6844 VDDD.n93 VDDD 0.0981562
R6845 VDDD.n3807 VDDD 0.0981562
R6846 VDDD.n3826 VDDD 0.0981562
R6847 VDDD.n3673 VDDD.n214 0.0968542
R6848 VDDD.n446 VDDD.n379 0.0968542
R6849 VDDD.n745 VDDD.n744 0.0968542
R6850 VDDD.n3126 VDDD 0.0968542
R6851 VDDD.n3060 VDDD.n756 0.0968542
R6852 VDDD.n3042 VDDD 0.0968542
R6853 VDDD.n1503 VDDD.n1328 0.0968542
R6854 VDDD.n1558 VDDD.n1557 0.0968542
R6855 VDDD.n1764 VDDD.n1763 0.0968542
R6856 VDDD.n1956 VDDD.n1955 0.0968542
R6857 VDDD.n2321 VDDD.n1966 0.0968542
R6858 VDDD.n202 VDDD.n201 0.0968542
R6859 VDDD.n3696 VDDD.n54 0.0950946
R6860 VDDD.n111 VDDD.n57 0.0950946
R6861 VDDD.n3724 VDDD.n39 0.0950946
R6862 VDDD.n3762 VDDD.n3761 0.0950946
R6863 VDDD.n3766 VDDD.n24 0.0950946
R6864 VDDD.n3572 VDDD.n3571 0.0950946
R6865 VDDD.n3576 VDDD.n359 0.0950946
R6866 VDDD.n3518 VDDD.n3517 0.0950946
R6867 VDDD.n3524 VDDD.n3523 0.0950946
R6868 VDDD.n3686 VDDD.n3685 0.0950946
R6869 VDDD.n3679 VDDD.n213 0.0950946
R6870 VDDD.n3622 VDDD.n3621 0.0950946
R6871 VDDD.n3627 VDDD.n3626 0.0950946
R6872 VDDD.n3469 VDDD.n3468 0.0950946
R6873 VDDD.n3459 VDDD.n3458 0.0950946
R6874 VDDD.n3284 VDDD.n484 0.0950946
R6875 VDDD.n559 VDDD.n487 0.0950946
R6876 VDDD.n437 VDDD.n436 0.0950946
R6877 VDDD.n445 VDDD.n383 0.0950946
R6878 VDDD.n3318 VDDD.n3317 0.0950946
R6879 VDDD.n3411 VDDD.n3315 0.0950946
R6880 VDDD.n3162 VDDD.n3161 0.0950946
R6881 VDDD.n3166 VDDD.n624 0.0950946
R6882 VDDD.n3114 VDDD.n3113 0.0950946
R6883 VDDD.n3120 VDDD.n3119 0.0950946
R6884 VDDD.n3077 VDDD.n691 0.0950946
R6885 VDDD.n746 VDDD.n694 0.0950946
R6886 VDDD.n3274 VDDD.n3273 0.0950946
R6887 VDDD.n3264 VDDD.n3263 0.0950946
R6888 VDDD.n867 VDDD.n866 0.0950946
R6889 VDDD.n1047 VDDD.n864 0.0950946
R6890 VDDD.n3024 VDDD.n822 0.0950946
R6891 VDDD.n1090 VDDD.n825 0.0950946
R6892 VDDD.n3072 VDDD.n3071 0.0950946
R6893 VDDD.n3065 VDDD.n755 0.0950946
R6894 VDDD.n900 VDDD.n899 0.0950946
R6895 VDDD.n1004 VDDD.n897 0.0950946
R6896 VDDD.n3015 VDDD.n3014 0.0950946
R6897 VDDD.n1109 VDDD.n1108 0.0950946
R6898 VDDD.n1426 VDDD.n1347 0.0950946
R6899 VDDD.n1421 VDDD.n1350 0.0950946
R6900 VDDD.n1515 VDDD.n1514 0.0950946
R6901 VDDD.n1508 VDDD.n1327 0.0950946
R6902 VDDD.n2969 VDDD.n1139 0.0950946
R6903 VDDD.n1234 VDDD.n1144 0.0950946
R6904 VDDD.n2797 VDDD.n2796 0.0950946
R6905 VDDD.n2851 VDDD.n1257 0.0950946
R6906 VDDD.n2755 VDDD.n2754 0.0950946
R6907 VDDD.n2759 VDDD.n1279 0.0950946
R6908 VDDD.n2716 VDDD.n1318 0.0950946
R6909 VDDD.n1559 VDDD.n1519 0.0950946
R6910 VDDD.n2962 VDDD.n2961 0.0950946
R6911 VDDD.n2953 VDDD.n2952 0.0950946
R6912 VDDD.n2580 VDDD.n2579 0.0950946
R6913 VDDD.n2571 VDDD.n2570 0.0950946
R6914 VDDD.n2207 VDDD.n2206 0.0950946
R6915 VDDD.n2213 VDDD.n2212 0.0950946
R6916 VDDD.n1630 VDDD.n1629 0.0950946
R6917 VDDD.n2586 VDDD.n2585 0.0950946
R6918 VDDD.n1880 VDDD.n1879 0.0950946
R6919 VDDD.n1872 VDDD.n1871 0.0950946
R6920 VDDD.n1770 VDDD.n1712 0.0950946
R6921 VDDD.n1765 VDDD.n1715 0.0950946
R6922 VDDD.n2705 VDDD.n2704 0.0950946
R6923 VDDD.n2689 VDDD.n2688 0.0950946
R6924 VDDD.n2153 VDDD.n2152 0.0950946
R6925 VDDD.n2157 VDDD.n2044 0.0950946
R6926 VDDD.n2424 VDDD.n2423 0.0950946
R6927 VDDD.n2483 VDDD.n1653 0.0950946
R6928 VDDD.n2338 VDDD.n1908 0.0950946
R6929 VDDD.n1957 VDDD.n1911 0.0950946
R6930 VDDD.n2375 VDDD.n2374 0.0950946
R6931 VDDD.n2380 VDDD.n1676 0.0950946
R6932 VDDD.n2095 VDDD.n2073 0.0950946
R6933 VDDD.n2103 VDDD.n2102 0.0950946
R6934 VDDD.n2333 VDDD.n2332 0.0950946
R6935 VDDD.n2326 VDDD.n1965 0.0950946
R6936 VDDD.n162 VDDD.n161 0.0950946
R6937 VDDD.n203 VDDD.n117 0.0950946
R6938 VDDD VDDD.n576 0.0930646
R6939 VDDD VDDD.n781 0.0930646
R6940 VDDD VDDD.n3719 0.0917162
R6941 VDDD.n1142 VDDD.n564 0.0909059
R6942 VDDD.n3018 VDDD.n626 0.0909059
R6943 VDDD.n3022 VDDD.n3021 0.0909059
R6944 VDDD.n3074 VDDD.n749 0.0909059
R6945 VDDD.n2795 VDDD 0.0851354
R6946 VDDD.n2583 VDDD.n1237 0.0848235
R6947 VDDD.n2708 VDDD.n2707 0.0848235
R6948 VDDD.n1882 VDDD.n1281 0.0848235
R6949 VDDD.n2711 VDDD.n1561 0.0848235
R6950 VDDD.n3684 VDDD.n3683 0.0838333
R6951 VDDD.n3516 VDDD.n3514 0.0838333
R6952 VDDD.n3525 VDDD.n3496 0.0838333
R6953 VDDD.n440 VDDD.n438 0.0838333
R6954 VDDD.n3285 VDDD.n483 0.0838333
R6955 VDDD.n558 VDDD.n494 0.0838333
R6956 VDDD.n702 VDDD.n698 0.0838333
R6957 VDDD.n3112 VDDD.n663 0.0838333
R6958 VDDD.n3121 VDDD.n655 0.0838333
R6959 VDDD.n3070 VDDD.n3069 0.0838333
R6960 VDDD.n3025 VDDD.n821 0.0838333
R6961 VDDD.n1009 VDDD.n895 0.0838333
R6962 VDDD.n1513 VDDD.n1512 0.0838333
R6963 VDDD.n1146 VDDD.n1145 0.0838333
R6964 VDDD.n2717 VDDD.n1317 0.0838333
R6965 VDDD.n2753 VDDD.n1283 0.0838333
R6966 VDDD.n2760 VDDD.n1278 0.0838333
R6967 VDDD.n1722 VDDD.n1720 0.0838333
R6968 VDDD.n1878 VDDD.n1680 0.0838333
R6969 VDDD.n1873 VDDD.n1867 0.0838333
R6970 VDDD.n2690 VDDD.n2684 0.0838333
R6971 VDDD.n2587 VDDD.n1579 0.0838333
R6972 VDDD.n1922 VDDD.n1918 0.0838333
R6973 VDDD.n2373 VDDD.n1674 0.0838333
R6974 VDDD.n2379 VDDD.n2378 0.0838333
R6975 VDDD.n1642 VDDD.n1638 0.0838333
R6976 VDDD.n2331 VDDD.n2330 0.0838333
R6977 VDDD.n2094 VDDD.n2092 0.0838333
R6978 VDDD.n2104 VDDD.n2068 0.0838333
R6979 VDDD.n167 VDDD.n121 0.0838333
R6980 VDDD.n3697 VDDD.n53 0.0838333
R6981 VDDD.n110 VDDD.n58 0.0838333
R6982 VDDD.n3713 VDDD.n3712 0.0838333
R6983 VDDD.n3771 VDDD.n22 0.0838333
R6984 VDDD.n1941 VDDD 0.082648
R6985 VDDD.n2043 VDDD 0.082648
R6986 VDDD VDDD.n3295 0.082648
R6987 VDDD.n1659 VDDD 0.082648
R6988 VDDD.n1633 VDDD 0.0823353
R6989 VDDD.n2155 VDDD 0.0823353
R6990 VDDD.n1883 VDDD 0.0823353
R6991 VDDD.n2335 VDDD 0.0823353
R6992 VDDD.n3620 VDDD.n3619 0.0812292
R6993 VDDD.n3272 VDDD.n3271 0.0812292
R6994 VDDD.n1010 VDDD.n894 0.0812292
R6995 VDDD.n2970 VDDD.n1138 0.0812292
R6996 VDDD.n2960 VDDD.n2959 0.0812292
R6997 VDDD.n1628 VDDD.n1627 0.0812292
R6998 VDDD.n2578 VDDD.n2577 0.0812292
R6999 VDDD.n2205 VDDD.n2204 0.0812292
R7000 VDDD.n3772 VDDD.n21 0.0812292
R7001 VDDD.n1354 VDDD 0.0799271
R7002 VDDD.n3610 VDDD.n343 0.0760208
R7003 VDDD.n3422 VDDD.n3310 0.0760208
R7004 VDDD.n898 VDDD.n890 0.0760208
R7005 VDDD.n1137 VDDD.n1135 0.0760208
R7006 VDDD.n1623 VDDD.n1584 0.0760208
R7007 VDDD.n2443 VDDD.n1635 0.0760208
R7008 VDDD.n2195 VDDD.n2031 0.0760208
R7009 VDDD.n3760 VDDD.n3758 0.0760208
R7010 VDDD.n211 VDDD.n209 0.0708125
R7011 VDDD.n3633 VDDD.n337 0.0708125
R7012 VDDD.n434 VDDD.n386 0.0708125
R7013 VDDD.n3467 VDDD.n366 0.0708125
R7014 VDDD.n3410 VDDD.n3409 0.0708125
R7015 VDDD.n3078 VDDD.n690 0.0708125
R7016 VDDD.n3265 VDDD.n3259 0.0708125
R7017 VDDD.n862 VDDD.n860 0.0708125
R7018 VDDD.n1003 VDDD.n1002 0.0708125
R7019 VDDD.n1325 VDDD.n1323 0.0708125
R7020 VDDD.n3013 VDDD.n1099 0.0708125
R7021 VDDD.n1233 VDDD.n1232 0.0708125
R7022 VDDD.n2718 VDDD.n1316 0.0708125
R7023 VDDD.n2794 VDDD.n1254 0.0708125
R7024 VDDD.n1771 VDDD.n1711 0.0708125
R7025 VDDD.n2592 VDDD.n1577 0.0708125
R7026 VDDD.n2339 VDDD.n1907 0.0708125
R7027 VDDD.n2421 VDDD.n1650 0.0708125
R7028 VDDD.n1963 VDDD.n1961 0.0708125
R7029 VDDD.n2151 VDDD.n2049 0.0708125
R7030 VDDD.n2220 VDDD.n2027 0.0708125
R7031 VDDD.n160 VDDD.n159 0.0708125
R7032 VDDD.n3718 VDDD.n45 0.0708125
R7033 VDDD.n3765 VDDD.n18 0.0708125
R7034 VDDD.n64 VDDD.n62 0.0680676
R7035 VDDD.n64 VDDD.n63 0.0680676
R7036 VDDD.n3711 VDDD.n44 0.0680676
R7037 VDDD.n3711 VDDD.n3710 0.0680676
R7038 VDDD.n3770 VDDD.n23 0.0680676
R7039 VDDD.n3770 VDDD.n3769 0.0680676
R7040 VDDD.n3478 VDDD.n3474 0.0680676
R7041 VDDD.n3478 VDDD.n3477 0.0680676
R7042 VDDD.n3502 VDDD.n3501 0.0680676
R7043 VDDD.n3501 VDDD.n3500 0.0680676
R7044 VDDD.n3682 VDDD.n210 0.0680676
R7045 VDDD.n3682 VDDD.n3681 0.0680676
R7046 VDDD.n3617 VDDD.n344 0.0680676
R7047 VDDD.n3617 VDDD.n339 0.0680676
R7048 VDDD.n3455 VDDD.n365 0.0680676
R7049 VDDD.n3457 VDDD.n3455 0.0680676
R7050 VDDD.n491 VDDD.n489 0.0680676
R7051 VDDD.n491 VDDD.n490 0.0680676
R7052 VDDD.n441 VDDD.n385 0.0680676
R7053 VDDD.n442 VDDD.n441 0.0680676
R7054 VDDD.n3415 VDDD.n3314 0.0680676
R7055 VDDD.n3415 VDDD.n3414 0.0680676
R7056 VDDD.n631 VDDD.n629 0.0680676
R7057 VDDD.n631 VDDD.n630 0.0680676
R7058 VDDD.n662 VDDD.n661 0.0680676
R7059 VDDD.n661 VDDD.n660 0.0680676
R7060 VDDD.n701 VDDD.n699 0.0680676
R7061 VDDD.n701 VDDD.n700 0.0680676
R7062 VDDD.n3260 VDDD.n567 0.0680676
R7063 VDDD.n3262 VDDD.n3260 0.0680676
R7064 VDDD.n1051 VDDD.n863 0.0680676
R7065 VDDD.n1051 VDDD.n1050 0.0680676
R7066 VDDD.n833 VDDD.n831 0.0680676
R7067 VDDD.n833 VDDD.n832 0.0680676
R7068 VDDD.n3068 VDDD.n752 0.0680676
R7069 VDDD.n3068 VDDD.n3067 0.0680676
R7070 VDDD.n1008 VDDD.n896 0.0680676
R7071 VDDD.n1008 VDDD.n1007 0.0680676
R7072 VDDD.n1105 VDDD.n1098 0.0680676
R7073 VDDD.n1105 VDDD.n1104 0.0680676
R7074 VDDD.n1358 VDDD.n1348 0.0680676
R7075 VDDD.n1358 VDDD.n1349 0.0680676
R7076 VDDD.n1511 VDDD.n1324 0.0680676
R7077 VDDD.n1511 VDDD.n1510 0.0680676
R7078 VDDD.n2968 VDDD.n1140 0.0680676
R7079 VDDD.n1143 VDDD.n1140 0.0680676
R7080 VDDD.n2855 VDDD.n1255 0.0680676
R7081 VDDD.n2855 VDDD.n2854 0.0680676
R7082 VDDD.n1287 VDDD.n1284 0.0680676
R7083 VDDD.n1287 VDDD.n1286 0.0680676
R7084 VDDD.n2715 VDDD.n1319 0.0680676
R7085 VDDD.n1518 VDDD.n1319 0.0680676
R7086 VDDD.n2949 VDDD.n1240 0.0680676
R7087 VDDD.n2951 VDDD.n2949 0.0680676
R7088 VDDD.n2567 VDDD.n1636 0.0680676
R7089 VDDD.n2569 VDDD.n2567 0.0680676
R7090 VDDD.n2202 VDDD.n2030 0.0680676
R7091 VDDD.n2202 VDDD.n2029 0.0680676
R7092 VDDD.n1586 VDDD.n1585 0.0680676
R7093 VDDD.n1585 VDDD.n1580 0.0680676
R7094 VDDD.n1868 VDDD.n1681 0.0680676
R7095 VDDD.n1870 VDDD.n1868 0.0680676
R7096 VDDD.n1721 VDDD.n1713 0.0680676
R7097 VDDD.n1721 VDDD.n1714 0.0680676
R7098 VDDD.n2685 VDDD.n1567 0.0680676
R7099 VDDD.n2687 VDDD.n2685 0.0680676
R7100 VDDD.n2053 VDDD.n2048 0.0680676
R7101 VDDD.n2053 VDDD.n2052 0.0680676
R7102 VDDD.n2487 VDDD.n1651 0.0680676
R7103 VDDD.n2487 VDDD.n2486 0.0680676
R7104 VDDD.n1921 VDDD.n1919 0.0680676
R7105 VDDD.n1921 VDDD.n1920 0.0680676
R7106 VDDD.n2384 VDDD.n1675 0.0680676
R7107 VDDD.n2384 VDDD.n2383 0.0680676
R7108 VDDD.n2097 VDDD.n2096 0.0680676
R7109 VDDD.n2096 VDDD.n2071 0.0680676
R7110 VDDD.n2329 VDDD.n1962 0.0680676
R7111 VDDD.n2329 VDDD.n2328 0.0680676
R7112 VDDD.n166 VDDD.n164 0.0680676
R7113 VDDD.n166 VDDD.n165 0.0680676
R7114 VDDD.n2964 VDDD.n1237 0.0665765
R7115 VDDD.n2708 VDDD.n1095 0.0665765
R7116 VDDD.n2757 VDDD.n1281 0.0665765
R7117 VDDD.n2712 VDDD.n2711 0.0665765
R7118 VDDD.n492 VDDD.n488 0.0656042
R7119 VDDD.n3111 VDDD.n659 0.0656042
R7120 VDDD.n834 VDDD.n830 0.0656042
R7121 VDDD.n1359 VDDD.n1357 0.0656042
R7122 VDDD.n2752 VDDD.n1288 0.0656042
R7123 VDDD.n1877 VDDD.n1682 0.0656042
R7124 VDDD.n2386 VDDD.n2385 0.0656042
R7125 VDDD.n2093 VDDD.n2070 0.0656042
R7126 VDDD.n65 VDDD.n61 0.0656042
R7127 VDDD.n2965 VDDD.n1142 0.0604941
R7128 VDDD.n3018 VDDD.n3017 0.0604941
R7129 VDDD.n3021 VDDD.n1092 0.0604941
R7130 VDDD.n1517 VDDD.n749 0.0604941
R7131 VDDD VDDD.n232 0.0603958
R7132 VDDD VDDD.n231 0.0603958
R7133 VDDD VDDD.n230 0.0603958
R7134 VDDD VDDD.n251 0.0603958
R7135 VDDD VDDD.n243 0.0603958
R7136 VDDD.n3678 VDDD.n212 0.0603958
R7137 VDDD.n3678 VDDD.n3677 0.0603958
R7138 VDDD.n228 VDDD 0.0603958
R7139 VDDD.n3505 VDDD 0.0603958
R7140 VDDD VDDD.n3483 0.0603958
R7141 VDDD.n3600 VDDD 0.0603958
R7142 VDDD VDDD.n346 0.0603958
R7143 VDDD VDDD.n332 0.0603958
R7144 VDDD.n406 VDDD 0.0603958
R7145 VDDD.n407 VDDD 0.0603958
R7146 VDDD.n408 VDDD 0.0603958
R7147 VDDD VDDD.n392 0.0603958
R7148 VDDD.n419 VDDD 0.0603958
R7149 VDDD.n439 VDDD.n382 0.0603958
R7150 VDDD.n447 VDDD.n382 0.0603958
R7151 VDDD.n467 VDDD 0.0603958
R7152 VDDD.n468 VDDD 0.0603958
R7153 VDDD.n478 VDDD 0.0603958
R7154 VDDD VDDD.n3286 0.0603958
R7155 VDDD.n551 VDDD 0.0603958
R7156 VDDD.n547 VDDD 0.0603958
R7157 VDDD.n533 VDDD 0.0603958
R7158 VDDD VDDD.n519 0.0603958
R7159 VDDD.n528 VDDD 0.0603958
R7160 VDDD.n3444 VDDD 0.0603958
R7161 VDDD.n3432 VDDD 0.0603958
R7162 VDDD VDDD.n3306 0.0603958
R7163 VDDD.n3307 VDDD 0.0603958
R7164 VDDD.n3417 VDDD 0.0603958
R7165 VDDD VDDD.n3323 0.0603958
R7166 VDDD.n3404 VDDD 0.0603958
R7167 VDDD.n3328 VDDD 0.0603958
R7168 VDDD.n3394 VDDD 0.0603958
R7169 VDDD.n678 VDDD 0.0603958
R7170 VDDD.n3097 VDDD 0.0603958
R7171 VDDD VDDD.n3096 0.0603958
R7172 VDDD.n3093 VDDD 0.0603958
R7173 VDDD.n682 VDDD 0.0603958
R7174 VDDD.n3084 VDDD 0.0603958
R7175 VDDD.n704 VDDD.n703 0.0603958
R7176 VDDD.n703 VDDD.n695 0.0603958
R7177 VDDD VDDD.n731 0.0603958
R7178 VDDD.n3102 VDDD 0.0603958
R7179 VDDD.n3103 VDDD 0.0603958
R7180 VDDD.n3107 VDDD 0.0603958
R7181 VDDD.n643 VDDD 0.0603958
R7182 VDDD.n3148 VDDD 0.0603958
R7183 VDDD.n3150 VDDD 0.0603958
R7184 VDDD VDDD.n618 0.0603958
R7185 VDDD.n608 VDDD 0.0603958
R7186 VDDD.n594 VDDD 0.0603958
R7187 VDDD VDDD.n575 0.0603958
R7188 VDDD.n3247 VDDD 0.0603958
R7189 VDDD VDDD.n3246 0.0603958
R7190 VDDD VDDD.n3238 0.0603958
R7191 VDDD.n783 VDDD 0.0603958
R7192 VDDD.n808 VDDD 0.0603958
R7193 VDDD VDDD.n801 0.0603958
R7194 VDDD.n753 VDDD 0.0603958
R7195 VDDD.n3064 VDDD.n754 0.0603958
R7196 VDDD.n3064 VDDD.n3063 0.0603958
R7197 VDDD.n3034 VDDD 0.0603958
R7198 VDDD VDDD.n3033 0.0603958
R7199 VDDD.n1079 VDDD 0.0603958
R7200 VDDD.n1076 VDDD 0.0603958
R7201 VDDD.n1042 VDDD 0.0603958
R7202 VDDD.n1036 VDDD 0.0603958
R7203 VDDD.n1030 VDDD 0.0603958
R7204 VDDD.n995 VDDD 0.0603958
R7205 VDDD VDDD.n994 0.0603958
R7206 VDDD.n989 VDDD 0.0603958
R7207 VDDD VDDD.n988 0.0603958
R7208 VDDD VDDD.n981 0.0603958
R7209 VDDD VDDD.n934 0.0603958
R7210 VDDD.n953 VDDD 0.0603958
R7211 VDDD.n1447 VDDD 0.0603958
R7212 VDDD.n1480 VDDD 0.0603958
R7213 VDDD VDDD.n1479 0.0603958
R7214 VDDD VDDD.n1478 0.0603958
R7215 VDDD.n1467 VDDD 0.0603958
R7216 VDDD.n1507 VDDD.n1326 0.0603958
R7217 VDDD.n1507 VDDD.n1506 0.0603958
R7218 VDDD VDDD.n1485 0.0603958
R7219 VDDD.n1341 VDDD 0.0603958
R7220 VDDD.n1434 VDDD 0.0603958
R7221 VDDD VDDD.n1433 0.0603958
R7222 VDDD.n1428 VDDD 0.0603958
R7223 VDDD.n1414 VDDD 0.0603958
R7224 VDDD.n1393 VDDD 0.0603958
R7225 VDDD VDDD.n1392 0.0603958
R7226 VDDD.n3005 VDDD 0.0603958
R7227 VDDD VDDD.n3004 0.0603958
R7228 VDDD VDDD.n2996 0.0603958
R7229 VDDD VDDD.n1128 0.0603958
R7230 VDDD.n2985 VDDD 0.0603958
R7231 VDDD VDDD.n2984 0.0603958
R7232 VDDD VDDD.n2976 0.0603958
R7233 VDDD VDDD.n1154 0.0603958
R7234 VDDD.n1221 VDDD 0.0603958
R7235 VDDD VDDD.n1220 0.0603958
R7236 VDDD.n1217 VDDD 0.0603958
R7237 VDDD.n1305 VDDD 0.0603958
R7238 VDDD.n2737 VDDD 0.0603958
R7239 VDDD VDDD.n2736 0.0603958
R7240 VDDD.n1523 VDDD.n1522 0.0603958
R7241 VDDD.n1522 VDDD.n1520 0.0603958
R7242 VDDD.n1546 VDDD 0.0603958
R7243 VDDD VDDD.n1545 0.0603958
R7244 VDDD VDDD.n1294 0.0603958
R7245 VDDD VDDD.n1292 0.0603958
R7246 VDDD.n2783 VDDD 0.0603958
R7247 VDDD VDDD.n1260 0.0603958
R7248 VDDD.n2790 VDDD 0.0603958
R7249 VDDD.n2822 VDDD 0.0603958
R7250 VDDD VDDD.n2821 0.0603958
R7251 VDDD VDDD.n2948 0.0603958
R7252 VDDD VDDD.n2941 0.0603958
R7253 VDDD.n1250 VDDD 0.0603958
R7254 VDDD.n2937 VDDD 0.0603958
R7255 VDDD.n2907 VDDD 0.0603958
R7256 VDDD.n2903 VDDD 0.0603958
R7257 VDDD.n2902 VDDD 0.0603958
R7258 VDDD.n2899 VDDD 0.0603958
R7259 VDDD.n1699 VDDD 0.0603958
R7260 VDDD.n1700 VDDD 0.0603958
R7261 VDDD.n1789 VDDD 0.0603958
R7262 VDDD VDDD.n1788 0.0603958
R7263 VDDD.n1783 VDDD 0.0603958
R7264 VDDD.n1724 VDDD.n1723 0.0603958
R7265 VDDD.n1723 VDDD.n1716 0.0603958
R7266 VDDD VDDD.n1745 0.0603958
R7267 VDDD.n1798 VDDD 0.0603958
R7268 VDDD.n1803 VDDD 0.0603958
R7269 VDDD.n1847 VDDD 0.0603958
R7270 VDDD VDDD.n1846 0.0603958
R7271 VDDD.n1599 VDDD 0.0603958
R7272 VDDD.n1606 VDDD 0.0603958
R7273 VDDD VDDD.n2602 0.0603958
R7274 VDDD.n2680 VDDD 0.0603958
R7275 VDDD VDDD.n2679 0.0603958
R7276 VDDD VDDD.n2603 0.0603958
R7277 VDDD.n2675 VDDD 0.0603958
R7278 VDDD.n2645 VDDD 0.0603958
R7279 VDDD.n2641 VDDD 0.0603958
R7280 VDDD.n2640 VDDD 0.0603958
R7281 VDDD.n2637 VDDD 0.0603958
R7282 VDDD.n1898 VDDD 0.0603958
R7283 VDDD.n1899 VDDD 0.0603958
R7284 VDDD.n2356 VDDD 0.0603958
R7285 VDDD.n1924 VDDD.n1923 0.0603958
R7286 VDDD.n1923 VDDD.n1912 0.0603958
R7287 VDDD VDDD.n1943 0.0603958
R7288 VDDD VDDD.n1888 0.0603958
R7289 VDDD.n2365 VDDD 0.0603958
R7290 VDDD.n2412 VDDD 0.0603958
R7291 VDDD VDDD.n1658 0.0603958
R7292 VDDD VDDD.n2480 0.0603958
R7293 VDDD.n2451 VDDD 0.0603958
R7294 VDDD VDDD.n2450 0.0603958
R7295 VDDD VDDD.n2449 0.0603958
R7296 VDDD VDDD.n2566 0.0603958
R7297 VDDD VDDD.n2565 0.0603958
R7298 VDDD VDDD.n1645 0.0603958
R7299 VDDD.n2554 VDDD 0.0603958
R7300 VDDD.n1995 VDDD 0.0603958
R7301 VDDD.n2019 VDDD 0.0603958
R7302 VDDD VDDD.n2017 0.0603958
R7303 VDDD.n2325 VDDD.n1964 0.0603958
R7304 VDDD.n2325 VDDD.n2324 0.0603958
R7305 VDDD.n2305 VDDD 0.0603958
R7306 VDDD VDDD.n2304 0.0603958
R7307 VDDD.n2081 VDDD 0.0603958
R7308 VDDD.n2083 VDDD 0.0603958
R7309 VDDD.n2091 VDDD 0.0603958
R7310 VDDD.n2140 VDDD 0.0603958
R7311 VDDD.n2144 VDDD 0.0603958
R7312 VDDD.n2166 VDDD 0.0603958
R7313 VDDD VDDD.n2024 0.0603958
R7314 VDDD.n2289 VDDD 0.0603958
R7315 VDDD VDDD.n136 0.0603958
R7316 VDDD.n137 VDDD 0.0603958
R7317 VDDD VDDD.n128 0.0603958
R7318 VDDD VDDD.n127 0.0603958
R7319 VDDD.n148 VDDD 0.0603958
R7320 VDDD.n169 VDDD.n168 0.0603958
R7321 VDDD.n168 VDDD.n118 0.0603958
R7322 VDDD VDDD.n3704 0.0603958
R7323 VDDD.n3698 VDDD 0.0603958
R7324 VDDD.n3727 VDDD 0.0603958
R7325 VDDD VDDD.n35 0.0603958
R7326 VDDD.n3782 VDDD 0.0603958
R7327 VDDD.n3783 VDDD 0.0603958
R7328 VDDD.n3784 VDDD 0.0603958
R7329 VDDD.n3787 VDDD 0.0603958
R7330 VDDD VDDD.n3476 0.0577917
R7331 VDDD.n3618 VDDD 0.0577917
R7332 VDDD VDDD.n3294 0.0577917
R7333 VDDD VDDD.n623 0.0577917
R7334 VDDD.n870 VDDD 0.0577917
R7335 VDDD.n1107 VDDD 0.0577917
R7336 VDDD.n1256 VDDD 0.0577917
R7337 VDDD VDDD.n1242 0.0577917
R7338 VDDD.n1652 VDDD 0.0577917
R7339 VDDD VDDD.n2051 0.0577917
R7340 VDDD.n2203 VDDD 0.0577917
R7341 VDDD.n56 VDDD.n55 0.0574697
R7342 VDDD.n42 VDDD.n40 0.0574697
R7343 VDDD.n3768 VDDD.n25 0.0574697
R7344 VDDD.n3472 VDDD.n360 0.0574697
R7345 VDDD.n3521 VDDD.n3520 0.0574697
R7346 VDDD.n3680 VDDD.n208 0.0574697
R7347 VDDD.n342 VDDD.n340 0.0574697
R7348 VDDD.n3456 VDDD.n363 0.0574697
R7349 VDDD.n486 VDDD.n485 0.0574697
R7350 VDDD.n443 VDDD.n384 0.0574697
R7351 VDDD.n3413 VDDD.n3320 0.0574697
R7352 VDDD.n627 VDDD.n625 0.0574697
R7353 VDDD.n3117 VDDD.n3116 0.0574697
R7354 VDDD.n693 VDDD.n692 0.0574697
R7355 VDDD.n3261 VDDD.n565 0.0574697
R7356 VDDD.n1049 VDDD.n869 0.0574697
R7357 VDDD.n824 VDDD.n823 0.0574697
R7358 VDDD.n3066 VDDD.n750 0.0574697
R7359 VDDD.n1006 VDDD.n902 0.0574697
R7360 VDDD.n1103 VDDD.n1096 0.0574697
R7361 VDDD.n1424 VDDD.n1423 0.0574697
R7362 VDDD.n1509 VDDD.n1322 0.0574697
R7363 VDDD.n2967 VDDD.n1141 0.0574697
R7364 VDDD.n2853 VDDD.n2799 0.0574697
R7365 VDDD.n1282 VDDD.n1280 0.0574697
R7366 VDDD.n2714 VDDD.n1320 0.0574697
R7367 VDDD.n2950 VDDD.n1238 0.0574697
R7368 VDDD.n2568 VDDD.n1634 0.0574697
R7369 VDDD.n2210 VDDD.n2209 0.0574697
R7370 VDDD.n1631 VDDD.n1583 0.0574697
R7371 VDDD.n2584 VDDD.n1581 0.0574697
R7372 VDDD.n1869 VDDD.n1679 0.0574697
R7373 VDDD.n1768 VDDD.n1767 0.0574697
R7374 VDDD.n2686 VDDD.n1565 0.0574697
R7375 VDDD.n2046 VDDD.n2045 0.0574697
R7376 VDDD.n2426 VDDD.n2425 0.0574697
R7377 VDDD.n2485 VDDD.n2484 0.0574697
R7378 VDDD.n1910 VDDD.n1909 0.0574697
R7379 VDDD.n2382 VDDD.n1677 0.0574697
R7380 VDDD.n2098 VDDD.n2072 0.0574697
R7381 VDDD.n2101 VDDD.n2100 0.0574697
R7382 VDDD.n2327 VDDD.n1960 0.0574697
R7383 VDDD.n163 VDDD.n115 0.0574697
R7384 VDDD.n204 VDDD.n116 0.0574697
R7385 VDDD.n3526 VDDD.n3499 0.0551875
R7386 VDDD.n493 VDDD.n492 0.0551875
R7387 VDDD.n3122 VDDD.n659 0.0551875
R7388 VDDD.n836 VDDD.n834 0.0551875
R7389 VDDD.n1361 VDDD.n1359 0.0551875
R7390 VDDD.n1288 VDDD.n1285 0.0551875
R7391 VDDD.n1874 VDDD.n1682 0.0551875
R7392 VDDD.n2385 VDDD.n1671 0.0551875
R7393 VDDD.n2105 VDDD.n2070 0.0551875
R7394 VDDD.n66 VDDD.n65 0.0551875
R7395 VDDD.n1089 VDDD 0.0525833
R7396 VDDD.n1420 VDDD 0.0525833
R7397 VDDD.n3325 VDDD.n3324 0.0512937
R7398 VDDD.n3465 VDDD.n3464 0.0510929
R7399 VDDD.n243 VDDD.n209 0.0499792
R7400 VDDD.n3570 VDDD.n3569 0.0499792
R7401 VDDD.n3629 VDDD.n337 0.0499792
R7402 VDDD.n434 VDDD.n433 0.0499792
R7403 VDDD.n3467 VDDD.n3466 0.0499792
R7404 VDDD.n3410 VDDD.n3322 0.0499792
R7405 VDDD.n3079 VDDD.n3078 0.0499792
R7406 VDDD.n3160 VDDD.n3159 0.0499792
R7407 VDDD.n3266 VDDD.n3265 0.0499792
R7408 VDDD.n1053 VDDD.n862 0.0499792
R7409 VDDD.n1003 VDDD.n903 0.0499792
R7410 VDDD.n1459 VDDD.n1323 0.0499792
R7411 VDDD.n3013 VDDD.n3012 0.0499792
R7412 VDDD.n1233 VDDD.n1147 0.0499792
R7413 VDDD.n1316 VDDD.n1313 0.0499792
R7414 VDDD.n2857 VDDD.n1254 0.0499792
R7415 VDDD.n1772 VDDD.n1771 0.0499792
R7416 VDDD.n2703 VDDD.n2702 0.0499792
R7417 VDDD.n2588 VDDD.n1577 0.0499792
R7418 VDDD.n2340 VDDD.n2339 0.0499792
R7419 VDDD.n2489 VDDD.n1650 0.0499792
R7420 VDDD.n2004 VDDD.n1961 0.0499792
R7421 VDDD.n2151 VDDD.n2150 0.0499792
R7422 VDDD.n2215 VDDD.n2027 0.0499792
R7423 VDDD.n160 VDDD.n158 0.0499792
R7424 VDDD.n3718 VDDD.n3717 0.0499792
R7425 VDDD.n3765 VDDD.n19 0.0499792
R7426 VDDD.n3616 VDDD.n343 0.0447708
R7427 VDDD.n3312 VDDD.n3310 0.0447708
R7428 VDDD.n568 VDDD.n566 0.0447708
R7429 VDDD.n898 VDDD.n891 0.0447708
R7430 VDDD.n2971 VDDD.n1137 0.0447708
R7431 VDDD.n1241 VDDD.n1239 0.0447708
R7432 VDDD.n1626 VDDD.n1584 0.0447708
R7433 VDDD.n1637 VDDD.n1635 0.0447708
R7434 VDDD.n2201 VDDD.n2031 0.0447708
R7435 VDDD.n3760 VDDD.n3759 0.0447708
R7436 VDDD VDDD.n3499 0.0434688
R7437 VDDD.n62 VDDD.n54 0.0410405
R7438 VDDD.n63 VDDD.n57 0.0410405
R7439 VDDD.n3719 VDDD.n44 0.0410405
R7440 VDDD.n3710 VDDD.n39 0.0410405
R7441 VDDD.n3761 VDDD.n23 0.0410405
R7442 VDDD.n3769 VDDD.n24 0.0410405
R7443 VDDD.n3571 VDDD.n3474 0.0410405
R7444 VDDD.n3477 VDDD.n359 0.0410405
R7445 VDDD.n3517 VDDD.n3502 0.0410405
R7446 VDDD.n3524 VDDD.n3500 0.0410405
R7447 VDDD.n3685 VDDD.n210 0.0410405
R7448 VDDD.n3681 VDDD.n3679 0.0410405
R7449 VDDD.n3621 VDDD.n344 0.0410405
R7450 VDDD.n3627 VDDD.n339 0.0410405
R7451 VDDD.n3468 VDDD.n365 0.0410405
R7452 VDDD.n3458 VDDD.n3457 0.0410405
R7453 VDDD.n489 VDDD.n484 0.0410405
R7454 VDDD.n490 VDDD.n487 0.0410405
R7455 VDDD.n437 VDDD.n385 0.0410405
R7456 VDDD.n442 VDDD.n383 0.0410405
R7457 VDDD.n3317 VDDD.n3314 0.0410405
R7458 VDDD.n3414 VDDD.n3315 0.0410405
R7459 VDDD.n3161 VDDD.n629 0.0410405
R7460 VDDD.n630 VDDD.n624 0.0410405
R7461 VDDD.n3113 VDDD.n662 0.0410405
R7462 VDDD.n3120 VDDD.n660 0.0410405
R7463 VDDD.n699 VDDD.n691 0.0410405
R7464 VDDD.n700 VDDD.n694 0.0410405
R7465 VDDD.n3273 VDDD.n567 0.0410405
R7466 VDDD.n3263 VDDD.n3262 0.0410405
R7467 VDDD.n866 VDDD.n863 0.0410405
R7468 VDDD.n1050 VDDD.n864 0.0410405
R7469 VDDD.n831 VDDD.n822 0.0410405
R7470 VDDD.n832 VDDD.n825 0.0410405
R7471 VDDD.n3071 VDDD.n752 0.0410405
R7472 VDDD.n3067 VDDD.n3065 0.0410405
R7473 VDDD.n899 VDDD.n896 0.0410405
R7474 VDDD.n1007 VDDD.n897 0.0410405
R7475 VDDD.n3014 VDDD.n1098 0.0410405
R7476 VDDD.n1108 VDDD.n1104 0.0410405
R7477 VDDD.n1348 VDDD.n1347 0.0410405
R7478 VDDD.n1350 VDDD.n1349 0.0410405
R7479 VDDD.n1514 VDDD.n1324 0.0410405
R7480 VDDD.n1510 VDDD.n1508 0.0410405
R7481 VDDD.n2969 VDDD.n2968 0.0410405
R7482 VDDD.n1144 VDDD.n1143 0.0410405
R7483 VDDD.n2796 VDDD.n1255 0.0410405
R7484 VDDD.n2854 VDDD.n1257 0.0410405
R7485 VDDD.n2754 VDDD.n1284 0.0410405
R7486 VDDD.n1286 VDDD.n1279 0.0410405
R7487 VDDD.n2716 VDDD.n2715 0.0410405
R7488 VDDD.n1519 VDDD.n1518 0.0410405
R7489 VDDD.n2961 VDDD.n1240 0.0410405
R7490 VDDD.n2952 VDDD.n2951 0.0410405
R7491 VDDD.n2579 VDDD.n1636 0.0410405
R7492 VDDD.n2570 VDDD.n2569 0.0410405
R7493 VDDD.n2206 VDDD.n2030 0.0410405
R7494 VDDD.n2213 VDDD.n2029 0.0410405
R7495 VDDD.n1629 VDDD.n1586 0.0410405
R7496 VDDD.n2586 VDDD.n1580 0.0410405
R7497 VDDD.n1879 VDDD.n1681 0.0410405
R7498 VDDD.n1872 VDDD.n1870 0.0410405
R7499 VDDD.n1713 VDDD.n1712 0.0410405
R7500 VDDD.n1715 VDDD.n1714 0.0410405
R7501 VDDD.n2704 VDDD.n1567 0.0410405
R7502 VDDD.n2689 VDDD.n2687 0.0410405
R7503 VDDD.n2152 VDDD.n2048 0.0410405
R7504 VDDD.n2052 VDDD.n2044 0.0410405
R7505 VDDD.n2423 VDDD.n1651 0.0410405
R7506 VDDD.n2486 VDDD.n1653 0.0410405
R7507 VDDD.n1919 VDDD.n1908 0.0410405
R7508 VDDD.n1920 VDDD.n1911 0.0410405
R7509 VDDD.n2374 VDDD.n1675 0.0410405
R7510 VDDD.n2383 VDDD.n1676 0.0410405
R7511 VDDD.n2097 VDDD.n2095 0.0410405
R7512 VDDD.n2103 VDDD.n2071 0.0410405
R7513 VDDD.n2332 VDDD.n1962 0.0410405
R7514 VDDD.n2328 VDDD.n2326 0.0410405
R7515 VDDD.n164 VDDD.n162 0.0410405
R7516 VDDD.n165 VDDD.n117 0.0410405
R7517 VDDD.n3578 VDDD.n3577 0.0395625
R7518 VDDD.n3620 VDDD.n3616 0.0395625
R7519 VDDD.n3460 VDDD.n3453 0.0395625
R7520 VDDD.n3272 VDDD.n568 0.0395625
R7521 VDDD.n1046 VDDD.n1045 0.0395625
R7522 VDDD.n894 VDDD.n891 0.0395625
R7523 VDDD.n1111 VDDD.n1110 0.0395625
R7524 VDDD.n2971 VDDD.n2970 0.0395625
R7525 VDDD.n2850 VDDD.n2849 0.0395625
R7526 VDDD.n2960 VDDD.n1241 0.0395625
R7527 VDDD.n2693 VDDD.n1571 0.0395625
R7528 VDDD.n1628 VDDD.n1626 0.0395625
R7529 VDDD.n2482 VDDD.n2481 0.0395625
R7530 VDDD.n2578 VDDD.n1637 0.0395625
R7531 VDDD.n2159 VDDD.n2158 0.0395625
R7532 VDDD.n2205 VDDD.n2201 0.0395625
R7533 VDDD.n3726 VDDD.n3725 0.0395625
R7534 VDDD.n3759 VDDD.n21 0.0395625
R7535 VDDD.n3277 VDDD.n3276 0.0361647
R7536 VDDD.n3164 VDDD.n362 0.0361647
R7537 VDDD.n3281 VDDD.n561 0.0361647
R7538 VDDD.n3075 VDDD.n562 0.0361647
R7539 VDDD.n3629 VDDD.n3628 0.0343542
R7540 VDDD.n3322 VDDD.n3321 0.0343542
R7541 VDDD.n3266 VDDD.n572 0.0343542
R7542 VDDD.n903 VDDD.n895 0.0343542
R7543 VDDD.n1147 VDDD.n1146 0.0343542
R7544 VDDD.n2955 VDDD.n1245 0.0343542
R7545 VDDD.n2588 VDDD.n2587 0.0343542
R7546 VDDD.n2573 VDDD.n1642 0.0343542
R7547 VDDD.n2215 VDDD.n2214 0.0343542
R7548 VDDD.n22 VDDD.n19 0.0343542
R7549 VDDD.n3104 VDDD 0.0330521
R7550 VDDD.n993 VDDD 0.0330521
R7551 VDDD VDDD.n1351 0.0330521
R7552 VDDD.n2815 VDDD 0.0330521
R7553 VDDD.n1799 VDDD 0.0330521
R7554 VDDD.n232 VDDD 0.03175
R7555 VDDD.n231 VDDD 0.03175
R7556 VDDD VDDD.n230 0.03175
R7557 VDDD VDDD.n228 0.03175
R7558 VDDD.n3569 VDDD 0.03175
R7559 VDDD.n3475 VDDD 0.03175
R7560 VDDD.n3600 VDDD 0.03175
R7561 VDDD.n333 VDDD 0.03175
R7562 VDDD VDDD.n406 0.03175
R7563 VDDD VDDD.n407 0.03175
R7564 VDDD VDDD.n467 0.03175
R7565 VDDD VDDD.n478 0.03175
R7566 VDDD.n3461 VDDD 0.03175
R7567 VDDD VDDD.n3328 0.03175
R7568 VDDD VDDD.n678 0.03175
R7569 VDDD.n3097 VDDD 0.03175
R7570 VDDD.n3096 VDDD 0.03175
R7571 VDDD VDDD.n3102 0.03175
R7572 VDDD VDDD.n3148 0.03175
R7573 VDDD.n3168 VDDD 0.03175
R7574 VDDD.n3247 VDDD 0.03175
R7575 VDDD VDDD.n783 0.03175
R7576 VDDD.n808 VDDD 0.03175
R7577 VDDD.n3034 VDDD 0.03175
R7578 VDDD.n835 VDDD 0.03175
R7579 VDDD VDDD.n871 0.03175
R7580 VDDD.n1045 VDDD 0.03175
R7581 VDDD.n989 VDDD 0.03175
R7582 VDDD VDDD.n1447 0.03175
R7583 VDDD.n1480 VDDD 0.03175
R7584 VDDD.n1479 VDDD 0.03175
R7585 VDDD VDDD.n1341 0.03175
R7586 VDDD.n1434 VDDD 0.03175
R7587 VDDD.n1360 VDDD 0.03175
R7588 VDDD VDDD.n1102 0.03175
R7589 VDDD.n3005 VDDD 0.03175
R7590 VDDD.n2985 VDDD 0.03175
R7591 VDDD.n1221 VDDD 0.03175
R7592 VDDD VDDD.n1305 0.03175
R7593 VDDD.n2737 VDDD 0.03175
R7594 VDDD.n1294 VDDD 0.03175
R7595 VDDD VDDD.n1252 0.03175
R7596 VDDD.n2955 VDDD 0.03175
R7597 VDDD VDDD.n1250 0.03175
R7598 VDDD VDDD.n1699 0.03175
R7599 VDDD VDDD.n1700 0.03175
R7600 VDDD.n1789 VDDD 0.03175
R7601 VDDD VDDD.n1797 0.03175
R7602 VDDD.n1847 VDDD 0.03175
R7603 VDDD.n2691 VDDD 0.03175
R7604 VDDD VDDD.n2693 0.03175
R7605 VDDD.n2680 VDDD 0.03175
R7606 VDDD VDDD.n1898 0.03175
R7607 VDDD VDDD.n1899 0.03175
R7608 VDDD.n1888 VDDD 0.03175
R7609 VDDD.n2412 VDDD 0.03175
R7610 VDDD VDDD.n1648 0.03175
R7611 VDDD.n2481 VDDD 0.03175
R7612 VDDD.n2450 VDDD 0.03175
R7613 VDDD.n2566 VDDD 0.03175
R7614 VDDD.n1646 VDDD 0.03175
R7615 VDDD VDDD.n1995 0.03175
R7616 VDDD.n2019 VDDD 0.03175
R7617 VDDD.n2305 VDDD 0.03175
R7618 VDDD VDDD.n1979 0.03175
R7619 VDDD.n2050 VDDD 0.03175
R7620 VDDD.n2228 VDDD 0.03175
R7621 VDDD.n137 VDDD 0.03175
R7622 VDDD.n128 VDDD 0.03175
R7623 VDDD.n3705 VDDD 0.03175
R7624 VDDD.n3714 VDDD 0.03175
R7625 VDDD VDDD.n3726 0.03175
R7626 VDDD VDDD.n3782 0.03175
R7627 VDDD VDDD.n3783 0.03175
R7628 VDDD.n3784 VDDD 0.03175
R7629 VDDD VDDD.n569 0.0304479
R7630 VDDD.n2209 VDDD.n2208 0.0292489
R7631 VDDD.n2211 VDDD.n2210 0.0292489
R7632 VDDD.n2581 VDDD.n1634 0.0292489
R7633 VDDD.n2568 VDDD.n1632 0.0292489
R7634 VDDD.n2963 VDDD.n1238 0.0292489
R7635 VDDD.n2950 VDDD.n1236 0.0292489
R7636 VDDD.n2967 VDDD.n2966 0.0292489
R7637 VDDD.n1235 VDDD.n1141 0.0292489
R7638 VDDD.n902 VDDD.n901 0.0292489
R7639 VDDD.n1006 VDDD.n1005 0.0292489
R7640 VDDD.n3275 VDDD.n565 0.0292489
R7641 VDDD.n3261 VDDD.n563 0.0292489
R7642 VDDD.n3320 VDDD.n3319 0.0292489
R7643 VDDD.n3413 VDDD.n3412 0.0292489
R7644 VDDD.n3623 VDDD.n342 0.0292489
R7645 VDDD.n3625 VDDD.n340 0.0292489
R7646 VDDD.n3763 VDDD.n25 0.0292489
R7647 VDDD.n3768 VDDD.n3767 0.0292489
R7648 VDDD.n1582 VDDD.n1581 0.0292489
R7649 VDDD.n1583 VDDD.n1582 0.0292489
R7650 VDDD.n2154 VDDD.n2046 0.0292489
R7651 VDDD.n2156 VDDD.n2045 0.0292489
R7652 VDDD.n2706 VDDD.n1565 0.0292489
R7653 VDDD.n2686 VDDD.n1563 0.0292489
R7654 VDDD.n2799 VDDD.n2798 0.0292489
R7655 VDDD.n2853 VDDD.n2852 0.0292489
R7656 VDDD.n3016 VDDD.n1096 0.0292489
R7657 VDDD.n1103 VDDD.n1094 0.0292489
R7658 VDDD.n869 VDDD.n868 0.0292489
R7659 VDDD.n1049 VDDD.n1048 0.0292489
R7660 VDDD.n3163 VDDD.n627 0.0292489
R7661 VDDD.n3165 VDDD.n625 0.0292489
R7662 VDDD.n3470 VDDD.n363 0.0292489
R7663 VDDD.n3456 VDDD.n361 0.0292489
R7664 VDDD.n3573 VDDD.n3472 0.0292489
R7665 VDDD.n3575 VDDD.n360 0.0292489
R7666 VDDD.n3721 VDDD.n42 0.0292489
R7667 VDDD.n3723 VDDD.n40 0.0292489
R7668 VDDD.n2485 VDDD.n2427 0.0292489
R7669 VDDD.n2427 VDDD.n2426 0.0292489
R7670 VDDD.n2376 VDDD.n1677 0.0292489
R7671 VDDD.n2382 VDDD.n2381 0.0292489
R7672 VDDD.n1881 VDDD.n1679 0.0292489
R7673 VDDD.n1869 VDDD.n1678 0.0292489
R7674 VDDD.n2756 VDDD.n1282 0.0292489
R7675 VDDD.n2758 VDDD.n1280 0.0292489
R7676 VDDD.n1425 VDDD.n1424 0.0292489
R7677 VDDD.n1423 VDDD.n1422 0.0292489
R7678 VDDD.n3023 VDDD.n823 0.0292489
R7679 VDDD.n1091 VDDD.n824 0.0292489
R7680 VDDD.n3116 VDDD.n3115 0.0292489
R7681 VDDD.n3118 VDDD.n3117 0.0292489
R7682 VDDD.n3283 VDDD.n485 0.0292489
R7683 VDDD.n560 VDDD.n486 0.0292489
R7684 VDDD.n3520 VDDD.n3519 0.0292489
R7685 VDDD.n3522 VDDD.n3521 0.0292489
R7686 VDDD.n3695 VDDD.n55 0.0292489
R7687 VDDD.n112 VDDD.n56 0.0292489
R7688 VDDD.n2100 VDDD.n2099 0.0292489
R7689 VDDD.n2099 VDDD.n2098 0.0292489
R7690 VDDD.n2334 VDDD.n1960 0.0292489
R7691 VDDD.n2327 VDDD.n1959 0.0292489
R7692 VDDD.n2337 VDDD.n1909 0.0292489
R7693 VDDD.n1958 VDDD.n1910 0.0292489
R7694 VDDD.n1769 VDDD.n1768 0.0292489
R7695 VDDD.n1767 VDDD.n1766 0.0292489
R7696 VDDD.n2714 VDDD.n2713 0.0292489
R7697 VDDD.n1560 VDDD.n1320 0.0292489
R7698 VDDD.n1516 VDDD.n1322 0.0292489
R7699 VDDD.n1509 VDDD.n1321 0.0292489
R7700 VDDD.n3073 VDDD.n750 0.0292489
R7701 VDDD.n3066 VDDD.n748 0.0292489
R7702 VDDD.n3076 VDDD.n692 0.0292489
R7703 VDDD.n747 VDDD.n693 0.0292489
R7704 VDDD.n435 VDDD.n384 0.0292489
R7705 VDDD.n444 VDDD.n443 0.0292489
R7706 VDDD.n3687 VDDD.n208 0.0292489
R7707 VDDD.n3680 VDDD.n206 0.0292489
R7708 VDDD.n116 VDDD.n114 0.0292489
R7709 VDDD.n163 VDDD.n114 0.0292489
R7710 VDDD.n3526 VDDD.n3525 0.0291458
R7711 VDDD.n494 VDDD.n493 0.0291458
R7712 VDDD.n3416 VDDD 0.0291458
R7713 VDDD.n836 VDDD.n835 0.0291458
R7714 VDDD.n1285 VDDD.n1278 0.0291458
R7715 VDDD.n1874 VDDD.n1873 0.0291458
R7716 VDDD.n2378 VDDD.n1671 0.0291458
R7717 VDDD.n2105 VDDD.n2104 0.0291458
R7718 VDDD.n66 VDDD.n58 0.0291458
R7719 VDDD VDDD.n751 0.0278438
R7720 VDDD VDDD.n2572 0.0278438
R7721 VDDD.n3479 VDDD 0.0265417
R7722 VDDD.n3628 VDDD 0.0265417
R7723 VDDD.n3454 VDDD 0.0265417
R7724 VDDD.n3321 VDDD 0.0265417
R7725 VDDD.n632 VDDD 0.0265417
R7726 VDDD.n572 VDDD 0.0265417
R7727 VDDD.n1052 VDDD 0.0265417
R7728 VDDD VDDD.n1106 0.0265417
R7729 VDDD.n2856 VDDD 0.0265417
R7730 VDDD.n1245 VDDD 0.0265417
R7731 VDDD.n2488 VDDD 0.0265417
R7732 VDDD.n2054 VDDD 0.0265417
R7733 VDDD.n2214 VDDD 0.0265417
R7734 VDDD.n3683 VDDD.n212 0.0239375
R7735 VDDD.n3677 VDDD.n214 0.0239375
R7736 VDDD.n440 VDDD.n439 0.0239375
R7737 VDDD.n447 VDDD.n446 0.0239375
R7738 VDDD.n704 VDDD.n702 0.0239375
R7739 VDDD.n745 VDDD.n695 0.0239375
R7740 VDDD VDDD.n3125 0.0239375
R7741 VDDD.n3069 VDDD.n754 0.0239375
R7742 VDDD.n3063 VDDD.n756 0.0239375
R7743 VDDD VDDD.n766 0.0239375
R7744 VDDD.n1512 VDDD.n1326 0.0239375
R7745 VDDD.n1506 VDDD.n1328 0.0239375
R7746 VDDD VDDD.n1111 0.0239375
R7747 VDDD.n1523 VDDD.n1317 0.0239375
R7748 VDDD.n1558 VDDD.n1520 0.0239375
R7749 VDDD.n1724 VDDD.n1722 0.0239375
R7750 VDDD.n1764 VDDD.n1716 0.0239375
R7751 VDDD.n1924 VDDD.n1922 0.0239375
R7752 VDDD.n1956 VDDD.n1912 0.0239375
R7753 VDDD.n2330 VDDD.n1964 0.0239375
R7754 VDDD.n2324 VDDD.n1966 0.0239375
R7755 VDDD.n169 VDDD.n167 0.0239375
R7756 VDDD.n202 VDDD.n118 0.0239375
R7757 VDDD.n244 VDDD 0.0226354
R7758 VDDD.n3660 VDDD 0.0226354
R7759 VDDD VDDD.n226 0.0226354
R7760 VDDD.n3515 VDDD 0.0226354
R7761 VDDD.n3554 VDDD 0.0226354
R7762 VDDD.n3566 VDDD 0.0226354
R7763 VDDD.n3578 VDDD 0.0226354
R7764 VDDD VDDD.n3599 0.0226354
R7765 VDDD.n3640 VDDD 0.0226354
R7766 VDDD VDDD.n277 0.0226354
R7767 VDDD.n408 VDDD 0.0226354
R7768 VDDD VDDD.n418 0.0226354
R7769 VDDD.n453 VDDD 0.0226354
R7770 VDDD VDDD.n466 0.0226354
R7771 VDDD VDDD.n477 0.0226354
R7772 VDDD VDDD.n495 0.0226354
R7773 VDDD.n550 VDDD 0.0226354
R7774 VDDD.n547 VDDD 0.0226354
R7775 VDDD.n536 VDDD 0.0226354
R7776 VDDD.n533 VDDD 0.0226354
R7777 VDDD.n3466 VDDD 0.0226354
R7778 VDDD.n3444 VDDD 0.0226354
R7779 VDDD.n3437 VDDD 0.0226354
R7780 VDDD.n3432 VDDD 0.0226354
R7781 VDDD VDDD.n3312 0.0226354
R7782 VDDD VDDD.n3327 0.0226354
R7783 VDDD.n3394 VDDD 0.0226354
R7784 VDDD VDDD.n3342 0.0226354
R7785 VDDD.n3092 VDDD 0.0226354
R7786 VDDD.n3087 VDDD 0.0226354
R7787 VDDD.n732 VDDD 0.0226354
R7788 VDDD.n725 VDDD 0.0226354
R7789 VDDD VDDD.n3107 0.0226354
R7790 VDDD.n3122 VDDD 0.0226354
R7791 VDDD.n3153 VDDD 0.0226354
R7792 VDDD.n3159 VDDD 0.0226354
R7793 VDDD.n618 VDDD 0.0226354
R7794 VDDD.n612 VDDD 0.0226354
R7795 VDDD.n608 VDDD 0.0226354
R7796 VDDD.n3246 VDDD 0.0226354
R7797 VDDD.n3238 VDDD 0.0226354
R7798 VDDD VDDD.n3178 0.0226354
R7799 VDDD.n3197 VDDD 0.0226354
R7800 VDDD.n794 VDDD 0.0226354
R7801 VDDD.n3047 VDDD 0.0226354
R7802 VDDD VDDD.n769 0.0226354
R7803 VDDD.n3033 VDDD 0.0226354
R7804 VDDD.n1053 VDDD 0.0226354
R7805 VDDD VDDD.n874 0.0226354
R7806 VDDD.n1036 VDDD 0.0226354
R7807 VDDD VDDD.n878 0.0226354
R7808 VDDD.n1030 VDDD 0.0226354
R7809 VDDD.n988 VDDD 0.0226354
R7810 VDDD.n982 VDDD 0.0226354
R7811 VDDD.n981 VDDD 0.0226354
R7812 VDDD.n946 VDDD 0.0226354
R7813 VDDD.n1470 VDDD 0.0226354
R7814 VDDD.n1495 VDDD 0.0226354
R7815 VDDD.n1486 VDDD 0.0226354
R7816 VDDD.n1485 VDDD 0.0226354
R7817 VDDD.n1432 VDDD 0.0226354
R7818 VDDD.n1361 VDDD 0.0226354
R7819 VDDD.n1414 VDDD 0.0226354
R7820 VDDD.n3012 VDDD 0.0226354
R7821 VDDD.n2997 VDDD 0.0226354
R7822 VDDD.n2996 VDDD 0.0226354
R7823 VDDD.n2977 VDDD 0.0226354
R7824 VDDD.n1220 VDDD 0.0226354
R7825 VDDD.n1200 VDDD 0.0226354
R7826 VDDD.n1180 VDDD 0.0226354
R7827 VDDD.n1549 VDDD 0.0226354
R7828 VDDD.n1546 VDDD 0.0226354
R7829 VDDD.n1538 VDDD 0.0226354
R7830 VDDD VDDD.n2782 0.0226354
R7831 VDDD.n2783 VDDD 0.0226354
R7832 VDDD VDDD.n2789 0.0226354
R7833 VDDD.n2790 VDDD 0.0226354
R7834 VDDD.n2857 VDDD 0.0226354
R7835 VDDD.n2849 VDDD 0.0226354
R7836 VDDD.n2942 VDDD 0.0226354
R7837 VDDD.n2941 VDDD 0.0226354
R7838 VDDD.n2937 VDDD 0.0226354
R7839 VDDD VDDD.n2883 0.0226354
R7840 VDDD.n1787 VDDD 0.0226354
R7841 VDDD VDDD.n1717 0.0226354
R7842 VDDD.n1746 VDDD 0.0226354
R7843 VDDD.n1738 VDDD 0.0226354
R7844 VDDD.n1851 VDDD 0.0226354
R7845 VDDD.n1835 VDDD 0.0226354
R7846 VDDD.n1831 VDDD 0.0226354
R7847 VDDD.n2702 VDDD 0.0226354
R7848 VDDD.n1599 VDDD 0.0226354
R7849 VDDD VDDD.n1605 0.0226354
R7850 VDDD.n1606 VDDD 0.0226354
R7851 VDDD.n2679 VDDD 0.0226354
R7852 VDDD.n2675 VDDD 0.0226354
R7853 VDDD.n2636 VDDD 0.0226354
R7854 VDDD.n1944 VDDD 0.0226354
R7855 VDDD.n1943 VDDD 0.0226354
R7856 VDDD VDDD.n2411 0.0226354
R7857 VDDD.n1658 VDDD 0.0226354
R7858 VDDD.n2489 VDDD 0.0226354
R7859 VDDD.n2573 VDDD 0.0226354
R7860 VDDD.n2559 VDDD 0.0226354
R7861 VDDD VDDD.n1645 0.0226354
R7862 VDDD.n2537 VDDD 0.0226354
R7863 VDDD.n2517 VDDD 0.0226354
R7864 VDDD.n2320 VDDD 0.0226354
R7865 VDDD VDDD.n1973 0.0226354
R7866 VDDD.n2297 VDDD 0.0226354
R7867 VDDD VDDD.n2082 0.0226354
R7868 VDDD.n2083 VDDD 0.0226354
R7869 VDDD.n2123 VDDD 0.0226354
R7870 VDDD.n2150 VDDD 0.0226354
R7871 VDDD.n2159 VDDD 0.0226354
R7872 VDDD.n2185 VDDD 0.0226354
R7873 VDDD VDDD.n2227 0.0226354
R7874 VDDD VDDD.n2024 0.0226354
R7875 VDDD.n2272 VDDD 0.0226354
R7876 VDDD.n2252 VDDD 0.0226354
R7877 VDDD.n145 VDDD 0.0226354
R7878 VDDD VDDD.n119 0.0226354
R7879 VDDD.n179 VDDD 0.0226354
R7880 VDDD VDDD.n49 0.0226354
R7881 VDDD.n96 VDDD 0.0226354
R7882 VDDD.n3717 VDDD 0.0226354
R7883 VDDD.n3734 VDDD 0.0226354
R7884 VDDD.n3779 VDDD 0.0226354
R7885 VDDD.n3804 VDDD 0.0226354
R7886 VDDD VDDD.n3825 0.0226354
R7887 VDDD VDDD.n3832 0.0226354
R7888 VDDD.n3577 VDDD 0.0213333
R7889 VDDD VDDD.n3460 0.0213333
R7890 VDDD.n3316 VDDD 0.0213333
R7891 VDDD VDDD.n3167 0.0213333
R7892 VDDD.n1046 VDDD 0.0213333
R7893 VDDD.n1110 VDDD 0.0213333
R7894 VDDD.n2850 VDDD 0.0213333
R7895 VDDD VDDD.n1571 0.0213333
R7896 VDDD.n2482 VDDD 0.0213333
R7897 VDDD.n2158 VDDD 0.0213333
R7898 VDDD.n3725 VDDD 0.0213333
R7899 VDDD.n3514 VDDD.n3513 0.0187292
R7900 VDDD.n3516 VDDD.n3515 0.0187292
R7901 VDDD.n3286 VDDD.n3285 0.0187292
R7902 VDDD.n488 VDDD.n483 0.0187292
R7903 VDDD.n3108 VDDD.n663 0.0187292
R7904 VDDD.n3112 VDDD.n3111 0.0187292
R7905 VDDD.n3026 VDDD.n3025 0.0187292
R7906 VDDD.n830 VDDD.n821 0.0187292
R7907 VDDD.n1428 VDDD.n1427 0.0187292
R7908 VDDD.n1357 VDDD.n1354 0.0187292
R7909 VDDD.n2748 VDDD.n1283 0.0187292
R7910 VDDD.n2753 VDDD.n2752 0.0187292
R7911 VDDD VDDD.n2954 0.0187292
R7912 VDDD.n1804 VDDD.n1680 0.0187292
R7913 VDDD.n1878 VDDD.n1877 0.0187292
R7914 VDDD.n2373 VDDD.n2372 0.0187292
R7915 VDDD.n2386 VDDD.n1674 0.0187292
R7916 VDDD.n2092 VDDD.n2091 0.0187292
R7917 VDDD.n2094 VDDD.n2093 0.0187292
R7918 VDDD.n3698 VDDD.n3697 0.0187292
R7919 VDDD.n61 VDDD.n53 0.0187292
R7920 VDDD.n3316 VDDD 0.0174271
R7921 VDDD VDDD.n566 0.016125
R7922 VDDD VDDD.n1239 0.016125
R7923 VDDD.n3684 VDDD.n211 0.0135208
R7924 VDDD.n3566 VDDD.n3473 0.0135208
R7925 VDDD.n438 VDDD.n386 0.0135208
R7926 VDDD.n366 VDDD.n364 0.0135208
R7927 VDDD.n698 VDDD.n690 0.0135208
R7928 VDDD.n3153 VDDD.n628 0.0135208
R7929 VDDD.n3070 VDDD.n753 0.0135208
R7930 VDDD.n865 VDDD.n860 0.0135208
R7931 VDDD.n1513 VDDD.n1325 0.0135208
R7932 VDDD.n1099 VDDD.n1097 0.0135208
R7933 VDDD.n2718 VDDD.n2717 0.0135208
R7934 VDDD.n2795 VDDD.n2794 0.0135208
R7935 VDDD.n1720 VDDD.n1711 0.0135208
R7936 VDDD.n1831 VDDD.n1566 0.0135208
R7937 VDDD.n1918 VDDD.n1907 0.0135208
R7938 VDDD.n2422 VDDD.n2421 0.0135208
R7939 VDDD.n2331 VDDD.n1963 0.0135208
R7940 VDDD.n2049 VDDD.n2047 0.0135208
R7941 VDDD.n159 VDDD.n121 0.0135208
R7942 VDDD.n45 VDDD.n43 0.0135208
R7943 VDDD.n3454 VDDD 0.0122188
R7944 VDDD VDDD.n632 0.0122188
R7945 VDDD VDDD.n1052 0.0122188
R7946 VDDD.n1106 VDDD 0.0122188
R7947 VDDD VDDD.n2856 0.0122188
R7948 VDDD.n2684 VDDD 0.0122188
R7949 VDDD VDDD.n2488 0.0122188
R7950 VDDD VDDD.n2054 0.0122188
R7951 VDDD.n3712 VDDD 0.0122188
R7952 VDDD.n3624 VDDD.n26 0.0118353
R7953 VDDD.n3574 VDDD.n41 0.0118353
R7954 VDDD.n3693 VDDD.n113 0.0118353
R7955 VDDD.n3689 VDDD.n3688 0.0118353
R7956 VDDD.n3570 VDDD 0.0109167
R7957 VDDD.n3160 VDDD 0.0109167
R7958 VDDD VDDD.n751 0.0109167
R7959 VDDD.n2954 VDDD 0.0109167
R7960 VDDD.n2703 VDDD 0.0109167
R7961 VDDD.n2572 VDDD 0.0109167
R7962 VDDD.n3531 VDDD.n3496 0.0083125
R7963 VDDD.n558 VDDD.n557 0.0083125
R7964 VDDD.n3125 VDDD.n655 0.0083125
R7965 VDDD.n1089 VDDD.n1088 0.0083125
R7966 VDDD.n1420 VDDD.n1419 0.0083125
R7967 VDDD.n2761 VDDD.n2760 0.0083125
R7968 VDDD.n1867 VDDD.n1866 0.0083125
R7969 VDDD.n2379 VDDD.n1670 0.0083125
R7970 VDDD.n2110 VDDD.n2068 0.0083125
R7971 VDDD.n110 VDDD.n109 0.0083125
R7972 VDDD VDDD.n3121 0.00701042
R7973 VDDD VDDD.n1360 0.00701042
R7974 VDDD.n1427 VDDD 0.00440625
R7975 VDDD.n3720 VDDD 0.00387838
R7976 VDDD VDDD.n3479 0.00310417
R7977 VDDD.n3476 VDDD.n3475 0.00310417
R7978 VDDD.n3619 VDDD.n3618 0.00310417
R7979 VDDD.n3461 VDDD.n3294 0.00310417
R7980 VDDD.n3417 VDDD.n3416 0.00310417
R7981 VDDD.n3168 VDDD.n623 0.00310417
R7982 VDDD.n3271 VDDD.n569 0.00310417
R7983 VDDD.n871 VDDD.n870 0.00310417
R7984 VDDD.n1010 VDDD.n1009 0.00310417
R7985 VDDD.n1107 VDDD.n1102 0.00310417
R7986 VDDD.n1145 VDDD.n1138 0.00310417
R7987 VDDD.n1256 VDDD.n1252 0.00310417
R7988 VDDD.n2959 VDDD.n1242 0.00310417
R7989 VDDD.n2691 VDDD.n2690 0.00310417
R7990 VDDD.n1627 VDDD.n1579 0.00310417
R7991 VDDD.n1652 VDDD.n1648 0.00310417
R7992 VDDD.n2577 VDDD.n1638 0.00310417
R7993 VDDD.n2051 VDDD.n2050 0.00310417
R7994 VDDD.n2204 VDDD.n2203 0.00310417
R7995 VDDD.n3714 VDDD.n3713 0.00310417
R7996 VDDD.n3772 VDDD.n3771 0.00310417
R7997 a_1835_9813.n3 a_1835_9813.n0 807.871
R7998 a_1835_9813.n4 a_1835_9813.t5 389.183
R7999 a_1835_9813.n5 a_1835_9813.n4 251.167
R8000 a_1835_9813.t0 a_1835_9813.n5 223.571
R8001 a_1835_9813.n2 a_1835_9813.t8 212.081
R8002 a_1835_9813.n1 a_1835_9813.t6 212.081
R8003 a_1835_9813.n3 a_1835_9813.n2 176.576
R8004 a_1835_9813.n4 a_1835_9813.t3 174.891
R8005 a_1835_9813.n2 a_1835_9813.t7 139.78
R8006 a_1835_9813.n1 a_1835_9813.t4 139.78
R8007 a_1835_9813.n0 a_1835_9813.t2 63.3219
R8008 a_1835_9813.n0 a_1835_9813.t1 63.3219
R8009 a_1835_9813.n2 a_1835_9813.n1 61.346
R8010 a_1835_9813.n5 a_1835_9813.n3 37.5061
R8011 a_4739_10625.n1 a_4739_10625.t3 530.01
R8012 a_4739_10625.t0 a_4739_10625.n5 421.021
R8013 a_4739_10625.n0 a_4739_10625.t7 337.171
R8014 a_4739_10625.n3 a_4739_10625.t1 280.223
R8015 a_4739_10625.n4 a_4739_10625.t6 263.173
R8016 a_4739_10625.n4 a_4739_10625.t2 227.826
R8017 a_4739_10625.n0 a_4739_10625.t5 199.762
R8018 a_4739_10625.n2 a_4739_10625.n1 170.81
R8019 a_4739_10625.n2 a_4739_10625.n0 167.321
R8020 a_4739_10625.n5 a_4739_10625.n4 152
R8021 a_4739_10625.n1 a_4739_10625.t4 141.923
R8022 a_4739_10625.n3 a_4739_10625.n2 10.8376
R8023 a_4739_10625.n5 a_4739_10625.n3 2.50485
R8024 a_4700_10499.t0 a_4700_10499.n3 370.026
R8025 a_4700_10499.n0 a_4700_10499.t3 351.356
R8026 a_4700_10499.n1 a_4700_10499.t5 334.717
R8027 a_4700_10499.n3 a_4700_10499.t1 325.971
R8028 a_4700_10499.n1 a_4700_10499.t2 309.935
R8029 a_4700_10499.n0 a_4700_10499.t4 305.683
R8030 a_4700_10499.n2 a_4700_10499.n0 16.879
R8031 a_4700_10499.n3 a_4700_10499.n2 10.8867
R8032 a_4700_10499.n2 a_4700_10499.n1 9.3005
R8033 VSSD.n3666 VSSD.n46 25423.7
R8034 VSSD.n3658 VSSD 8566
R8035 VSSD VSSD.t1393 4897.32
R8036 VSSD VSSD.t1448 4888.89
R8037 VSSD VSSD.n3397 4522.16
R8038 VSSD.n3666 VSSD.n3665 4490.81
R8039 VSSD.n3665 VSSD.n3664 4490.81
R8040 VSSD.n3664 VSSD.n3663 4490.81
R8041 VSSD.n3663 VSSD.n3662 4490.81
R8042 VSSD.n3662 VSSD.n3661 4490.81
R8043 VSSD.n3661 VSSD.n3660 4490.81
R8044 VSSD.n3660 VSSD.n3659 4490.81
R8045 VSSD.n3659 VSSD.n3658 4490.81
R8046 VSSD.n3390 VSSD.n46 4424.4
R8047 VSSD.n3391 VSSD.n3390 4424.4
R8048 VSSD.n3392 VSSD.n3391 4424.4
R8049 VSSD.n3393 VSSD.n3392 4424.4
R8050 VSSD.n3394 VSSD.n3393 4424.4
R8051 VSSD.n3395 VSSD.n3394 4424.4
R8052 VSSD.n3396 VSSD.n3395 4424.4
R8053 VSSD.n3397 VSSD.n3396 4424.4
R8054 VSSD.t1448 VSSD 4408.43
R8055 VSSD.t1393 VSSD 4408.43
R8056 VSSD VSSD.t1490 4408.43
R8057 VSSD VSSD.t1473 4408.43
R8058 VSSD VSSD.t1434 4408.43
R8059 VSSD.t1195 VSSD.t1454 3101.92
R8060 VSSD VSSD.t1505 2857.47
R8061 VSSD.t1431 VSSD 2857.47
R8062 VSSD VSSD.t1310 2562.45
R8063 VSSD.t306 VSSD.t1269 2410.73
R8064 VSSD.t123 VSSD.t1367 2410.73
R8065 VSSD.t311 VSSD.t1318 2410.73
R8066 VSSD.t1493 VSSD.t1378 2326.44
R8067 VSSD.t1094 VSSD.t129 2149.43
R8068 VSSD.t901 VSSD.t919 2149.43
R8069 VSSD.t520 VSSD.t525 2149.43
R8070 VSSD.t344 VSSD.t751 2149.43
R8071 VSSD VSSD.t869 2149.43
R8072 VSSD.t78 VSSD.t1705 2149.43
R8073 VSSD.t111 VSSD.t1721 2149.43
R8074 VSSD.t1578 VSSD.t1623 2149.43
R8075 VSSD.t1618 VSSD.t1106 2149.43
R8076 VSSD.t70 VSSD.t518 2149.43
R8077 VSSD.t817 VSSD.t943 2149.43
R8078 VSSD.t1280 VSSD 2081.99
R8079 VSSD.t1378 VSSD 2081.99
R8080 VSSD.t342 VSSD.t1510 2022.99
R8081 VSSD.t1829 VSSD.t763 1980.84
R8082 VSSD.n3389 VSSD.t1459 1938.7
R8083 VSSD.n3056 VSSD.t1298 1938.7
R8084 VSSD VSSD.t528 1845.98
R8085 VSSD.t443 VSSD 1837.55
R8086 VSSD VSSD.t1370 1795.4
R8087 VSSD.t1505 VSSD 1795.4
R8088 VSSD VSSD.t1516 1795.4
R8089 VSSD VSSD.t1547 1786.97
R8090 VSSD VSSD.t1216 1786.97
R8091 VSSD.t1295 VSSD 1786.97
R8092 VSSD.t982 VSSD.t435 1753.26
R8093 VSSD.t1018 VSSD.t304 1753.26
R8094 VSSD.t1587 VSSD.t340 1753.26
R8095 VSSD.t1762 VSSD.t1759 1753.26
R8096 VSSD.t13 VSSD.t1172 1753.26
R8097 VSSD.t718 VSSD.t1843 1753.26
R8098 VSSD.t80 VSSD.t1820 1753.26
R8099 VSSD.t825 VSSD.t986 1753.26
R8100 VSSD.t1726 VSSD.t313 1753.26
R8101 VSSD.t538 VSSD.t182 1753.26
R8102 VSSD.t961 VSSD.t1712 1719.54
R8103 VSSD.t650 VSSD.t1470 1711.11
R8104 VSSD.t1272 VSSD 1702.68
R8105 VSSD VSSD.t1213 1702.68
R8106 VSSD VSSD.t1321 1702.68
R8107 VSSD VSSD.t1422 1702.68
R8108 VSSD VSSD.t1437 1702.68
R8109 VSSD VSSD.t1254 1702.68
R8110 VSSD VSSD.t1263 1702.68
R8111 VSSD.t1462 VSSD 1702.68
R8112 VSSD VSSD.t1228 1702.68
R8113 VSSD.t177 VSSD.t1275 1601.53
R8114 VSSD.t1440 VSSD.t632 1601.53
R8115 VSSD VSSD.t1085 1559.39
R8116 VSSD.t1537 VSSD.t1242 1550.96
R8117 VSSD.t1216 VSSD.t1354 1550.96
R8118 VSSD.t1283 VSSD.t1443 1550.96
R8119 VSSD.t1357 VSSD.t1198 1550.96
R8120 VSSD.t1390 VSSD.t1295 1550.96
R8121 VSSD.n672 VSSD.t1373 1550.96
R8122 VSSD.t1516 VSSD.t1431 1550.96
R8123 VSSD.t1334 VSSD.t641 1534.1
R8124 VSSD.t1465 VSSD.t716 1534.1
R8125 VSSD.t1814 VSSD.t1248 1534.1
R8126 VSSD.t488 VSSD 1525.67
R8127 VSSD.t656 VSSD 1483.52
R8128 VSSD VSSD.t246 1432.95
R8129 VSSD VSSD.t1405 1407.66
R8130 VSSD VSSD.t1411 1407.66
R8131 VSSD VSSD.t1222 1407.66
R8132 VSSD VSSD.t1231 1407.66
R8133 VSSD VSSD.t1351 1407.66
R8134 VSSD VSSD.t1479 1407.66
R8135 VSSD VSSD.t1257 1407.66
R8136 VSSD VSSD.t1234 1407.66
R8137 VSSD VSSD.t1301 1407.66
R8138 VSSD.t1029 VSSD.t185 1399.23
R8139 VSSD.t730 VSSD.t1813 1399.23
R8140 VSSD.t66 VSSD.t12 1399.23
R8141 VSSD.t952 VSSD.t1030 1399.23
R8142 VSSD.t275 VSSD.t1819 1399.23
R8143 VSSD.t268 VSSD.t532 1399.23
R8144 VSSD.t862 VSSD.t724 1399.23
R8145 VSSD.t550 VSSD.t227 1399.23
R8146 VSSD.t103 VSSD.t589 1399.23
R8147 VSSD.t790 VSSD.t1176 1399.23
R8148 VSSD.t1692 VSSD.t580 1399.23
R8149 VSSD.t1807 VSSD.t51 1399.23
R8150 VSSD.t1127 VSSD.t1027 1399.23
R8151 VSSD.t964 VSSD.n1617 1382.38
R8152 VSSD.t1083 VSSD.t1775 1373.95
R8153 VSSD.t839 VSSD.t637 1373.95
R8154 VSSD.t1119 VSSD.t627 1373.95
R8155 VSSD.t613 VSSD.t837 1314.94
R8156 VSSD VSSD.t1459 1306.51
R8157 VSSD.t1242 VSSD 1306.51
R8158 VSSD.t1547 VSSD 1306.51
R8159 VSSD.t1354 VSSD 1306.51
R8160 VSSD.t1348 VSSD 1306.51
R8161 VSSD.t1269 VSSD 1306.51
R8162 VSSD VSSD.t1283 1306.51
R8163 VSSD.t1298 VSSD 1306.51
R8164 VSSD.t1286 VSSD 1306.51
R8165 VSSD.t1367 VSSD 1306.51
R8166 VSSD VSSD.t1357 1306.51
R8167 VSSD.t1318 VSSD 1306.51
R8168 VSSD VSSD.t1195 1306.51
R8169 VSSD.t1408 VSSD 1306.51
R8170 VSSD.t1769 VSSD 1289.66
R8171 VSSD.t1189 VSSD 1289.66
R8172 VSSD.t298 VSSD.t1089 1281.23
R8173 VSSD.t639 VSSD.t1593 1255.94
R8174 VSSD.t410 VSSD.t504 1255.94
R8175 VSSD.t1058 VSSD.t1714 1255.94
R8176 VSSD.t1139 VSSD.t980 1255.94
R8177 VSSD.t308 VSSD.t489 1255.94
R8178 VSSD.t1591 VSSD.t183 1255.94
R8179 VSSD.t675 VSSD.t478 1255.94
R8180 VSSD.t1682 VSSD.t1764 1255.94
R8181 VSSD.t590 VSSD.t506 1255.94
R8182 VSSD.t569 VSSD.t1670 1255.94
R8183 VSSD.t558 VSSD.t404 1255.94
R8184 VSSD.t669 VSSD.t1648 1255.94
R8185 VSSD.t331 VSSD.t1660 1255.94
R8186 VSSD.t1778 VSSD.t805 1255.94
R8187 VSSD.t500 VSSD.n171 1247.51
R8188 VSSD.t349 VSSD 1239.08
R8189 VSSD.t1192 VSSD.t581 1230.65
R8190 VSSD.t1396 VSSD.t760 1230.65
R8191 VSSD.t1425 VSSD.t121 1230.65
R8192 VSSD.t811 VSSD 1230.65
R8193 VSSD.t1245 VSSD.t935 1230.65
R8194 VSSD.t1646 VSSD.t1343 1230.65
R8195 VSSD.t127 VSSD.t110 1213.79
R8196 VSSD.t202 VSSD.t992 1213.79
R8197 VSSD.n933 VSSD.n866 1198.25
R8198 VSSD.n3305 VSSD.n3304 1198.25
R8199 VSSD.n2693 VSSD.n1329 1198.25
R8200 VSSD.n2456 VSSD.n2455 1198.25
R8201 VSSD.n1489 VSSD.n1482 1198.25
R8202 VSSD.n2106 VSSD.n2105 1198.25
R8203 VSSD.n3408 VSSD.n3398 1198.25
R8204 VSSD.n3473 VSSD.n96 1198.25
R8205 VSSD.n3534 VSSD.n73 1198.25
R8206 VSSD.n3657 VSSD.n3656 1198.25
R8207 VSSD.n248 VSSD.n214 1198.25
R8208 VSSD.n2454 VSSD.n2453 1197.79
R8209 VSSD.n3303 VSSD.n3302 1195.68
R8210 VSSD.n311 VSSD.n249 1195.68
R8211 VSSD.n3667 VSSD.n15 1194.5
R8212 VSSD.n673 VSSD.n672 1194.5
R8213 VSSD.n826 VSSD.n825 1194.5
R8214 VSSD.n987 VSSD.n827 1194.5
R8215 VSSD.n3389 VSSD.n3388 1194.5
R8216 VSSD.n1295 VSSD.n1294 1194.5
R8217 VSSD.n1296 VSSD.t1289 1194.5
R8218 VSSD.n3116 VSSD.n3056 1194.5
R8219 VSSD.n2951 VSSD.n1099 1194.5
R8220 VSSD.n3055 VSSD.n3054 1194.5
R8221 VSSD.n2869 VSSD.n2861 1194.5
R8222 VSSD.n2770 VSSD.n2694 1194.5
R8223 VSSD.t958 VSSD.n2692 1194.5
R8224 VSSD.n2567 VSSD.n2566 1194.5
R8225 VSSD.n1481 VSSD.n1382 1194.5
R8226 VSSD.n2215 VSSD.n2140 1194.5
R8227 VSSD.n2280 VSSD.n2107 1194.5
R8228 VSSD.n1971 VSSD.n1970 1194.5
R8229 VSSD.n1769 VSSD.n1693 1194.5
R8230 VSSD.n1829 VSSD.n1657 1194.5
R8231 VSSD.n1616 VSSD.n1615 1194.5
R8232 VSSD.n1888 VSSD.n1617 1194.5
R8233 VSSD.n422 VSSD.n171 1194.5
R8234 VSSD.n490 VSSD.n489 1194.5
R8235 VSSD VSSD.t607 1188.51
R8236 VSSD.t1327 VSSD.t1482 1163.22
R8237 VSSD.n2861 VSSD.t1402 1163.22
R8238 VSSD.t267 VSSD.t310 1163.22
R8239 VSSD.t463 VSSD.t98 1163.22
R8240 VSSD.t1260 VSSD.t1519 1163.22
R8241 VSSD.t1476 VSSD.n1616 1163.22
R8242 VSSD.t1513 VSSD.t1225 1163.22
R8243 VSSD.n1693 VSSD.t1384 1163.22
R8244 VSSD.t883 VSSD.t1799 1146.36
R8245 VSSD.t34 VSSD.t695 1146.36
R8246 VSSD.t853 VSSD.t917 1112.64
R8247 VSSD.t1141 VSSD.t578 1112.64
R8248 VSSD.t1848 VSSD.t1589 1112.64
R8249 VSSD.t1656 VSSD.t990 1112.64
R8250 VSSD.t399 VSSD.t162 1112.64
R8251 VSSD.t514 VSSD.t293 1112.64
R8252 VSSD.t788 VSSD.t269 1112.64
R8253 VSSD.t1131 VSSD.t171 1112.64
R8254 VSSD.t1680 VSSD.t329 1112.64
R8255 VSSD.t115 VSSD.t242 1112.64
R8256 VSSD.t234 VSSD.t446 1112.64
R8257 VSSD.t236 VSSD.t771 1112.64
R8258 VSSD.t712 VSSD.t897 1112.64
R8259 VSSD.t1674 VSSD.t424 1112.64
R8260 VSSD.t62 VSSD.t889 1112.64
R8261 VSSD.t319 VSSD.t493 1112.64
R8262 VSSD.t945 VSSD.t512 1112.64
R8263 VSSD.t416 VSSD 1104.21
R8264 VSSD.t198 VSSD 1104.21
R8265 VSSD VSSD.t1816 1104.21
R8266 VSSD VSSD.t8 1095.79
R8267 VSSD.t1672 VSSD.t264 1053.64
R8268 VSSD VSSD.t1219 1048.99
R8269 VSSD VSSD.t1399 1048.99
R8270 VSSD VSSD.t1183 1048.99
R8271 VSSD VSSD.t1532 1048.99
R8272 VSSD VSSD.t1304 1048.99
R8273 VSSD VSSD.t1555 1048.99
R8274 VSSD.t1522 VSSD 1048.99
R8275 VSSD.t1550 VSSD 1047.19
R8276 VSSD.t1676 VSSD.t667 1036.78
R8277 VSSD.t1443 VSSD 1011.49
R8278 VSSD VSSD.t1210 1011.49
R8279 VSSD.t1502 VSSD 1011.49
R8280 VSSD.t442 VSSD.t336 1003.07
R8281 VSSD.t857 VSSD.t499 1003.07
R8282 VSSD.t1251 VSSD.t868 994.636
R8283 VSSD.t1635 VSSD.t1201 994.636
R8284 VSSD.t773 VSSD.t1062 977.779
R8285 VSSD.t947 VSSD.t346 977.779
R8286 VSSD.t725 VSSD.t1040 977.779
R8287 VSSD.t1219 VSSD 944.277
R8288 VSSD.t1399 VSSD 944.277
R8289 VSSD.t1183 VSSD 944.277
R8290 VSSD.t1532 VSSD 944.277
R8291 VSSD.t1304 VSSD 944.277
R8292 VSSD.t1555 VSSD 944.277
R8293 VSSD VSSD.t1550 944.277
R8294 VSSD VSSD.t1522 944.277
R8295 VSSD.t474 VSSD.t228 944.062
R8296 VSSD.t452 VSSD.t1662 944.062
R8297 VSSD.t1684 VSSD.t114 944.062
R8298 VSSD VSSD.n3055 927.203
R8299 VSSD.n2566 VSSD 927.203
R8300 VSSD VSSD.n2693 927.203
R8301 VSSD VSSD.n2107 927.203
R8302 VSSD VSSD.n1657 927.203
R8303 VSSD VSSD.n671 927.203
R8304 VSSD.t1028 VSSD.t1149 918.774
R8305 VSSD.t719 VSSD.t1031 918.774
R8306 VSSD.t1405 VSSD 918.774
R8307 VSSD.t1289 VSSD 918.774
R8308 VSSD.t139 VSSD.t156 918.774
R8309 VSSD.t1482 VSSD 918.774
R8310 VSSD.n3303 VSSD 918.774
R8311 VSSD.t1411 VSSD 918.774
R8312 VSSD.t1021 VSSD.t723 918.774
R8313 VSSD.t549 VSSD.t523 918.774
R8314 VSSD.t1510 VSSD 918.774
R8315 VSSD.n2694 VSSD 918.774
R8316 VSSD.t1222 VSSD 918.774
R8317 VSSD.t775 VSSD.t50 918.774
R8318 VSSD.t1231 VSSD 918.774
R8319 VSSD VSSD.t1260 918.774
R8320 VSSD.t1126 VSSD.t942 918.774
R8321 VSSD.t1351 VSSD 918.774
R8322 VSSD.t102 VSSD.t297 918.774
R8323 VSSD.t471 VSSD.t445 918.774
R8324 VSSD VSSD.t1513 918.774
R8325 VSSD.t477 VSSD.t398 918.774
R8326 VSSD.t831 VSSD.t707 918.774
R8327 VSSD.n1693 VSSD 918.774
R8328 VSSD.t1479 VSSD 918.774
R8329 VSSD.n249 VSSD 918.774
R8330 VSSD.t1257 VSSD 918.774
R8331 VSSD VSSD.t1307 918.774
R8332 VSSD.t1373 VSSD 918.774
R8333 VSSD.t960 VSSD.t1737 918.774
R8334 VSSD.n3668 VSSD 918.774
R8335 VSSD.t672 VSSD.t1 918.774
R8336 VSSD.t1234 VSSD 918.774
R8337 VSSD.t1301 VSSD 918.774
R8338 VSSD.t556 VSSD.t958 910.346
R8339 VSSD.t1068 VSSD.t1105 910.346
R8340 VSSD.t246 VSSD 893.487
R8341 VSSD.t748 VSSD 885.058
R8342 VSSD.t1112 VSSD.t100 876.629
R8343 VSSD.t1596 VSSD.t1414 876.629
R8344 VSSD.t170 VSSD.t1696 876.629
R8345 VSSD.t1292 VSSD.t1771 859.77
R8346 VSSD.t75 VSSD.t1493 859.77
R8347 VSSD.t929 VSSD.t1189 859.77
R8348 VSSD.t1454 VSSD.t586 859.77
R8349 VSSD.n3390 VSSD 851.341
R8350 VSSD.n3391 VSSD 851.341
R8351 VSSD.n3392 VSSD 851.341
R8352 VSSD.n3393 VSSD 851.341
R8353 VSSD.n3394 VSSD 851.341
R8354 VSSD.t458 VSSD 851.341
R8355 VSSD.t677 VSSD.t533 851.341
R8356 VSSD.n3395 VSSD 851.341
R8357 VSSD.n3396 VSSD 851.341
R8358 VSSD.n3397 VSSD 851.341
R8359 VSSD VSSD.n46 851.341
R8360 VSSD.t791 VSSD.t83 842.913
R8361 VSSD.t685 VSSD.t1598 842.913
R8362 VSSD.t43 VSSD.t933 842.913
R8363 VSSD.t175 VSSD.t155 842.913
R8364 VSSD.t195 VSSD.t194 834.484
R8365 VSSD.t666 VSSD.t157 834.484
R8366 VSSD.t156 VSSD.t853 834.484
R8367 VSSD.t578 VSSD.t1167 834.484
R8368 VSSD.t293 VSSD.t549 834.484
R8369 VSSD.t171 VSSD.t441 834.484
R8370 VSSD.t849 VSSD.t677 834.484
R8371 VSSD.t329 VSSD.t775 834.484
R8372 VSSD.t951 VSSD.t115 834.484
R8373 VSSD.t942 VSSD.t748 834.484
R8374 VSSD.t446 VSSD.t1806 834.484
R8375 VSSD.t771 VSSD.t225 834.484
R8376 VSSD.t117 VSSD.t122 834.484
R8377 VSSD.t984 VSSD.t1753 834.484
R8378 VSSD.t1746 VSSD.t175 834.484
R8379 VSSD.t1097 VSSD.t64 834.484
R8380 VSSD.t476 VSSD.t1610 834.484
R8381 VSSD.t1 VSSD.t945 834.484
R8382 VSSD.t1419 VSSD.t1577 826.054
R8383 VSSD.t1032 VSSD.t1408 826.054
R8384 VSSD.t1149 VSSD.t639 809.196
R8385 VSSD.t100 VSSD.t738 809.196
R8386 VSSD.t1811 VSSD.t131 809.196
R8387 VSSD.t1793 VSSD.t730 809.196
R8388 VSSD.t664 VSSD.t448 809.196
R8389 VSSD.t1714 VSSD.t719 809.196
R8390 VSSD.t206 VSSD.t809 809.196
R8391 VSSD.t1752 VSSD.t810 809.196
R8392 VSSD.t980 VSSD.t139 809.196
R8393 VSSD.t532 VSSD.t1023 809.196
R8394 VSSD.t522 VSSD.t1168 809.196
R8395 VSSD.t1617 VSSD.t308 809.196
R8396 VSSD.t183 VSSD.t1021 809.196
R8397 VSSD.t724 VSSD.t1833 809.196
R8398 VSSD.t524 VSSD.t550 809.196
R8399 VSSD.t523 VSSD.t675 809.196
R8400 VSSD.t729 VSSD.t334 809.196
R8401 VSSD.t1764 VSSD.t1742 809.196
R8402 VSSD.t1063 VSSD.t1171 809.196
R8403 VSSD.t77 VSSD.t590 809.196
R8404 VSSD.t885 VSSD.t2 809.196
R8405 VSSD.t450 VSSD.t569 809.196
R8406 VSSD.t1090 VSSD.t39 809.196
R8407 VSSD.t49 VSSD.t790 809.196
R8408 VSSD.t50 VSSD.t1841 809.196
R8409 VSSD VSSD.t254 809.196
R8410 VSSD.t580 VSSD.t161 809.196
R8411 VSSD.t1577 VSSD.t669 809.196
R8412 VSSD.t1620 VSSD.t226 809.196
R8413 VSSD.t1614 VSSD.t331 809.196
R8414 VSSD.t536 VSSD.t562 809.196
R8415 VSSD.t805 VSSD.t960 809.196
R8416 VSSD.t1027 VSSD.t517 809.196
R8417 VSSD.t125 VSSD.t74 809.196
R8418 VSSD.t1035 VSSD.t1797 809.196
R8419 VSSD.t584 VSSD.t72 809.196
R8420 VSSD.t0 VSSD.t671 809.196
R8421 VSSD.t1023 VSSD.t901 800.766
R8422 VSSD.t525 VSSD.t522 800.766
R8423 VSSD.t751 VSSD.t524 800.766
R8424 VSSD.t1705 VSSD.t1063 800.766
R8425 VSSD.t776 VSSD.t873 800.766
R8426 VSSD.t1085 VSSD.t49 800.766
R8427 VSSD.t1117 VSSD.t325 800.766
R8428 VSSD.t1721 VSSD.t551 800.766
R8429 VSSD.t161 VSSD.t1108 800.766
R8430 VSSD.t999 VSSD.t1823 800.766
R8431 VSSD.t765 VSSD.t543 800.766
R8432 VSSD.t1623 VSSD.t1580 800.766
R8433 VSSD.t362 VSSD.t300 800.766
R8434 VSSD.t1106 VSSD.t1620 800.766
R8435 VSSD.t1678 VSSD 800.766
R8436 VSSD.t173 VSSD.t1034 800.766
R8437 VSSD.t998 VSSD.t1740 800.766
R8438 VSSD.t671 VSSD.t817 800.766
R8439 VSSD.t843 VSSD.t495 792.337
R8440 VSSD.t475 VSSD.t1811 792.337
R8441 VSSD.t244 VSSD.t1008 783.909
R8442 VSSD.t230 VSSD.t378 783.909
R8443 VSSD.t438 VSSD.t315 783.909
R8444 VSSD.t1310 VSSD.t1348 775.48
R8445 VSSD.t338 VSSD.t1083 775.48
R8446 VSSD.t1818 VSSD.t1571 775.48
R8447 VSSD.t1735 VSSD.t1576 775.48
R8448 VSSD.t1165 VSSD.t700 775.48
R8449 VSSD.t1734 VSSD.t548 775.48
R8450 VSSD.t1777 VSSD.t1794 775.48
R8451 VSSD.t6 VSSD.t614 775.48
R8452 VSSD.t1210 VSSD.t1286 775.48
R8453 VSSD.t1079 VSSD.t971 775.48
R8454 VSSD.t1720 VSSD.t881 775.48
R8455 VSSD.t203 VSSD.t432 775.48
R8456 VSSD.t903 VSSD.t1789 775.48
R8457 VSSD.t1711 VSSD.t431 775.48
R8458 VSSD.t636 VSSD.t882 775.48
R8459 VSSD.t108 VSSD.t839 775.48
R8460 VSSD.t1370 VSSD.t1280 775.48
R8461 VSSD.t398 VSSD.t832 775.48
R8462 VSSD.t396 VSSD.t831 775.48
R8463 VSSD.t1755 VSSD.t352 775.48
R8464 VSSD.t1694 VSSD.t1121 775.48
R8465 VSSD.t472 VSSD.t855 775.48
R8466 VSSD.t1718 VSSD.t582 775.48
R8467 VSSD.t473 VSSD.t856 775.48
R8468 VSSD.t1768 VSSD.t1118 775.48
R8469 VSSD.t627 VSSD.t30 775.48
R8470 VSSD.t1593 VSSD.t1026 767.051
R8471 VSSD.t1060 VSSD.t682 767.051
R8472 VSSD.t868 VSSD.t1058 767.051
R8473 VSSD.t435 VSSD.t1139 767.051
R8474 VSSD.t489 VSSD.t1018 767.051
R8475 VSSD.t863 VSSD.t1591 767.051
R8476 VSSD.t965 VSSD.t266 767.051
R8477 VSSD.t99 VSSD.t289 767.051
R8478 VSSD.t987 VSSD.t252 767.051
R8479 VSSD.t1062 VSSD.t260 767.051
R8480 VSSD.t478 VSSD.t1587 767.051
R8481 VSSD.t346 VSSD.t1137 767.051
R8482 VSSD.t288 VSSD.t166 767.051
R8483 VSSD.t1759 VSSD.t1682 767.051
R8484 VSSD.t506 VSSD.t13 767.051
R8485 VSSD.t1175 VSSD.t244 767.051
R8486 VSSD.t221 VSSD.t1716 767.051
R8487 VSSD.t1666 VSSD.t1635 767.051
R8488 VSSD.t254 VSSD.t718 767.051
R8489 VSSD.t401 VSSD.t230 767.051
R8490 VSSD.t753 VSSD.t211 767.051
R8491 VSSD.t1823 VSSD.t753 767.051
R8492 VSSD.t1154 VSSD.t558 767.051
R8493 VSSD.t315 VSSD.t1736 767.051
R8494 VSSD.t1648 VSSD.t349 767.051
R8495 VSSD.t1660 VSSD.t1726 767.051
R8496 VSSD.t256 VSSD.t725 767.051
R8497 VSSD.t238 VSSD.t67 767.051
R8498 VSSD.t897 VSSD.t516 767.051
R8499 VSSD.t963 VSSD.t1674 767.051
R8500 VSSD.t182 VSSD.t1678 767.051
R8501 VSSD.t1704 VSSD.t1778 767.051
R8502 VSSD.t1150 VSSD.t871 758.621
R8503 VSSD.t504 VSSD.t530 758.621
R8504 VSSD.t899 VSSD.t1251 758.621
R8505 VSSD.t1825 VSSD 758.621
R8506 VSSD.t1201 VSSD.t815 758.621
R8507 VSSD.t611 VSSD.t733 758.621
R8508 VSSD VSSD.t954 758.621
R8509 VSSD.t915 VSSD.t776 750.192
R8510 VSSD.t1640 VSSD.t1117 750.192
R8511 VSSD VSSD.t1154 750.192
R8512 VSSD.t543 VSSD.t366 750.192
R8513 VSSD VSSD.t1654 750.192
R8514 VSSD.t683 VSSD.t81 741.763
R8515 VSSD.t684 VSSD.t395 741.763
R8516 VSSD.t1803 VSSD.t996 741.763
R8517 VSSD.t1128 VSSD.t604 741.763
R8518 VSSD.t743 VSSD.t1717 741.763
R8519 VSSD.t41 VSSD.t1751 741.763
R8520 VSSD.t179 VSSD 733.333
R8521 VSSD.t652 VSSD.t819 724.904
R8522 VSSD.t819 VSSD.t372 724.904
R8523 VSSD.t374 VSSD.t90 724.904
R8524 VSSD.t90 VSSD.t370 724.904
R8525 VSSD.t370 VSSD.t92 724.904
R8526 VSSD.t658 VSSD.t88 724.904
R8527 VSSD.t88 VSSD.t821 724.904
R8528 VSSD.t821 VSSD.t660 724.904
R8529 VSSD.t823 VSSD.t662 724.904
R8530 VSSD.t186 VSSD.t190 724.904
R8531 VSSD.t135 VSSD.t186 724.904
R8532 VSSD.t137 VSSD.t188 724.904
R8533 VSSD.t1145 VSSD.t133 724.904
R8534 VSSD.t1697 VSSD.t1690 724.904
R8535 VSSD.t484 VSSD.t609 724.904
R8536 VSSD.t609 VSSD.t284 724.904
R8537 VSSD.t286 VSSD.t1606 724.904
R8538 VSSD.t1604 VSSD.t1608 724.904
R8539 VSSD.t486 VSSD.t276 724.904
R8540 VSSD.t26 VSSD.t605 724.904
R8541 VSSD.t1239 VSSD.t1126 724.904
R8542 VSSD.t879 VSSD.t96 716.476
R8543 VSSD.t973 VSSD.t137 716.476
R8544 VSSD.t1700 VSSD.t394 716.476
R8545 VSSD.t455 VSSD.t451 716.476
R8546 VSSD.t744 VSSD.t704 716.476
R8547 VSSD.t641 VSSD.t416 708.047
R8548 VSSD.t736 VSSD.t1791 708.047
R8549 VSSD.t321 VSSD.t408 708.047
R8550 VSSD.t716 VSSD.t714 708.047
R8551 VSSD.t1712 VSSD.t899 708.047
R8552 VSSD.t204 VSSD.t961 708.047
R8553 VSSD.t528 VSSD.t598 708.047
R8554 VSSD.t8 VSSD.t982 708.047
R8555 VSSD.t919 VSSD.t144 708.047
R8556 VSSD.t565 VSSD.t380 708.047
R8557 VSSD.t380 VSSD.t420 708.047
R8558 VSSD.t420 VSSD.t1177 708.047
R8559 VSSD.t1177 VSSD.t1629 708.047
R8560 VSSD.t1010 VSSD.t546 708.047
R8561 VSSD.t546 VSSD.t1012 708.047
R8562 VSSD.t1709 VSSD.t646 708.047
R8563 VSSD.t602 VSSD.t520 708.047
R8564 VSSD.t1771 VSSD.t1769 708.047
R8565 VSSD.t1103 VSSD.t1099 708.047
R8566 VSSD.t1099 VSSD.t1101 708.047
R8567 VSSD.t756 VSSD.t1831 708.047
R8568 VSSD.t1831 VSSD.t758 708.047
R8569 VSSD.t1775 VSSD.t20 708.047
R8570 VSSD.t616 VSSD.t773 708.047
R8571 VSSD.t1839 VSSD.t4 708.047
R8572 VSSD.t1160 VSSD.t344 708.047
R8573 VSSD.t340 VSSD.t342 708.047
R8574 VSSD.t1081 VSSD.t1077 708.047
R8575 VSSD.t949 VSSD.t947 708.047
R8576 VSSD.t637 VSSD.t142 708.047
R8577 VSSD.t390 VSSD.t1585 708.047
R8578 VSSD.t1092 VSSD.t149 708.047
R8579 VSSD.t106 VSSD.t909 708.047
R8580 VSSD.t911 VSSD.t106 708.047
R8581 VSSD.t1834 VSSD.t78 708.047
R8582 VSSD.t83 VSSD.t85 708.047
R8583 VSSD.t575 VSSD.t464 708.047
R8584 VSSD.t777 VSSD.t1006 708.047
R8585 VSSD.t1621 VSSD.t1048 708.047
R8586 VSSD.t1843 VSSD.t75 708.047
R8587 VSSD.t1598 VSSD.t1600 708.047
R8588 VSSD.t1801 VSSD.t468 708.047
R8589 VSSD.t426 VSSD.t111 708.047
R8590 VSSD.t927 VSSD.t877 708.047
R8591 VSSD.t323 VSSD.t541 708.047
R8592 VSSD.t1638 VSSD.t1749 708.047
R8593 VSSD.t45 VSSD.t43 708.047
R8594 VSSD.t933 VSSD.t929 708.047
R8595 VSSD.t18 VSSD.t16 708.047
R8596 VSSD.t466 VSSD.t1578 708.047
R8597 VSSD.t297 VSSD.t459 708.047
R8598 VSSD.t1723 VSSD.t1693 708.047
R8599 VSSD.t1129 VSSD.t443 708.047
R8600 VSSD.t1820 VSSD.t1732 708.047
R8601 VSSD.t829 VSSD.t825 708.047
R8602 VSSD.t741 VSSD.t1618 708.047
R8603 VSSD.t354 VSSD.t356 708.047
R8604 VSSD.t1040 VSSD.t1046 708.047
R8605 VSSD.t52 VSSD.t1119 708.047
R8606 VSSD.t413 VSSD.t1002 708.047
R8607 VSSD.t56 VSSD.t327 708.047
R8608 VSSD.t632 VSSD.t54 708.047
R8609 VSSD.t691 VSSD.t693 708.047
R8610 VSSD.t586 VSSD.t538 708.047
R8611 VSSD.t1816 VSSD.t1814 708.047
R8612 VSSD.t518 VSSD.t731 708.047
R8613 VSSD.t600 VSSD.t1032 708.047
R8614 VSSD.t1760 VSSD.t584 708.047
R8615 VSSD.t72 VSSD.t782 708.047
R8616 VSSD.t302 VSSD.t678 699.617
R8617 VSSD.t24 VSSD.t1738 699.617
R8618 VSSD VSSD.t795 699.617
R8619 VSSD.t1110 VSSD.t62 699.617
R8620 VSSD.t1729 VSSD.t480 699.617
R8621 VSSD.t1787 VSSD.t482 699.617
R8622 VSSD VSSD.t679 691.188
R8623 VSSD.t1558 VSSD.t306 691.188
R8624 VSSD.t1147 VSSD.t197 691.188
R8625 VSSD.t728 VSSD.t975 691.188
R8626 VSSD.t869 VSSD.t1563 691.188
R8627 VSSD.t1381 VSSD.t123 691.188
R8628 VSSD.t895 VSSD.t834 691.188
R8629 VSSD.t665 VSSD.t213 691.188
R8630 VSSD.t1204 VSSD.t311 691.188
R8631 VSSD.t723 VSSD.t1485 682.76
R8632 VSSD.t588 VSSD.t1207 682.76
R8633 VSSD.t1096 VSSD.t140 674.331
R8634 VSSD.t621 VSSD.t206 674.331
R8635 VSSD.t913 VSSD.t1625 674.331
R8636 VSSD.t32 VSSD.t827 674.331
R8637 VSSD.t94 VSSD.t132 665.9
R8638 VSSD.t740 VSSD.t1153 665.9
R8639 VSSD.t1819 VSSD.t807 657.471
R8640 VSSD.t1785 VSSD.t799 657.471
R8641 VSSD.t1156 VSSD.t684 657.471
R8642 VSSD.t861 VSSD.t1128 657.471
R8643 VSSD.t1717 VSSD.t1091 657.471
R8644 VSSD.t412 VSSD.t368 657.471
R8645 VSSD.t985 VSSD.t1773 657.471
R8646 VSSD.t415 VSSD.t577 657.471
R8647 VSSD.t937 VSSD.t1774 657.471
R8648 VSSD.t762 VSSD.t796 649.043
R8649 VSSD.t977 VSSD.t510 649.043
R8650 VSSD.n2694 VSSD 649.043
R8651 VSSD.t571 VSSD.t232 649.043
R8652 VSSD.t69 VSSD.t619 640.614
R8653 VSSD.t1691 VSSD.t37 640.614
R8654 VSSD.t68 VSSD.t278 640.614
R8655 VSSD.t1124 VSSD.t835 640.614
R8656 VSSD VSSD.t1272 632.184
R8657 VSSD.n826 VSSD 632.184
R8658 VSSD.n827 VSSD 632.184
R8659 VSSD.n866 VSSD 632.184
R8660 VSSD.t1213 VSSD 632.184
R8661 VSSD VSSD.n1295 632.184
R8662 VSSD VSSD.t374 632.184
R8663 VSSD.t662 VSSD 632.184
R8664 VSSD.t646 VSSD 632.184
R8665 VSSD VSSD.n3303 632.184
R8666 VSSD.t1321 VSSD 632.184
R8667 VSSD VSSD.n1099 632.184
R8668 VSSD.n3055 VSSD 632.184
R8669 VSSD.t1422 VSSD 632.184
R8670 VSSD.t958 VSSD 632.184
R8671 VSSD.t1437 VSSD 632.184
R8672 VSSD.t1757 VSSD.t747 632.184
R8673 VSSD VSSD.n1481 632.184
R8674 VSSD.t1795 VSSD 632.184
R8675 VSSD.t1254 VSSD 632.184
R8676 VSSD.t535 VSSD.t1116 632.184
R8677 VSSD.n2107 VSSD 632.184
R8678 VSSD.n2140 VSSD 632.184
R8679 VSSD.t540 VSSD.t120 632.184
R8680 VSSD.t1263 VSSD 632.184
R8681 VSSD.n1657 VSSD 632.184
R8682 VSSD VSSD.t1462 632.184
R8683 VSSD.n171 VSSD 632.184
R8684 VSSD.n249 VSSD 632.184
R8685 VSSD.t1228 VSSD 632.184
R8686 VSSD.t1740 VSSD.t1760 632.184
R8687 VSSD VSSD.n3389 623.755
R8688 VSSD.t1289 VSSD 623.755
R8689 VSSD.t1167 VSSD 623.755
R8690 VSSD.n2861 VSSD 623.755
R8691 VSSD.t1647 VSSD.t1735 623.755
R8692 VSSD.n2566 VSSD 623.755
R8693 VSSD.t645 VSSD.t1711 623.755
R8694 VSSD VSSD.t588 623.755
R8695 VSSD.t441 VSSD 623.755
R8696 VSSD.n1970 VSSD 623.755
R8697 VSSD VSSD.t951 623.755
R8698 VSSD.t941 VSSD.t386 623.755
R8699 VSSD.n1616 VSSD 623.755
R8700 VSSD.t225 VSSD 623.755
R8701 VSSD VSSD.n490 623.755
R8702 VSSD.t856 VSSD.t303 623.755
R8703 VSSD.n671 VSSD 623.755
R8704 VSSD.t1307 VSSD 623.755
R8705 VSSD.n3668 VSSD 623.755
R8706 VSSD VSSD.n3667 623.755
R8707 VSSD.t1169 VSSD 623.755
R8708 VSSD.t1042 VSSD 615.327
R8709 VSSD.t813 VSSD 615.327
R8710 VSSD.t211 VSSD.t1124 615.327
R8711 VSSD.t779 VSSD.t508 606.898
R8712 VSSD.t47 VSSD 606.898
R8713 VSSD.n866 VSSD.t69 606.898
R8714 VSSD.t917 VSSD.t268 606.898
R8715 VSSD.t581 VSSD.t1141 606.898
R8716 VSSD.t1589 VSSD.t862 606.898
R8717 VSSD.t1652 VSSD.t1647 606.898
R8718 VSSD.t250 VSSD.t335 606.898
R8719 VSSD.t227 VSSD.t514 606.898
R8720 VSSD.t497 VSSD.t1796 606.898
R8721 VSSD.t164 VSSD.t645 606.898
R8722 VSSD.t347 VSSD.t977 606.898
R8723 VSSD.t760 VSSD.t1785 606.898
R8724 VSSD.t392 VSSD.t726 606.898
R8725 VSSD.t121 VSSD.t1131 606.898
R8726 VSSD.t1799 VSSD.t1810 606.898
R8727 VSSD.t219 VSSD.t442 606.898
R8728 VSSD.t499 VSSD.t271 606.898
R8729 VSSD.t761 VSSD.t1676 606.898
R8730 VSSD.t1699 VSSD.t891 606.898
R8731 VSSD.t607 VSSD.t1499 606.898
R8732 VSSD.t1686 VSSD.t613 606.898
R8733 VSSD.t51 VSSD.t234 606.898
R8734 VSSD.t453 VSSD.t571 606.898
R8735 VSSD.t1089 VSSD.t258 606.898
R8736 VSSD.t935 VSSD.t236 606.898
R8737 VSSD.t979 VSSD.t240 606.898
R8738 VSSD.t303 VSSD.t248 606.898
R8739 VSSD.t262 VSSD.t635 606.898
R8740 VSSD.t953 VSSD.t1658 606.898
R8741 VSSD.t493 VSSD.t1127 606.898
R8742 VSSD.t512 VSSD.t1646 606.898
R8743 VSSD.n671 VSSD.n670 599.125
R8744 VSSD.n3669 VSSD.n3668 599.125
R8745 VSSD.t873 VSSD.t575 598.467
R8746 VSSD.t325 VSSD.t1801 598.467
R8747 VSSD.t1749 VSSD.t765 598.467
R8748 VSSD.t967 VSSD.t267 590.038
R8749 VSSD.t98 VSSD.t1581 590.038
R8750 VSSD.t702 VSSD 590.038
R8751 VSSD.t35 VSSD.t470 590.038
R8752 VSSD.n248 VSSD.t634 590.038
R8753 VSSD.t1781 VSSD.t621 581.61
R8754 VSSD.t1064 VSSD.t864 581.61
R8755 VSSD VSSD.t927 581.61
R8756 VSSD.t541 VSSD 581.61
R8757 VSSD.t1496 VSSD.t1793 573.181
R8758 VSSD.t567 VSSD.t1052 573.181
R8759 VSSD.t1073 VSSD.t1143 573.181
R8760 VSSD.t596 VSSD.t360 573.181
R8761 VSSD.t1069 VSSD.t643 573.181
R8762 VSSD.t1075 VSSD.t358 573.181
R8763 VSSD.t1071 VSSD.t803 573.181
R8764 VSSD.t350 VSSD.t797 573.181
R8765 VSSD.t1615 VSSD.t1135 573.181
R8766 VSSD.t841 VSSD.t1038 573.181
R8767 VSSD.t517 VSSD.t1428 573.181
R8768 VSSD.t1813 VSSD 564.751
R8769 VSSD.n3665 VSSD 564.751
R8770 VSSD.t1707 VSSD.t1066 564.751
R8771 VSSD.t648 VSSD.t689 564.751
R8772 VSSD.n3664 VSSD 564.751
R8773 VSSD.n3663 VSSD 564.751
R8774 VSSD.t801 VSSD.t333 564.751
R8775 VSSD.n3662 VSSD 564.751
R8776 VSSD.t2 VSSD 564.751
R8777 VSSD.n3661 VSSD 564.751
R8778 VSSD.n3660 VSSD 564.751
R8779 VSSD.n3659 VSSD 564.751
R8780 VSSD.n3658 VSSD 564.751
R8781 VSSD VSSD.n3666 564.751
R8782 VSSD.t527 VSSD.t851 556.322
R8783 VSSD VSSD.t428 556.322
R8784 VSSD.t1387 VSSD.t488 556.322
R8785 VSSD.t1650 VSSD.t1850 556.322
R8786 VSSD.t1134 VSSD.t631 556.322
R8787 VSSD VSSD.t786 547.894
R8788 VSSD VSSD.t784 547.894
R8789 VSSD VSSD.t382 547.894
R8790 VSSD.t936 VSSD.t666 547.894
R8791 VSSD.t598 VSSD 547.894
R8792 VSSD.t144 VSSD 547.894
R8793 VSSD.t147 VSSD 547.894
R8794 VSSD.t1836 VSSD 547.894
R8795 VSSD VSSD.t1162 547.894
R8796 VSSD.t464 VSSD 547.894
R8797 VSSD.t1006 VSSD 547.894
R8798 VSSD.t388 VSSD 547.894
R8799 VSSD.t1275 VSSD.t1825 547.894
R8800 VSSD.t815 VSSD 547.894
R8801 VSSD.t468 VSSD 547.894
R8802 VSSD.t1004 VSSD 547.894
R8803 VSSD VSSD.t426 547.894
R8804 VSSD.t406 VSSD 547.894
R8805 VSSD VSSD.t466 547.894
R8806 VSSD VSSD.t1129 547.894
R8807 VSSD VSSD.t32 547.894
R8808 VSSD VSSD.t58 547.894
R8809 VSSD VSSD.t56 547.894
R8810 VSSD VSSD.t939 547.894
R8811 VSSD.t954 VSSD.t1440 547.894
R8812 VSSD.t731 VSSD 547.894
R8813 VSSD.t780 VSSD 547.894
R8814 VSSD.t408 VSSD.t779 539.465
R8815 VSSD.t96 VSSD.t567 539.465
R8816 VSSD VSSD.t687 539.465
R8817 VSSD.t1019 VSSD.t845 539.465
R8818 VSSD.t1158 VSSD.t847 539.465
R8819 VSSD.t754 VSSD.t180 539.465
R8820 VSSD.t1135 VSSD.t219 539.465
R8821 VSSD.t271 VSSD.t841 539.465
R8822 VSSD.t110 VSSD.t1155 539.465
R8823 VSSD.t434 VSSD.t202 539.465
R8824 VSSD.t92 VSSD.t1186 531.034
R8825 VSSD.t87 VSSD.t1056 531.034
R8826 VSSD.t215 VSSD.t1157 531.034
R8827 VSSD VSSD.t1390 531.034
R8828 VSSD.t269 VSSD 522.606
R8829 VSSD.t956 VSSD 522.606
R8830 VSSD.t544 VSSD.t433 522.606
R8831 VSSD.t1164 VSSD.t994 522.606
R8832 VSSD VSSD.t204 514.177
R8833 VSSD.t1783 VSSD.t1122 514.177
R8834 VSSD.t1402 VSSD 514.177
R8835 VSSD VSSD.t1827 514.177
R8836 VSSD VSSD.t1583 514.177
R8837 VSSD.t552 VSSD.t683 514.177
R8838 VSSD.t273 VSSD.t1803 514.177
R8839 VSSD.t284 VSSD 514.177
R8840 VSSD.t1608 VSSD.t921 514.177
R8841 VSSD.t1024 VSSD.t1604 514.177
R8842 VSSD.t1751 VSSD.t209 514.177
R8843 VSSD VSSD.t18 514.177
R8844 VSSD VSSD.t502 514.177
R8845 VSSD.t1048 VSSD.t761 505.748
R8846 VSSD.t282 VSSD.t925 505.748
R8847 VSSD.t714 VSSD.t47 497.318
R8848 VSSD.t660 VSSD 497.318
R8849 VSSD.t893 VSSD.t1688 497.318
R8850 VSSD.t969 VSSD.t1695 488.889
R8851 VSSD.t699 VSSD.t291 488.889
R8852 VSSD.t589 VSSD.t153 488.889
R8853 VSSD.t1114 VSSD 488.889
R8854 VSSD.t1105 VSSD.t706 488.889
R8855 VSSD.t872 VSSD.t1068 488.889
R8856 VSSD VSSD.t1094 480.461
R8857 VSSD.t65 VSSD.t1451 480.461
R8858 VSSD.t697 VSSD 480.461
R8859 VSSD.t252 VSSD.t6 480.461
R8860 VSSD.t166 VSSD.t1079 480.461
R8861 VSSD.t1702 VSSD 480.461
R8862 VSSD VSSD.t160 480.461
R8863 VSSD.t352 VSSD.t238 480.461
R8864 VSSD VSSD.t1766 480.461
R8865 VSSD.t943 VSSD 480.461
R8866 VSSD.t168 VSSD.t384 472.031
R8867 VSSD.t382 VSSD.t491 472.031
R8868 VSSD VSSD.t1014 472.031
R8869 VSSD VSSD.t1036 472.031
R8870 VSSD.n3056 VSSD.t1839 472.031
R8871 VSSD.t623 VSSD 472.031
R8872 VSSD.t1008 VSSD.t439 472.031
R8873 VSSD.n1481 VSSD.t887 472.031
R8874 VSSD.n1970 VSSD.t1050 472.031
R8875 VSSD.t378 VSSD.t295 472.031
R8876 VSSD.t931 VSSD.t438 472.031
R8877 VSSD.t232 VSSD 472.031
R8878 VSSD.t364 VSSD 472.031
R8879 VSSD.n490 VSSD.t356 472.031
R8880 VSSD.t738 VSSD.t843 463.603
R8881 VSSD VSSD.t863 463.603
R8882 VSSD VSSD.t594 463.603
R8883 VSSD.t1572 VSSD.t135 463.603
R8884 VSSD.t317 VSSD.t554 463.603
R8885 VSSD.t799 VSSD.t60 455.173
R8886 VSSD.t228 VSSD.t1758 455.173
R8887 VSSD.t887 VSSD 455.173
R8888 VSSD.t1050 VSSD 455.173
R8889 VSSD.t1662 VSSD.t159 455.173
R8890 VSSD.t119 VSSD.t1684 455.173
R8891 VSSD.t1664 VSSD 455.173
R8892 VSSD.t745 VSSD.t477 455.173
R8893 VSSD.t707 VSSD.t859 455.173
R8894 VSSD VSSD.t536 455.173
R8895 VSSD VSSD.t1054 455.173
R8896 VSSD.t1574 VSSD.t192 446.743
R8897 VSSD.t1841 VSSD 446.743
R8898 VSSD.t113 VSSD.t1602 446.743
R8899 VSSD.t1580 VSSD 446.743
R8900 VSSD VSSD.t198 446.743
R8901 VSSD VSSD.t500 446.743
R8902 VSSD VSSD.t1028 438.315
R8903 VSSD.t1451 VSSD.t664 438.315
R8904 VSSD VSSD.t65 438.315
R8905 VSSD.t1470 VSSD.t697 438.315
R8906 VSSD.t104 VSSD.t629 438.315
R8907 VSSD.t909 VSSD.t1743 438.315
R8908 VSSD.t217 VSSD.t1808 438.315
R8909 VSSD.t708 VSSD 438.315
R8910 VSSD.t1668 VSSD.t1016 438.315
R8911 VSSD.t551 VSSD 438.315
R8912 VSSD.t1151 VSSD.t223 438.315
R8913 VSSD.t770 VSSD.t625 438.315
R8914 VSSD.t1737 VSSD 438.315
R8915 VSSD.t1845 VSSD.t866 429.885
R8916 VSSD.t1804 VSSD.t720 429.885
R8917 VSSD.t1642 VSSD.t652 429.885
R8918 VSSD.t457 VSSD.t1000 429.885
R8919 VSSD.t14 VSSD.t618 429.885
R8920 VSSD.n2106 VSSD.t280 421.457
R8921 VSSD.t834 VSSD.t734 421.457
R8922 VSSD.t418 VSSD.t665 421.457
R8923 VSSD.t1179 VSSD.t376 413.027
R8924 VSSD.t151 VSSD.t1087 413.027
R8925 VSSD.t560 VSSD.t24 413.027
R8926 VSSD VSSD.t14 413.027
R8927 VSSD.t208 VSSD 413.027
R8928 VSSD.t480 VSSD.t1097 413.027
R8929 VSSD.t1610 VSSD.t1787 413.027
R8930 VSSD.t1727 VSSD.t736 404.599
R8931 VSSD.n3304 VSSD.t654 404.599
R8932 VSSD.n1482 VSSD.t791 404.599
R8933 VSSD.t709 VSSD.t1725 404.599
R8934 VSSD.t1725 VSSD.t3 404.599
R8935 VSSD.t3 VSSD.t101 404.599
R8936 VSSD.n2455 VSSD.t1044 404.599
R8937 VSSD.t1025 VSSD.t573 404.599
R8938 VSSD.t445 VSSD.t1025 404.599
R8939 VSSD.t1791 VSSD 396.17
R8940 VSSD.t10 VSSD 396.17
R8941 VSSD.t1633 VSSD.t461 396.17
R8942 VSSD.t394 VSSD.t217 396.17
R8943 VSSD.t336 VSSD.t709 396.17
R8944 VSSD.t101 VSSD.t857 396.17
R8945 VSSD.t451 VSSD.t1668 396.17
R8946 VSSD.t223 VSSD.t744 396.17
R8947 VSSD VSSD.t319 396.17
R8948 VSSD.n1295 VSSD.t1327 387.74
R8949 VSSD.t1745 VSSD.t151 387.74
R8950 VSSD.n672 VSSD.t1340 387.74
R8951 VSSD VSSD.t988 379.31
R8952 VSSD VSSD.t10 379.31
R8953 VSSD.t866 VSSD.t66 379.31
R8954 VSSD.t1030 VSSD.t1804 379.31
R8955 VSSD.t1627 VSSD.t28 379.31
R8956 VSSD.t734 VSSD.t745 379.31
R8957 VSSD.t859 VSSD.t418 379.31
R8958 VSSD.t12 VSSD.t721 370.882
R8959 VSSD.t720 VSSD.t1845 370.882
R8960 VSSD.t1846 VSSD.t952 370.882
R8961 VSSD.t430 VSSD.t936 370.882
R8962 VSSD.t39 VSSD.t1699 370.882
R8963 VSSD.t1636 VSSD.n2454 370.882
R8964 VSSD VSSD.t208 370.882
R8965 VSSD.n2140 VSSD.t406 370.882
R8966 VSSD.n1617 VSSD.t200 370.882
R8967 VSSD VSSD.t1566 364.712
R8968 VSSD.t907 VSSD.t1631 362.452
R8969 VSSD.t1631 VSSD.t905 362.452
R8970 VSSD.t923 VSSD.t486 362.452
R8971 VSSD.t1602 VSSD.t923 362.452
R8972 VSSD VSSD.t1807 362.452
R8973 VSSD VSSD.t708 354.024
R8974 VSSD.n1528 VSSD.n1513 352
R8975 VSSD.t905 VSSD.t1627 345.594
R8976 VSSD.t194 VSSD 337.166
R8977 VSSD.t700 VSSD.t250 337.166
R8978 VSSD.t1789 VSSD.t497 337.166
R8979 VSSD.n2454 VSSD.t702 337.166
R8980 VSSD.t240 VSSD.t1718 337.166
R8981 VSSD.t889 VSSD.t563 337.166
R8982 VSSD.n3398 VSSD.t1266 332.212
R8983 VSSD.n96 VSSD.t1324 332.212
R8984 VSSD.n73 VSSD.t1313 332.212
R8985 VSSD.t28 VSSD.t1633 328.736
R8986 VSSD.t1833 VSSD 328.736
R8987 VSSD VSSD.t1081 328.736
R8988 VSSD VSSD.t729 328.736
R8989 VSSD VSSD.t1174 328.736
R8990 VSSD.t1054 VSSD 328.736
R8991 VSSD VSSD.t1060 320.307
R8992 VSSD.n3304 VSSD.t823 320.307
R8993 VSSD.t153 VSSD.t1745 320.307
R8994 VSSD.t793 VSSD 320.307
R8995 VSSD.t1176 VSSD.t1527 320.307
R8996 VSSD.t1337 VSSD.t1692 320.307
R8997 VSSD VSSD.t1664 320.307
R8998 VSSD.t461 VSSD.t1179 311.877
R8999 VSSD.t1036 VSSD 311.877
R9000 VSSD.t763 VSSD.t969 311.877
R9001 VSSD.t291 VSSD.t650 311.877
R9002 VSSD.t22 VSSD.t560 311.877
R9003 VSSD VSSD.t364 311.877
R9004 VSSD VSSD.t80 311.877
R9005 VSSD.t379 VSSD 311.877
R9006 VSSD.n968 VSSD.t1805 307.536
R9007 VSSD.n974 VSSD.t867 307.536
R9008 VSSD.n815 VSSD.t531 307.536
R9009 VSSD.n3342 VSSD.t844 307.536
R9010 VSSD.n881 VSSD.t1123 307.536
R9011 VSSD.n1199 VSSD.t902 307.536
R9012 VSSD.n1199 VSSD.t1133 307.536
R9013 VSSD.n1094 VSSD.t764 307.536
R9014 VSSD.n3036 VSSD.t1084 307.536
R9015 VSSD.n3035 VSSD.t339 307.536
R9016 VSSD.n3063 VSSD.t752 307.536
R9017 VSSD.n3063 VSSD.t1009 307.536
R9018 VSSD.n2536 VSSD.t109 307.536
R9019 VSSD.n2616 VSSD.t840 307.536
R9020 VSSD.n2820 VSSD.t624 307.536
R9021 VSSD.n2810 VSSD.t1088 307.536
R9022 VSSD.n1396 VSSD.t858 307.536
R9023 VSSD.n2488 VSSD.t337 307.536
R9024 VSSD.n1535 VSSD.t916 307.536
R9025 VSSD.n1461 VSSD.t1641 307.536
R9026 VSSD.n2255 VSSD.t1824 307.536
R9027 VSSD.n2204 VSSD.t367 307.536
R9028 VSSD.n1686 VSSD.t860 307.536
R9029 VSSD.n1810 VSSD.t746 307.536
R9030 VSSD.n1861 VSSD.t363 307.536
R9031 VSSD.n448 VSSD.t628 307.536
R9032 VSSD.n160 VSSD.t31 307.536
R9033 VSSD.n3724 VSSD.t1741 307.536
R9034 VSSD.n883 VSSD.t437 306.988
R9035 VSSD.n1639 VSSD.t365 306.988
R9036 VSSD.n3008 VSSD.t651 306.983
R9037 VSSD.n707 VSSD.t71 304.238
R9038 VSSD.n778 VSSD.t130 304.238
R9039 VSSD.n3295 VSSD.t526 304.238
R9040 VSSD.n2928 VSSD.t1037 304.238
R9041 VSSD.n2760 VSSD.t1706 304.238
R9042 VSSD.n2326 VSSD.t1826 304.238
R9043 VSSD.n2338 VSSD.t668 304.238
R9044 VSSD.n1509 VSSD.t874 304.238
R9045 VSSD.n2388 VSSD.t1086 304.238
R9046 VSSD.n2014 VSSD.t326 304.238
R9047 VSSD.n2072 VSSD.t1722 304.238
R9048 VSSD.n2108 VSSD.t1109 304.238
R9049 VSSD.n2206 VSSD.t766 304.238
R9050 VSSD.n1700 VSSD.t1107 304.238
R9051 VSSD.n1915 VSSD.t1624 304.238
R9052 VSSD.n185 VSSD.t713 304.238
R9053 VSSD.n198 VSSD.t425 304.238
R9054 VSSD.n370 VSSD.t955 304.238
R9055 VSSD.n356 VSSD.t1111 304.238
R9056 VSSD.n3678 VSSD.t174 304.238
R9057 VSSD.n9 VSSD.t818 304.238
R9058 VSSD.t673 VSSD.t1727 303.449
R9059 VSSD.t185 VSSD.t673 303.449
R9060 VSSD.t448 VSSD.n827 303.449
R9061 VSSD.t436 VSSD 303.449
R9062 VSSD.t1014 VSSD 303.449
R9063 VSSD.n1482 VSSD.t793 303.449
R9064 VSSD.t1810 VSSD.t317 303.449
R9065 VSSD.n2455 VSSD.t1042 303.449
R9066 VSSD.t1606 VSSD.n2106 303.449
R9067 VSSD.t635 VSSD.t117 303.449
R9068 VSSD.t1753 VSSD.t953 303.449
R9069 VSSD.n3667 VSSD.t1169 303.449
R9070 VSSD.t1364 VSSD 301.519
R9071 VSSD.t376 VSSD.t1642 295.019
R9072 VSSD VSSD.t1617 295.019
R9073 VSSD.t428 VSSD.t457 295.019
R9074 VSSD.t1087 VSSD.t911 295.019
R9075 VSSD.t1742 VSSD 295.019
R9076 VSSD VSSD.t77 295.019
R9077 VSSD.t439 VSSD.t552 295.019
R9078 VSSD VSSD.t777 295.019
R9079 VSSD.t295 VSSD.t273 295.019
R9080 VSSD VSSD.t1114 295.019
R9081 VSSD.t618 VSSD.t22 295.019
R9082 VSSD.t160 VSSD 295.019
R9083 VSSD.t209 VSSD.t931 295.019
R9084 VSSD VSSD.t964 295.019
R9085 VSSD VSSD.t1614 295.019
R9086 VSSD.t810 VSSD.t1783 286.591
R9087 VSSD VSSD.t450 286.591
R9088 VSSD.t1527 VSSD.t1680 286.591
R9089 VSSD.t242 VSSD.t1337 286.591
R9090 VSSD.t1034 VSSD.t544 286.591
R9091 VSSD.t994 VSSD.t998 286.591
R9092 VSSD.n3213 VSSD.t647 286.433
R9093 VSSD.n3206 VSSD.t1708 285.481
R9094 VSSD.n3184 VSSD.t688 284.067
R9095 VSSD.n3212 VSSD.t690 284.024
R9096 VSSD VSSD.t1612 278.161
R9097 VSSD.t1827 VSSD 278.161
R9098 VSSD.t188 VSSD.t1574 278.161
R9099 VSSD.t891 VSSD.t221 278.161
R9100 VSSD.t278 VSSD.t113 278.161
R9101 VSSD.t809 VSSD.t762 269.733
R9102 VSSD VSSD.t907 269.733
R9103 VSSD.t1000 VSSD 269.733
R9104 VSSD.t60 VSSD.t801 269.733
R9105 VSSD.t1743 VSSD.t104 269.733
R9106 VSSD.t516 VSSD.t413 269.733
R9107 VSSD.t327 VSSD.t963 269.733
R9108 VSSD.t563 VSSD.t770 269.733
R9109 VSSD.t155 VSSD.t893 269.733
R9110 VSSD.n674 VSSD.t1971 266.474
R9111 VSSD.n1148 VSSD.t1975 266.474
R9112 VSSD.n2287 VSSD.t1865 266.474
R9113 VSSD.n3247 VSSD.t1891 265.317
R9114 VSSD.n2712 VSSD.t1917 265.317
R9115 VSSD.n1711 VSSD.t1974 265.317
R9116 VSSD.n567 VSSD.t1863 265.055
R9117 VSSD.n561 VSSD.t1889 262.784
R9118 VSSD.n562 VSSD.t1893 262.784
R9119 VSSD.n554 VSSD.t1978 262.784
R9120 VSSD.n887 VSSD.t1902 262.784
R9121 VSSD.n888 VSSD.t1943 262.784
R9122 VSSD.n492 VSSD.t1950 262.784
R9123 VSSD.n494 VSSD.t1857 262.784
R9124 VSSD.n1228 VSSD.t1866 262.784
R9125 VSSD.n1140 VSSD.t1915 262.784
R9126 VSSD.n1142 VSSD.t1874 262.784
R9127 VSSD.n3251 VSSD.t1864 262.784
R9128 VSSD.n3252 VSSD.t1941 262.784
R9129 VSSD.n2863 VSSD.t1934 262.784
R9130 VSSD.n2864 VSSD.t1936 262.784
R9131 VSSD.n3077 VSSD.t1862 262.784
R9132 VSSD.n3078 VSSD.t1869 262.784
R9133 VSSD.n2559 VSSD.t1884 262.784
R9134 VSSD.n2561 VSSD.t1897 262.784
R9135 VSSD.n2716 VSSD.t1954 262.784
R9136 VSSD.n2717 VSSD.t1970 262.784
R9137 VSSD.n1483 VSSD.t1886 262.784
R9138 VSSD.n1484 VSSD.t1898 262.784
R9139 VSSD.n2403 VSSD.t1959 262.784
R9140 VSSD.n2404 VSSD.t1973 262.784
R9141 VSSD.n1964 VSSD.t1987 262.784
R9142 VSSD.n1965 VSSD.t1855 262.784
R9143 VSSD.n1441 VSSD.t1986 262.784
R9144 VSSD.n2165 VSSD.t1921 262.784
R9145 VSSD.n2166 VSSD.t1922 262.784
R9146 VSSD.n1715 VSSD.t1878 262.784
R9147 VSSD.n1717 VSSD.t1883 262.784
R9148 VSSD.n1600 VSSD.t1946 262.784
R9149 VSSD.n1601 VSSD.t1948 262.784
R9150 VSSD.n267 VSSD.t1980 262.784
R9151 VSSD.n268 VSSD.t1984 262.784
R9152 VSSD.n134 VSSD.t1907 262.784
R9153 VSSD.n135 VSSD.t1912 262.784
R9154 VSSD.n3788 VSSD.t1977 262.784
R9155 VSSD.n3789 VSSD.t1982 262.784
R9156 VSSD.n717 VSSD.t1963 262.719
R9157 VSSD.n687 VSSD.t1881 262.719
R9158 VSSD.n641 VSSD.t1942 262.719
R9159 VSSD.n630 VSSD.t1923 262.719
R9160 VSSD.n619 VSSD.t1958 262.719
R9161 VSSD.n943 VSSD.t1858 262.719
R9162 VSSD.n3363 VSSD.t1972 262.719
R9163 VSSD.n3238 VSSD.t1877 262.719
R9164 VSSD.n1117 VSSD.t1885 262.719
R9165 VSSD.n1369 VSSD.t1856 262.719
R9166 VSSD.n2703 VSSD.t1900 262.719
R9167 VSSD.n2392 VSSD.t1894 262.719
R9168 VSSD.n2413 VSSD.t1905 262.719
R9169 VSSD.n1750 VSSD.t1960 262.719
R9170 VSSD.n1926 VSSD.t1930 262.719
R9171 VSSD.n1904 VSSD.t1867 262.719
R9172 VSSD.n116 VSSD.t1852 262.719
R9173 VSSD.n109 VSSD.t1927 262.719
R9174 VSSD.n88 VSSD.t1870 262.719
R9175 VSSD.n75 VSSD.t1880 262.719
R9176 VSSD.n65 VSSD.t1964 262.719
R9177 VSSD.n49 VSSD.t1875 262.719
R9178 VSSD.n3597 VSSD.t1876 262.719
R9179 VSSD.n3604 VSSD.t1888 262.719
R9180 VSSD.n318 VSSD.t1911 262.719
R9181 VSSD.n257 VSSD.t1920 262.719
R9182 VSSD.n257 VSSD.t1913 262.719
R9183 VSSD.n264 VSSD.t1933 262.719
R9184 VSSD.n264 VSSD.t1928 262.719
R9185 VSSD.n3751 VSSD.t1853 262.719
R9186 VSSD.n2 VSSD.t1931 262.719
R9187 VSSD.t384 VSSD 261.303
R9188 VSSD VSSD.t602 261.303
R9189 VSSD VSSD.t710 261.303
R9190 VSSD.t1583 VSSD 261.303
R9191 VSSD VSSD.t1160 261.303
R9192 VSSD.t192 VSSD.t1572 261.303
R9193 VSSD.t629 VSSD 261.303
R9194 VSSD VSSD.t1834 261.303
R9195 VSSD VSSD.t422 261.303
R9196 VSSD VSSD.t956 261.303
R9197 VSSD VSSD.t1636 261.303
R9198 VSSD.t877 VSSD 261.303
R9199 VSSD.t875 VSSD 261.303
R9200 VSSD VSSD.t1638 261.303
R9201 VSSD.t200 VSSD 261.303
R9202 VSSD.t258 VSSD.t362 261.303
R9203 VSSD.t1625 VSSD 261.303
R9204 VSSD VSSD.t741 261.303
R9205 VSSD.t502 VSSD 261.303
R9206 VSSD.t1002 VSSD 261.303
R9207 VSSD.t122 VSSD.t985 261.303
R9208 VSSD.t577 VSSD.t984 261.303
R9209 VSSD.t625 VSSD 261.303
R9210 VSSD.n982 VSSD.t1932 259.082
R9211 VSSD.n802 VSSD.t1940 259.082
R9212 VSSD.n1297 VSSD.t1860 259.082
R9213 VSSD.n3014 VSSD.t1879 259.082
R9214 VSSD.n1653 VSSD.t1896 259.082
R9215 VSSD.n3401 VSSD.t1872 259.082
R9216 VSSD.n3411 VSSD.t1976 259.082
R9217 VSSD.n3476 VSSD.t1957 259.082
R9218 VSSD.n3537 VSSD.t1961 259.082
R9219 VSSD.n3610 VSSD.t1939 259.082
R9220 VSSD.n3768 VSSD.t1861 259.082
R9221 VSSD VSSD.t1103 252.875
R9222 VSSD.t1585 VSSD 252.875
R9223 VSSD VSSD.t883 252.875
R9224 VSSD VSSD.t685 252.875
R9225 VSSD.t631 VSSD.t740 252.875
R9226 VSSD.t695 VSSD.t1134 252.875
R9227 VSSD VSSD.t600 252.875
R9228 VSSD.n2690 VSSD.t1001 244.853
R9229 VSSD.t851 VSSD.t436 244.445
R9230 VSSD VSSD.t1537 244.445
R9231 VSSD VSSD.t1292 244.445
R9232 VSSD.t554 VSSD.t458 244.445
R9233 VSSD.t1519 VSSD 244.445
R9234 VSSD.t1198 VSSD 244.445
R9235 VSSD.t1225 VSSD 244.445
R9236 VSSD.t1490 VSSD 244.445
R9237 VSSD.t1473 VSSD 244.445
R9238 VSSD.t1434 VSSD 244.445
R9239 VSSD.t1340 VSSD 244.445
R9240 VSSD.n2667 VSSD.t351 243.495
R9241 VSSD.n2684 VSSD.t1144 240.948
R9242 VSSD.n2078 VSSD.t15 240.948
R9243 VSSD.n3164 VSSD.t657 240.757
R9244 VSSD.n1326 VSSD.t800 238.44
R9245 VSSD.n2024 VSSD.t608 238.44
R9246 VSSD.n999 VSSD.t715 238.083
R9247 VSSD.n752 VSSD.t409 238.083
R9248 VSSD.n932 VSSD.t620 238.083
R9249 VSSD.n1138 VSSD.t9 238.083
R9250 VSSD.n1138 VSSD.t1822 238.083
R9251 VSSD.n2966 VSSD.t970 238.083
R9252 VSSD.n3007 VSSD.t292 238.083
R9253 VSSD.n3118 VSSD.t617 238.083
R9254 VSSD.n3081 VSSD.t343 238.083
R9255 VSSD.n3081 VSSD.t769 238.083
R9256 VSSD.n2583 VSSD.t950 238.083
R9257 VSSD.n1480 VSSD.t794 238.083
R9258 VSSD.n1416 VSSD.t1043 238.083
R9259 VSSD.n1417 VSSD.t814 238.083
R9260 VSSD.n2236 VSSD.t838 238.083
R9261 VSSD.n1883 VSSD.t572 238.083
R9262 VSSD.n487 VSSD.t1047 238.083
R9263 VSSD.n226 VSSD.t692 238.083
R9264 VSSD.n3683 VSSD.t545 238.083
R9265 VSSD.n19 VSSD.t995 238.083
R9266 VSSD.n3723 VSSD.t1761 238.083
R9267 VSSD.n1239 VSSD.t908 237.381
R9268 VSSD.n2211 VSSD.t403 237.029
R9269 VSSD.n375 VSSD.t1748 237.029
R9270 VSSD.n2582 VSSD.t1082 236.26
R9271 VSSD.t1414 VSSD.t195 236.016
R9272 VSSD.t721 VSSD.t168 236.016
R9273 VSSD.t491 VSSD.t1846 236.016
R9274 VSSD.t1052 VSSD.t430 236.016
R9275 VSSD VSSD.t1542 236.016
R9276 VSSD.t687 VSSD 236.016
R9277 VSSD.t310 VSSD.t87 236.016
R9278 VSSD.t1157 VSSD.t463 236.016
R9279 VSSD.t782 VSSD.t379 236.016
R9280 VSSD.n679 VSSD.t1817 233.732
R9281 VSSD.n864 VSSD.t962 233.732
R9282 VSSD.n942 VSSD.t1713 233.732
R9283 VSSD.n521 VSSD.t737 233.732
R9284 VSSD.n514 VSSD.t417 233.732
R9285 VSSD.n3265 VSSD.t307 233.732
R9286 VSSD.n2896 VSSD.t1772 233.732
R9287 VSSD.n3117 VSSD.t1840 233.732
R9288 VSSD.n2662 VSSD.t1573 233.732
R9289 VSSD.n2776 VSSD.t870 233.732
R9290 VSSD.n2730 VSSD.t124 233.732
R9291 VSSD.n2367 VSSD.t38 233.732
R9292 VSSD.n1491 VSSD.t84 233.732
R9293 VSSD.n1384 VSSD.t888 233.732
R9294 VSSD.n2419 VSSD.t76 233.732
R9295 VSSD.n1962 VSSD.t1599 233.732
R9296 VSSD.n1963 VSSD.t1051 233.732
R9297 VSSD.n2048 VSSD.t926 233.732
R9298 VSSD.n2179 VSSD.t44 233.732
R9299 VSSD.n2162 VSSD.t930 233.732
R9300 VSSD.n1729 VSSD.t312 233.732
R9301 VSSD.n1692 VSSD.t830 233.732
R9302 VSSD.n1660 VSSD.t1733 233.732
R9303 VSSD.n1611 VSSD.t17 233.732
R9304 VSSD.n1618 VSSD.t199 233.732
R9305 VSSD.n180 VSSD.t501 233.732
R9306 VSSD.n324 VSSD.t587 233.732
R9307 VSSD.n488 VSSD.t357 233.732
R9308 VSSD.t129 VSSD.t1496 227.587
R9309 VSSD.t784 VSSD 227.587
R9310 VSSD VSSD.t654 227.587
R9311 VSSD VSSD.t147 227.587
R9312 VSSD VSSD.t1836 227.587
R9313 VSSD VSSD.t1044 227.587
R9314 VSSD VSSD.t1686 227.587
R9315 VSSD.t58 VSSD 227.587
R9316 VSSD.t939 VSSD 227.587
R9317 VSSD.t1428 VSSD.t70 227.587
R9318 VSSD VSSD.t780 227.587
R9319 VSSD.n820 VSSD.t322 226.882
R9320 VSSD.n3351 VSSD.t674 226.882
R9321 VSSD.n1304 VSSD.t1645 226.882
R9322 VSSD.n1304 VSSD.t983 226.882
R9323 VSSD.n2968 VSSD.t968 226.882
R9324 VSSD.n2995 VSSD.t1582 226.882
R9325 VSSD.n3120 VSSD.t774 226.882
R9326 VSSD.n3119 VSSD.t5 226.882
R9327 VSSD.n3075 VSSD.t341 226.882
R9328 VSSD.n3075 VSSD.t768 226.882
R9329 VSSD.n2545 VSSD.t1078 226.882
R9330 VSSD.n2587 VSSD.t948 226.882
R9331 VSSD.n2365 VSSD.t534 226.882
R9332 VSSD.n2507 VSSD.t884 226.882
R9333 VSSD.n1496 VSSD.t86 226.882
R9334 VSSD.n1980 VSSD.t1601 226.882
R9335 VSSD.n2124 VSSD.t387 226.882
R9336 VSSD.n2159 VSSD.t46 226.882
R9337 VSSD.n1879 VSSD.t460 226.882
R9338 VSSD.n483 VSSD.t1041 226.882
R9339 VSSD.n140 VSSD.t355 226.882
R9340 VSSD.n181 VSSD.t503 226.882
R9341 VSSD.n209 VSSD.t940 226.882
R9342 VSSD.n343 VSSD.t694 226.882
R9343 VSSD.n37 VSSD.t128 226.882
R9344 VSSD.n3718 VSSD.t993 226.882
R9345 VSSD.n3725 VSSD.t585 226.882
R9346 VSSD.n1415 VSSD.t1045 224.643
R9347 VSSD.n746 VSSD.t717 223.748
R9348 VSSD.n680 VSSD.t1815 223.315
R9349 VSSD.n935 VSSD.t205 223.315
R9350 VSSD.n863 VSSD.t900 223.315
R9351 VSSD.n3370 VSSD.t642 223.315
R9352 VSSD.n872 VSSD.t622 223.315
R9353 VSSD.n3267 VSSD.t305 223.315
R9354 VSSD.n1126 VSSD.t1770 223.315
R9355 VSSD.n2659 VSSD.t1575 223.315
R9356 VSSD.n2778 VSSD.t1763 223.315
R9357 VSSD.n2732 VSSD.t1173 223.315
R9358 VSSD.n2377 VSSD.t816 223.315
R9359 VSSD.n1490 VSSD.t792 223.315
R9360 VSSD.n2397 VSSD.t1844 223.315
R9361 VSSD.n1975 VSSD.t686 223.315
R9362 VSSD.n2098 VSSD.t922 223.315
R9363 VSSD.n2141 VSSD.t407 223.315
R9364 VSSD.n2177 VSSD.t934 223.315
R9365 VSSD.n1731 VSSD.t314 223.315
R9366 VSSD.n1774 VSSD.t826 223.315
R9367 VSSD.n1661 VSSD.t1821 223.315
R9368 VSSD.n1607 VSSD.t19 223.315
R9369 VSSD.n1625 VSSD.t201 223.315
R9370 VSSD.n244 VSSD.t539 223.315
R9371 VSSD.n313 VSSD.t1456 222.784
R9372 VSSD.n1654 VSSD.t1514 221.793
R9373 VSSD.n890 VSSD.t1859 220.952
R9374 VSSD.n501 VSSD.t1925 220.952
R9375 VSSD.n3057 VSSD.t1938 220.952
R9376 VSSD.n3058 VSSD.t1944 220.952
R9377 VSSD.n2571 VSSD.t1952 220.952
R9378 VSSD.n3765 VSSD.t1517 220.222
R9379 VSSD.n1206 VSSD.t1328 220.082
R9380 VSSD.t1026 VSSD.t1334 219.157
R9381 VSSD.t682 VSSD.t1465 219.157
R9382 VSSD.t1695 VSSD.t967 219.157
R9383 VSSD.t1581 VSSD.t699 219.157
R9384 VSSD.t678 VSSD.t1090 219.157
R9385 VSSD VSSD.t1004 219.157
R9386 VSSD.t925 VSSD.t286 219.157
R9387 VSSD.t1174 VSSD.t35 219.157
R9388 VSSD.t795 VSSD.n248 219.157
R9389 VSSD.t1248 VSSD.t1704 219.157
R9390 VSSD.n2873 VSSD.t1899 218.607
R9391 VSSD.n2879 VSSD.t1293 218.428
R9392 VSSD.n1656 VSSD.t1503 218.428
R9393 VSSD.n747 VSSD.t1924 218.308
R9394 VSSD.n3249 VSSD.t1956 218.308
R9395 VSSD.n1216 VSSD.t1985 218.308
R9396 VSSD.n2714 VSSD.t1903 218.308
R9397 VSSD.n2826 VSSD.t1909 218.308
R9398 VSSD.n2792 VSSD.t1979 218.308
R9399 VSSD.n2328 VSSD.t1983 218.308
R9400 VSSD.n2378 VSSD.t1981 218.308
R9401 VSSD.n2163 VSSD.t1868 218.308
R9402 VSSD.n1713 VSSD.t1969 218.308
R9403 VSSD.n1609 VSSD.t1916 218.308
R9404 VSSD.n1902 VSSD.t1918 218.308
R9405 VSSD.n368 VSSD.t1926 218.308
R9406 VSSD.n3677 VSSD.t1968 218.308
R9407 VSSD.n677 VSSD.t1249 217.977
R9408 VSSD.n675 VSSD.t1342 217.892
R9409 VSSD.n3375 VSSD.t1335 217.892
R9410 VSSD.n568 VSSD.t1308 217.516
R9411 VSSD.n439 VSSD.t1296 216.959
R9412 VSSD.n2546 VSSD.t1212 216.238
R9413 VSSD.n665 VSSD.t1506 215.992
R9414 VSSD.n1653 VSSD.t1515 215.905
R9415 VSSD.n561 VSSD.t1230 214.456
R9416 VSSD.n561 VSSD.t1229 214.456
R9417 VSSD.n562 VSSD.t1546 214.456
R9418 VSSD.n562 VSSD.t1545 214.456
R9419 VSSD.n3757 VSSD.t1345 214.456
R9420 VSSD.n3737 VSSD.t1344 214.456
R9421 VSSD.n39 VSSD.t1410 214.456
R9422 VSSD.n3675 VSSD.t1409 214.456
R9423 VSSD.n546 VSSD.t1250 214.456
R9424 VSSD.n711 VSSD.t1430 214.456
R9425 VSSD.n699 VSSD.t1429 214.456
R9426 VSSD.n554 VSSD.t1375 214.456
R9427 VSSD.n554 VSSD.t1374 214.456
R9428 VSSD.n596 VSSD.t1436 214.456
R9429 VSSD.n594 VSSD.t1341 214.456
R9430 VSSD.n590 VSSD.t1435 214.456
R9431 VSSD.n593 VSSD.t1475 214.456
R9432 VSSD.n589 VSSD.t1492 214.456
R9433 VSSD.n586 VSSD.t1474 214.456
R9434 VSSD.n585 VSSD.t1507 214.456
R9435 VSSD.n569 VSSD.t1491 214.456
R9436 VSSD.n567 VSSD.t1309 214.456
R9437 VSSD.n134 VSSD.t1464 214.456
R9438 VSSD.n134 VSSD.t1463 214.456
R9439 VSSD.n135 VSSD.t1489 214.456
R9440 VSSD.n135 VSSD.t1488 214.456
R9441 VSSD.n887 VSSD.t1509 214.456
R9442 VSSD.n887 VSSD.t1508 214.456
R9443 VSSD.n888 VSSD.t1407 214.456
R9444 VSSD.n888 VSSD.t1406 214.456
R9445 VSSD.n901 VSSD.t1538 214.456
R9446 VSSD.n890 VSSD.t1244 214.456
R9447 VSSD.n890 VSSD.t1243 214.456
R9448 VSSD.n894 VSSD.t1539 214.456
R9449 VSSD.n491 VSSD.t1553 214.456
R9450 VSSD.n501 VSSD.t1461 214.456
R9451 VSSD.n501 VSSD.t1460 214.456
R9452 VSSD.n512 VSSD.t1554 214.456
R9453 VSSD.n520 VSSD.t1336 214.456
R9454 VSSD.n801 VSSD.t1416 214.456
R9455 VSSD.n805 VSSD.t1415 214.456
R9456 VSSD.n776 VSSD.t1497 214.456
R9457 VSSD.n786 VSSD.t1498 214.456
R9458 VSSD.n748 VSSD.t1467 214.456
R9459 VSSD.n994 VSSD.t1466 214.456
R9460 VSSD.n981 VSSD.t1453 214.456
R9461 VSSD.n830 VSSD.t1452 214.456
R9462 VSSD.n936 VSSD.t1253 214.456
R9463 VSSD.n955 VSSD.t1252 214.456
R9464 VSSD.n492 VSSD.t1363 214.456
R9465 VSSD.n492 VSSD.t1362 214.456
R9466 VSSD.n494 VSSD.t1274 214.456
R9467 VSSD.n494 VSSD.t1273 214.456
R9468 VSSD.n3250 VSSD.t1271 214.456
R9469 VSSD.n3260 VSSD.t1270 214.456
R9470 VSSD.n3250 VSSD.t1560 214.456
R9471 VSSD.n3242 VSSD.t1559 214.456
R9472 VSSD.n3241 VSSD.t1194 214.456
R9473 VSSD.n3235 VSSD.t1193 214.456
R9474 VSSD.n3229 VSSD.t1350 214.456
R9475 VSSD.n3226 VSSD.t1312 214.456
R9476 VSSD.n3218 VSSD.t1311 214.456
R9477 VSSD.n3218 VSSD.t1349 214.456
R9478 VSSD.n1298 VSSD.t1291 214.456
R9479 VSSD.n1139 VSSD.t1290 214.456
R9480 VSSD.n1215 VSSD.t1549 214.456
R9481 VSSD.n1153 VSSD.t1548 214.456
R9482 VSSD.n1289 VSSD.t1543 214.456
R9483 VSSD.n1287 VSSD.t1329 214.456
R9484 VSSD.n1237 VSSD.t1544 214.456
R9485 VSSD.n1022 VSSD.t1187 214.456
R9486 VSSD.n1033 VSSD.t1188 214.456
R9487 VSSD.n3160 VSSD.t1217 214.456
R9488 VSSD.n3170 VSSD.t1355 214.456
R9489 VSSD.n3179 VSSD.t1218 214.456
R9490 VSSD.n3156 VSSD.t1356 214.456
R9491 VSSD.n1228 VSSD.t1484 214.456
R9492 VSSD.n1228 VSSD.t1483 214.456
R9493 VSSD.n1140 VSSD.t1331 214.456
R9494 VSSD.n1140 VSSD.t1330 214.456
R9495 VSSD.n1142 VSSD.t1215 214.456
R9496 VSSD.n1142 VSSD.t1214 214.456
R9497 VSSD.n3251 VSSD.t1526 214.456
R9498 VSSD.n3251 VSSD.t1525 214.456
R9499 VSSD.n3252 VSSD.t1413 214.456
R9500 VSSD.n3252 VSSD.t1412 214.456
R9501 VSSD.n3041 VSSD.t1285 214.456
R9502 VSSD.n3025 VSSD.t1445 214.456
R9503 VSSD.n3049 VSSD.t1284 214.456
R9504 VSSD.n1077 VSSD.t1444 214.456
R9505 VSSD.n3015 VSSD.t1472 214.456
R9506 VSSD.n1080 VSSD.t1471 214.456
R9507 VSSD.n1115 VSSD.t1487 214.456
R9508 VSSD.n1123 VSSD.t1486 214.456
R9509 VSSD.n1124 VSSD.t1294 214.456
R9510 VSSD.n2872 VSSD.t1404 214.456
R9511 VSSD.n2870 VSSD.t1403 214.456
R9512 VSSD.n2863 VSSD.t1323 214.456
R9513 VSSD.n2863 VSSD.t1322 214.456
R9514 VSSD.n2864 VSSD.t1333 214.456
R9515 VSSD.n2864 VSSD.t1332 214.456
R9516 VSSD.n3057 VSSD.t1300 214.456
R9517 VSSD.n3057 VSSD.t1299 214.456
R9518 VSSD.n3058 VSSD.t1317 214.456
R9519 VSSD.n3058 VSSD.t1316 214.456
R9520 VSSD.n3077 VSSD.t1512 214.456
R9521 VSSD.n3077 VSSD.t1511 214.456
R9522 VSSD.n3078 VSSD.t1531 214.456
R9523 VSSD.n3078 VSSD.t1530 214.456
R9524 VSSD.n2715 VSSD.t1369 214.456
R9525 VSSD.n2725 VSSD.t1368 214.456
R9526 VSSD.n2715 VSSD.t1383 214.456
R9527 VSSD.n2707 VSSD.t1382 214.456
R9528 VSSD.n2706 VSSD.t1427 214.456
R9529 VSSD.n2700 VSSD.t1426 214.456
R9530 VSSD.n2695 VSSD.t1565 214.456
R9531 VSSD.n1364 VSSD.t1564 214.456
R9532 VSSD.n2791 VSSD.t1209 214.456
R9533 VSSD.n1361 VSSD.t1208 214.456
R9534 VSSD.n2825 VSSD.t1398 214.456
R9535 VSSD.n1327 VSSD.t1397 214.456
R9536 VSSD.n2558 VSSD.t1211 214.456
R9537 VSSD.n2571 VSSD.t1288 214.456
R9538 VSSD.n2571 VSSD.t1287 214.456
R9539 VSSD.n2559 VSSD.t1424 214.456
R9540 VSSD.n2559 VSSD.t1423 214.456
R9541 VSSD.n2561 VSSD.t1447 214.456
R9542 VSSD.n2561 VSSD.t1446 214.456
R9543 VSSD.n2716 VSSD.t1224 214.456
R9544 VSSD.n2716 VSSD.t1223 214.456
R9545 VSSD.n2717 VSSD.t1238 214.456
R9546 VSSD.n2717 VSSD.t1237 214.456
R9547 VSSD.n1483 VSSD.t1536 214.456
R9548 VSSD.n1483 VSSD.t1535 214.456
R9549 VSSD.n1484 VSSD.t1439 214.456
R9550 VSSD.n1484 VSSD.t1438 214.456
R9551 VSSD.n2402 VSSD.t1495 214.456
R9552 VSSD.n2402 VSSD.t1380 214.456
R9553 VSSD.n2399 VSSD.t1379 214.456
R9554 VSSD.n2395 VSSD.t1494 214.456
R9555 VSSD.n2394 VSSD.t1529 214.456
R9556 VSSD.n2387 VSSD.t1528 214.456
R9557 VSSD.n2379 VSSD.t1203 214.456
R9558 VSSD.n1419 VSSD.t1202 214.456
R9559 VSSD.n2329 VSSD.t1277 214.456
R9560 VSSD.n2317 VSSD.t1276 214.456
R9561 VSSD.n2463 VSSD.t1388 214.456
R9562 VSSD.n1413 VSSD.t1389 214.456
R9563 VSSD.n2519 VSSD.t1372 214.456
R9564 VSSD.n2519 VSSD.t1282 214.456
R9565 VSSD.n1516 VSSD.t1281 214.456
R9566 VSSD.n1515 VSSD.t1371 214.456
R9567 VSSD.n2403 VSSD.t1347 214.456
R9568 VSSD.n2403 VSSD.t1346 214.456
R9569 VSSD.n2404 VSSD.t1233 214.456
R9570 VSSD.n2404 VSSD.t1232 214.456
R9571 VSSD.n2164 VSSD.t1191 214.456
R9572 VSSD.n2161 VSSD.t1190 214.456
R9573 VSSD.n2139 VSSD.t1241 214.456
R9574 VSSD.n2230 VSSD.t1240 214.456
R9575 VSSD.n2263 VSSD.t1339 214.456
R9576 VSSD.n2109 VSSD.t1338 214.456
R9577 VSSD.n2282 VSSD.t1521 214.456
R9578 VSSD.n2068 VSSD.t1520 214.456
R9579 VSSD.n2022 VSSD.t1500 214.456
R9580 VSSD.n2025 VSSD.t1501 214.456
R9581 VSSD.n1964 VSSD.t1256 214.456
R9582 VSSD.n1964 VSSD.t1255 214.456
R9583 VSSD.n1965 VSSD.t1541 214.456
R9584 VSSD.n1965 VSSD.t1540 214.456
R9585 VSSD.n1441 VSSD.t1262 214.456
R9586 VSSD.n1441 VSSD.t1261 214.456
R9587 VSSD.n2165 VSSD.t1458 214.456
R9588 VSSD.n2165 VSSD.t1457 214.456
R9589 VSSD.n2166 VSSD.t1353 214.456
R9590 VSSD.n2166 VSSD.t1352 214.456
R9591 VSSD.n1650 VSSD.t1226 214.456
R9592 VSSD.n1834 VSSD.t1227 214.456
R9593 VSSD.n1664 VSSD.t1504 214.456
R9594 VSSD.n1694 VSSD.t1386 214.456
R9595 VSSD.n1776 VSSD.t1385 214.456
R9596 VSSD.n1705 VSSD.t1247 214.456
R9597 VSSD.n1762 VSSD.t1246 214.456
R9598 VSSD.n1706 VSSD.t1205 214.456
R9599 VSSD.n1714 VSSD.t1320 214.456
R9600 VSSD.n1724 VSSD.t1319 214.456
R9601 VSSD.n1714 VSSD.t1206 214.456
R9602 VSSD.n1715 VSSD.t1562 214.456
R9603 VSSD.n1715 VSSD.t1561 214.456
R9604 VSSD.n1717 VSSD.t1481 214.456
R9605 VSSD.n1717 VSSD.t1480 214.456
R9606 VSSD.n1619 VSSD.t1200 214.456
R9607 VSSD.n1901 VSSD.t1359 214.456
R9608 VSSD.n1590 VSSD.t1358 214.456
R9609 VSSD.n1585 VSSD.t1199 214.456
R9610 VSSD.n1584 VSSD.t1421 214.456
R9611 VSSD.n1946 VSSD.t1420 214.456
R9612 VSSD.n1608 VSSD.t1478 214.456
R9613 VSSD.n1599 VSSD.t1477 214.456
R9614 VSSD.n1600 VSSD.t1361 214.456
R9615 VSSD.n1600 VSSD.t1360 214.456
R9616 VSSD.n1601 VSSD.t1265 214.456
R9617 VSSD.n1601 VSSD.t1264 214.456
R9618 VSSD.n3609 VSSD.t1366 214.456
R9619 VSSD.n3607 VSSD.t1365 214.456
R9620 VSSD.n3606 VSSD.t1524 214.456
R9621 VSSD.n3600 VSSD.t1523 214.456
R9622 VSSD.n3599 VSSD.t1552 214.456
R9623 VSSD.n3594 VSSD.t1551 214.456
R9624 VSSD.n3587 VSSD.t1557 214.456
R9625 VSSD.n53 VSSD.t1556 214.456
R9626 VSSD.n54 VSSD.t1306 214.456
R9627 VSSD.n69 VSSD.t1305 214.456
R9628 VSSD.n70 VSSD.t1315 214.456
R9629 VSSD.n3536 VSSD.t1314 214.456
R9630 VSSD.n3529 VSSD.t1534 214.456
R9631 VSSD.n3501 VSSD.t1533 214.456
R9632 VSSD.n86 VSSD.t1185 214.456
R9633 VSSD.n92 VSSD.t1184 214.456
R9634 VSSD.n93 VSSD.t1326 214.456
R9635 VSSD.n3475 VSSD.t1325 214.456
R9636 VSSD.n3461 VSSD.t1401 214.456
R9637 VSSD.n113 VSSD.t1400 214.456
R9638 VSSD.n114 VSSD.t1221 214.456
R9639 VSSD.n120 VSSD.t1220 214.456
R9640 VSSD.n130 VSSD.t1268 214.456
R9641 VSSD.n3410 VSSD.t1267 214.456
R9642 VSSD.n3403 VSSD.t1568 214.456
R9643 VSSD.n3400 VSSD.t1567 214.456
R9644 VSSD.n266 VSSD.t1395 214.456
R9645 VSSD.n260 VSSD.t1394 214.456
R9646 VSSD.n266 VSSD.t1418 214.456
R9647 VSSD.n260 VSSD.t1417 214.456
R9648 VSSD.n259 VSSD.t1450 214.456
R9649 VSSD.n253 VSSD.t1449 214.456
R9650 VSSD.n259 VSSD.t1469 214.456
R9651 VSSD.n253 VSSD.t1468 214.456
R9652 VSSD.n252 VSSD.t1197 214.456
R9653 VSSD.n245 VSSD.t1196 214.456
R9654 VSSD.n331 VSSD.t1455 214.456
R9655 VSSD.n367 VSSD.t1442 214.456
R9656 VSSD.n212 VSSD.t1441 214.456
R9657 VSSD.n418 VSSD.t1392 214.456
R9658 VSSD.n172 VSSD.t1297 214.456
R9659 VSSD.n163 VSSD.t1391 214.456
R9660 VSSD.n267 VSSD.t1259 214.456
R9661 VSSD.n267 VSSD.t1258 214.456
R9662 VSSD.n268 VSSD.t1279 214.456
R9663 VSSD.n268 VSSD.t1278 214.456
R9664 VSSD.n0 VSSD.t1518 214.456
R9665 VSSD.n0 VSSD.t1433 214.456
R9666 VSSD.n4 VSSD.t1432 214.456
R9667 VSSD.n5 VSSD.t1236 214.456
R9668 VSSD.n3767 VSSD.t1235 214.456
R9669 VSSD.n3788 VSSD.t1377 214.456
R9670 VSSD.n3788 VSSD.t1376 214.456
R9671 VSSD.n3789 VSSD.t1303 214.456
R9672 VSSD.n3789 VSSD.t1302 214.456
R9673 VSSD.t1670 VSSD.t1387 210.728
R9674 VSSD VSSD.t280 210.728
R9675 VSSD.t1850 VSSD.t1024 210.728
R9676 VSSD.n814 VSSD.n813 209.254
R9677 VSSD.n3345 VSSD.n3344 209.254
R9678 VSSD.n876 VSSD.n875 209.254
R9679 VSSD.n1178 VSSD.n1165 209.254
R9680 VSSD.n1178 VSSD.n1166 209.254
R9681 VSSD.n3126 VSSD.n1070 209.254
R9682 VSSD.n1072 VSSD.n1071 209.254
R9683 VSSD.n3073 VSSD.n3071 209.254
R9684 VSSD.n3073 VSSD.n3072 209.254
R9685 VSSD.n2652 VSSD.n2647 209.254
R9686 VSSD.n2543 VSSD.n2542 209.254
R9687 VSSD.n2594 VSSD.n2593 209.254
R9688 VSSD.n2357 VSSD.n2356 209.254
R9689 VSSD.n2501 VSSD.n2500 209.254
R9690 VSSD.n1561 VSSD.n1497 209.254
R9691 VSSD.n1501 VSSD.n1500 209.254
R9692 VSSD.n1993 VSSD.n1468 209.254
R9693 VSSD.n1470 VSSD.n1469 209.254
R9694 VSSD.n2156 VSSD.n2155 209.254
R9695 VSSD.n2185 VSSD.n2158 209.254
R9696 VSSD.n1882 VSSD.n1881 209.254
R9697 VSSD.n471 VSSD.n470 209.254
R9698 VSSD.n155 VSSD.n154 209.254
R9699 VSSD.n349 VSSD.n222 209.254
R9700 VSSD.n241 VSSD.n240 209.254
R9701 VSSD.n35 VSSD.n34 209.254
R9702 VSSD.n3710 VSSD.n3709 209.254
R9703 VSSD.n2430 VSSD.n2429 207.974
R9704 VSSD.n1044 VSSD.n1043 207.213
R9705 VSSD.n3191 VSSD.n3185 207.213
R9706 VSSD.n3205 VSSD.n1047 207.213
R9707 VSSD.n3207 VSSD.n1046 207.213
R9708 VSSD.n2675 VSSD.n2674 206.909
R9709 VSSD.n2680 VSSD.n2679 206.909
R9710 VSSD.n2686 VSSD.n2685 206.909
R9711 VSSD.n2084 VSSD.n2060 206.909
R9712 VSSD.n2080 VSSD.n2064 206.909
R9713 VSSD.n2976 VSSD.n2975 206.823
R9714 VSSD.n2985 VSSD.n2983 206.823
R9715 VSSD.n2644 VSSD.n2643 205.899
R9716 VSSD.n2052 VSSD.n2051 205.899
R9717 VSSD.n2653 VSSD.n2646 205.481
R9718 VSSD.n2649 VSSD.n2648 205.481
R9719 VSSD.n1035 VSSD.n1034 204.692
R9720 VSSD.n2836 VSSD.n1323 204.692
R9721 VSSD.n2670 VSSD.n2669 204.692
R9722 VSSD.n2637 VSSD.n2636 204.692
R9723 VSSD.n2678 VSSD.n2677 204.692
R9724 VSSD.n2634 VSSD.n2633 204.692
R9725 VSSD.n2059 VSSD.n2058 204.692
R9726 VSSD.n1251 VSSD.n1249 204.522
R9727 VSSD.n1388 VSSD.n1387 204.457
R9728 VSSD.n549 VSSD.n548 203.526
R9729 VSSD.n859 VSSD.n858 203.526
R9730 VSSD.n988 VSSD.n749 203.526
R9731 VSSD.n3362 VSSD.n518 203.526
R9732 VSSD.n870 VSSD.n869 203.526
R9733 VSSD.n3274 VSSD.n3244 203.526
R9734 VSSD.n2910 VSSD.n1122 203.526
R9735 VSSD.n2785 VSSD.n1366 203.526
R9736 VSSD.n2739 VSSD.n2709 203.526
R9737 VSSD.n1421 VSSD.n1420 203.526
R9738 VSSD.n2461 VSSD.n1412 203.526
R9739 VSSD.n2090 VSSD.n2055 203.526
R9740 VSSD.n2257 VSSD.n2122 203.526
R9741 VSSD.n2136 VSSD.n2135 203.526
R9742 VSSD.n1738 VSSD.n1708 203.526
R9743 VSSD.n1782 VSSD.n1689 203.526
R9744 VSSD.n1666 VSSD.n1665 203.526
R9745 VSSD.n1872 VSSD.n1631 203.526
R9746 VSSD.n1579 VSSD.n1578 203.526
R9747 VSSD.n188 VSSD.n187 203.526
R9748 VSSD.n196 VSSD.n195 203.526
R9749 VSSD.n3731 VSSD.n3730 203.526
R9750 VSSD.n1247 VSSD.n1246 202.724
R9751 VSSD.n1263 VSSD.n1242 202.724
R9752 VSSD.t85 VSSD.t1175 202.299
R9753 VSSD.t747 VSSD.t1700 202.299
R9754 VSSD.t1600 VSSD.t401 202.299
R9755 VSSD.t1116 VSSD.t455 202.299
R9756 VSSD.t921 VSSD.t282 202.299
R9757 VSSD.t704 VSSD.t540 202.299
R9758 VSSD.t1736 VSSD.t45 202.299
R9759 VSSD.t573 VSSD.t1672 202.299
R9760 VSSD.t1658 VSSD.t262 202.299
R9761 VSSD.n3319 VSSD.n1023 201.458
R9762 VSSD.n1027 VSSD.n1026 201.458
R9763 VSSD.n2660 VSSD.n2642 201.458
R9764 VSSD.n2099 VSSD.n2050 201.458
R9765 VSSD.n3306 VSSD.n1032 201.129
R9766 VSSD.n1031 VSSD.n1030 201.129
R9767 VSSD.n1450 VSSD.n1448 201.129
R9768 VSSD.n2104 VSSD.n2047 201.129
R9769 VSSD.n651 VSSD.n584 200.692
R9770 VSSD.n788 VSSD.n787 200.692
R9771 VSSD.n1276 VSSD.n1235 200.692
R9772 VSSD.n3311 VSSD.n1029 200.692
R9773 VSSD.n2901 VSSD.n2900 200.692
R9774 VSSD.n2221 VSSD.n2137 200.692
R9775 VSSD.n2265 VSSD.n2264 200.692
R9776 VSSD.n1821 VSSD.n1662 200.692
R9777 VSSD.n420 VSSD.n419 200.692
R9778 VSSD.n2953 VSSD.n2952 200.516
R9779 VSSD.n2819 VSSD.n1331 200.516
R9780 VSSD.n2817 VSSD.n1335 200.516
R9781 VSSD.n2811 VSSD.n1341 200.516
R9782 VSSD.n2809 VSSD.n1344 200.516
R9783 VSSD.n1255 VSSD.n1248 200.508
R9784 VSSD.n2640 VSSD.n2639 200.508
R9785 VSSD.n1450 VSSD.n1449 200.508
R9786 VSSD.n2091 VSSD.n2054 200.508
R9787 VSSD.n2691 VSSD.n2631 200.105
R9788 VSSD.n811 VSSD.n810 199.739
R9789 VSSD.n761 VSSD.n758 199.739
R9790 VSSD.n921 VSSD.n877 199.739
R9791 VSSD.n914 VSSD.n880 199.739
R9792 VSSD.n907 VSSD.n906 199.739
R9793 VSSD.n1157 VSSD.n1155 199.739
R9794 VSSD.n1157 VSSD.n1156 199.739
R9795 VSSD.n1187 VSSD.n1185 199.739
R9796 VSSD.n1187 VSSD.n1186 199.739
R9797 VSSD.n2976 VSSD.n2974 199.739
R9798 VSSD.n2985 VSSD.n2984 199.739
R9799 VSSD.n3038 VSSD.n3028 199.739
R9800 VSSD.n3037 VSSD.n3031 199.739
R9801 VSSD.n3135 VSSD.n1066 199.739
R9802 VSSD.n3133 VSSD.n1067 199.739
R9803 VSSD.n3111 VSSD.n3060 199.739
R9804 VSSD.n3111 VSSD.n3062 199.739
R9805 VSSD.n3098 VSSD.n3067 199.739
R9806 VSSD.n3098 VSSD.n3068 199.739
R9807 VSSD.n2602 VSSD.n2601 199.739
R9808 VSSD.n2605 VSSD.n2604 199.739
R9809 VSSD.n2618 VSSD.n2617 199.739
R9810 VSSD.n2620 VSSD.n2619 199.739
R9811 VSSD.n2818 VSSD.n1332 199.739
R9812 VSSD.n2321 VSSD.n2320 199.739
R9813 VSSD.n2334 VSSD.n2315 199.739
R9814 VSSD.n2360 VSSD.n2359 199.739
R9815 VSSD.n1503 VSSD.n1502 199.739
R9816 VSSD.n1542 VSSD.n1505 199.739
R9817 VSSD.n2453 VSSD.n2384 199.739
R9818 VSSD.n1458 VSSD.n1457 199.739
R9819 VSSD.n2002 VSSD.n2001 199.739
R9820 VSSD.n1999 VSSD.n1465 199.739
R9821 VSSD.n2062 VSSD.n2061 199.739
R9822 VSSD.n2211 VSSD.n2142 199.739
R9823 VSSD.n2197 VSSD.n2150 199.739
R9824 VSSD.n2154 VSSD.n2153 199.739
R9825 VSSD.n1792 VSSD.n1791 199.739
R9826 VSSD.n1805 VSSD.n1804 199.739
R9827 VSSD.n1638 VSSD.n1637 199.739
R9828 VSSD.n1635 VSSD.n1634 199.739
R9829 VSSD.n445 VSSD.n444 199.739
R9830 VSSD.n447 VSSD.n446 199.739
R9831 VSSD.n460 VSSD.n459 199.739
R9832 VSSD.n463 VSSD.n462 199.739
R9833 VSSD.n413 VSSD.n184 199.739
R9834 VSSD.n401 VSSD.n191 199.739
R9835 VSSD.n399 VSSD.n192 199.739
R9836 VSSD.n200 VSSD.n199 199.739
R9837 VSSD.n375 VSSD.n210 199.739
R9838 VSSD.n361 VSSD.n216 199.739
R9839 VSSD.n224 VSSD.n223 199.739
R9840 VSSD.n3691 VSSD.n3690 199.739
R9841 VSSD.n3712 VSSD.n3711 199.739
R9842 VSSD.n17 VSSD.n16 199.739
R9843 VSSD.n2132 VSSD.n2131 199.536
R9844 VSSD.n179 VSSD.n177 198.696
R9845 VSSD VSSD.n3657 198.606
R9846 VSSD.n1244 VSSD.n1243 197.219
R9847 VSSD.n1264 VSSD.n1241 197.219
R9848 VSSD.n1274 VSSD.n1236 197.219
R9849 VSSD.n1114 VSSD.n1113 197.219
R9850 VSSD.n2934 VSSD.n1112 197.219
R9851 VSSD.n1101 VSSD.n1100 197.219
R9852 VSSD.n2959 VSSD.n1097 197.219
R9853 VSSD.n1337 VSSD.n1336 197.219
R9854 VSSD.t1266 VSSD 196.799
R9855 VSSD.t1324 VSSD 196.799
R9856 VSSD.t1313 VSSD 196.799
R9857 VSSD VSSD.t1364 196.799
R9858 VSSD.n1269 VSSD.n1238 196.782
R9859 VSSD.n710 VSSD.n709 196.442
R9860 VSSD.n698 VSSD.n697 196.442
R9861 VSSD.n886 VSSD.n885 196.442
R9862 VSSD.n849 VSSD.n848 196.442
R9863 VSSD.n847 VSSD.n846 196.442
R9864 VSSD.n832 VSSD.n831 196.442
R9865 VSSD.n835 VSSD.n834 196.442
R9866 VSSD.n803 VSSD.n773 196.442
R9867 VSSD.n751 VSSD.n750 196.442
R9868 VSSD.n524 VSSD.n523 196.442
R9869 VSSD.n3284 VSSD.n3240 196.442
R9870 VSSD.n2918 VSSD.n1119 196.442
R9871 VSSD.n2939 VSSD.n2935 196.442
R9872 VSSD.n2960 VSSD.n1096 196.442
R9873 VSSD.n1325 VSSD.n1324 196.442
R9874 VSSD.n1340 VSSD.n1339 196.442
R9875 VSSD.n1362 VSSD.n1360 196.442
R9876 VSSD.n2749 VSSD.n2705 196.442
R9877 VSSD.n2337 VSSD.n2336 196.442
R9878 VSSD.n2477 VSSD.n1398 196.442
R9879 VSSD.n1400 VSSD.n1399 196.442
R9880 VSSD.n1391 VSSD.n1390 196.442
R9881 VSSD.n2490 VSSD.n1393 196.442
R9882 VSSD.n1530 VSSD.n1511 196.442
R9883 VSSD.n2440 VSSD.n2391 196.442
R9884 VSSD.n2016 VSSD.n1460 196.442
R9885 VSSD.n1440 VSSD.n1439 196.442
R9886 VSSD.n1444 VSSD.n1443 196.442
R9887 VSSD.n2114 VSSD.n2113 196.442
R9888 VSSD.n2121 VSSD.n2120 196.442
R9889 VSSD.n2145 VSSD.n2144 196.442
R9890 VSSD.n1748 VSSD.n1703 196.442
R9891 VSSD.n1783 VSSD.n1688 196.442
R9892 VSSD.n1669 VSSD.n1668 196.442
R9893 VSSD.n1842 VSSD.n1652 196.442
R9894 VSSD.n1873 VSSD.n1630 196.442
R9895 VSSD.n1927 VSSD.n1582 196.442
R9896 VSSD.n1589 VSSD.n1588 196.442
R9897 VSSD.n218 VSSD.n217 196.442
R9898 VSSD.n3743 VSSD.n13 196.442
R9899 VSSD.t758 VSSD 193.87
R9900 VSSD.t1569 VSSD 193.87
R9901 VSSD.n653 VSSD.n652 190.399
R9902 VSSD.n781 VSSD.n780 190.399
R9903 VSSD.n1278 VSSD.n1277 190.399
R9904 VSSD.n3313 VSSD.n3312 190.399
R9905 VSSD.n2897 VSSD.n1127 190.399
R9906 VSSD.n2223 VSSD.n2222 190.399
R9907 VSSD.n2117 VSSD.n2116 190.399
R9908 VSSD.n1823 VSSD.n1822 190.399
R9909 VSSD.n3232 VSSD.n3231 189.556
R9910 VSSD.n2697 VSSD.n2696 189.556
R9911 VSSD.n1764 VSSD.n1696 189.556
R9912 VSSD.n783 VSSD.n782 189.481
R9913 VSSD.n3018 VSSD.n3017 189.481
R9914 VSSD.n42 VSSD.n41 189.481
R9915 VSSD.n3759 VSSD.n3758 189.481
R9916 VSSD.n1513 VSSD.n1512 189.201
R9917 VSSD.n1280 VSSD.n1279 188.429
R9918 VSSD.t1186 VSSD.t658 185.441
R9919 VSSD VSSD.t177 185.441
R9920 VSSD.t301 VSSD.t1621 185.441
R9921 VSSD.t386 VSSD.t999 185.441
R9922 VSSD.t433 VSSD.t127 185.441
R9923 VSSD.t992 VSSD.t1164 185.441
R9924 VSSD VSSD.t672 185.441
R9925 VSSD.t81 VSSD.t1757 177.012
R9926 VSSD.t996 VSSD.t535 177.012
R9927 VSSD.t120 VSSD.t41 177.012
R9928 VSSD.t988 VSSD.t94 168.583
R9929 VSSD.t1168 VSSD.t1192 168.583
R9930 VSSD.t1101 VSSD.t1019 168.583
R9931 VSSD.t845 VSSD.t1158 168.583
R9932 VSSD.t710 VSSD.t754 168.583
R9933 VSSD.t180 VSSD.t1829 168.583
R9934 VSSD.t335 VSSD.t1652 168.583
R9935 VSSD.t1796 VSSD.t164 168.583
R9936 VSSD.t594 VSSD 168.583
R9937 VSSD.t334 VSSD.t1396 168.583
R9938 VSSD.t1171 VSSD.t1425 168.583
R9939 VSSD.t1808 VSSD.t474 168.583
R9940 VSSD.t37 VSSD.t811 168.583
R9941 VSSD.t1016 VSSD.t452 168.583
R9942 VSSD.t276 VSSD.t1650 168.583
R9943 VSSD.t114 VSSD.t1151 168.583
R9944 VSSD.t226 VSSD.t1245 168.583
R9945 VSSD.t248 VSSD.t979 168.583
R9946 VSSD.t1343 VSSD.t0 168.583
R9947 VSSD.t333 VSSD.t1145 160.154
R9948 VSSD.n2693 VSSD.t623 160.154
R9949 VSSD VSSD.t885 160.154
R9950 VSSD VSSD.t813 160.154
R9951 VSSD VSSD.t402 160.154
R9952 VSSD.t1747 VSSD 160.154
R9953 VSSD.n1000 VSSD.t48 158.361
R9954 VSSD.n1048 VSSD.t865 157.291
R9955 VSSD.n3192 VSSD.t1613 155.286
R9956 VSSD.n2880 VSSD.t247 153.631
R9957 VSSD.n651 VSSD.n650 152
R9958 VSSD.n789 VSSD.n788 152
R9959 VSSD.n3311 VSSD.n3310 152
R9960 VSSD.n1276 VSSD.n1275 152
R9961 VSSD.n2900 VSSD.n2899 152
R9962 VSSD.n2266 VSSD.n2265 152
R9963 VSSD.n2221 VSSD.n2220 152
R9964 VSSD.n1821 VSSD.n1820 152
R9965 VSSD.n421 VSSD.n420 152
R9966 VSSD.t131 VSSD.t321 151.725
R9967 VSSD.t807 VSSD.t527 151.725
R9968 VSSD.t1485 VSSD.t1848 151.725
R9969 VSSD.t1143 VSSD.t592 151.725
R9970 VSSD.t360 VSSD.t1073 151.725
R9971 VSSD.t643 VSSD.t596 151.725
R9972 VSSD.t358 VSSD.t1069 151.725
R9973 VSSD.t803 VSSD.t1075 151.725
R9974 VSSD.t797 VSSD.t1071 151.725
R9975 VSSD.t190 VSSD.t350 151.725
R9976 VSSD.t1207 VSSD.t788 151.725
R9977 VSSD.t1758 VSSD.t1156 151.725
R9978 VSSD VSSD.t1795 151.725
R9979 VSSD.t159 VSSD.t861 151.725
R9980 VSSD.t1091 VSSD.t119 151.725
R9981 VSSD.t1773 VSSD.t412 151.725
R9982 VSSD.t1774 VSSD.t415 151.725
R9983 VSSD.n2962 VSSD.t1830 149.762
R9984 VSSD.n1345 VSSD.t154 149.762
R9985 VSSD.n1256 VSSD.t1643 146.464
R9986 VSSD.t1031 VSSD 143.296
R9987 VSSD.t1012 VSSD.t1707 143.296
R9988 VSSD.t1066 VSSD.t648 143.296
R9989 VSSD.t689 VSSD.t1709 143.296
R9990 VSSD.t1794 VSSD.t1734 143.296
R9991 VSSD.t881 VSSD.t203 143.296
R9992 VSSD.t855 VSSD.t1694 143.296
R9993 VSSD.t368 VSSD.t712 143.296
R9994 VSSD.t424 VSSD.t937 143.296
R9995 VSSD.t1566 VSSD 135.412
R9996 VSSD VSSD.n96 135.412
R9997 VSSD VSSD.n73 135.412
R9998 VSSD.n3657 VSSD 135.412
R9999 VSSD.t140 VSSD.t410 134.867
R10000 VSSD.t422 VSSD.t1615 134.867
R10001 VSSD.t1038 VSSD.t388 134.867
R10002 VSSD.t1153 VSSD.t1110 134.867
R10003 VSSD.t562 VSSD.t691 134.867
R10004 VSSD.n3398 VSSD 133.607
R10005 VSSD.t619 VSSD.t1781 126.438
R10006 VSSD.t1612 VSSD.t1064 126.438
R10007 VSSD.t864 VSSD.t1010 126.438
R10008 VSSD.t1693 VSSD.t102 126.438
R10009 VSSD.n1413 VSSD.t1910 121.927
R10010 VSSD.n2025 VSSD.t1904 121.927
R10011 VSSD.t796 VSSD.t879 118.008
R10012 VSSD.t592 VSSD 118.008
R10013 VSSD.t975 VSSD.t347 118.008
R10014 VSSD.t1499 VSSD.t484 118.008
R10015 VSSD.t470 VSSD.t298 118.008
R10016 VSSD.t706 VSSD.t895 118.008
R10017 VSSD.t213 VSSD.t872 118.008
R10018 VSSD.n783 VSSD.n742 117.334
R10019 VSSD.n3019 VSSD.n3018 117.334
R10020 VSSD.n43 VSSD.n42 117.334
R10021 VSSD.n3759 VSSD.n7 117.334
R10022 VSSD.n3225 VSSD.t1951 116.734
R10023 VSSD.n2520 VSSD.t1955 116.734
R10024 VSSD.n2401 VSSD.t1919 116.734
R10025 VSSD.n1769 VSSD.t1906 116.734
R10026 VSSD.n165 VSSD.t1967 116.734
R10027 VSSD.n3042 VSSD.t1953 112.349
R10028 VSSD.t1690 VSSD.t302 109.579
R10029 VSSD.t1688 VSSD.t34 109.579
R10030 VSSD.n894 VSSD.t1895 102.695
R10031 VSSD.n251 VSSD.t1871 102.379
R10032 VSSD.t508 VSSD.n826 101.15
R10033 VSSD.t726 VSSD.t390 101.15
R10034 VSSD.t1162 VSSD.t392 101.15
R10035 VSSD.t402 VSSD.t323 101.15
R10036 VSSD.t459 VSSD.t453 101.15
R10037 VSSD.t54 VSSD.t1747 101.15
R10038 VSSD.t74 VSSD.t1035 101.15
R10039 VSSD.n3301 VSSD.n3232 100.572
R10040 VSSD.n2766 VSSD.n2697 100.572
R10041 VSSD.n1765 VSSD.n1764 100.572
R10042 VSSD.n2546 VSSD.t1962 100.209
R10043 VSSD.n548 VSSD.t1779 100.001
R10044 VSSD.n858 VSSD.t1059 100.001
R10045 VSSD.n749 VSSD.t1061 100.001
R10046 VSSD.n813 VSSD.t505 100.001
R10047 VSSD.n3344 VSSD.t496 100.001
R10048 VSSD.n518 VSSD.t1594 100.001
R10049 VSSD.n869 VSSD.t1782 100.001
R10050 VSSD.n875 VSSD.t880 100.001
R10051 VSSD.n1165 VSSD.t1588 100.001
R10052 VSSD.n1166 VSSD.t1140 100.001
R10053 VSSD.n3244 VSSD.t490 100.001
R10054 VSSD.n1122 VSSD.t1592 100.001
R10055 VSSD.n2975 VSSD.t1057 100.001
R10056 VSSD.n2983 VSSD.t216 100.001
R10057 VSSD.n1070 VSSD.t253 100.001
R10058 VSSD.n1071 VSSD.t261 100.001
R10059 VSSD.n3071 VSSD.t479 100.001
R10060 VSSD.n3072 VSSD.t1595 100.001
R10061 VSSD.n2647 VSSD.t511 100.001
R10062 VSSD.n2542 VSSD.t1138 100.001
R10063 VSSD.n2593 VSSD.t167 100.001
R10064 VSSD.n1366 VSSD.t1683 100.001
R10065 VSSD.n2709 VSSD.t507 100.001
R10066 VSSD.n2429 VSSD.t255 100.001
R10067 VSSD.n2356 VSSD.t222 100.001
R10068 VSSD.n1420 VSSD.t1667 100.001
R10069 VSSD.n1412 VSSD.t1671 100.001
R10070 VSSD.n2500 VSSD.t555 100.001
R10071 VSSD.n1497 VSSD.t245 100.001
R10072 VSSD.n1500 VSSD.t553 100.001
R10073 VSSD.n1468 VSSD.t274 100.001
R10074 VSSD.n1469 VSSD.t231 100.001
R10075 VSSD.n2055 VSSD.t1651 100.001
R10076 VSSD.n2122 VSSD.t212 100.001
R10077 VSSD.n2135 VSSD.t559 100.001
R10078 VSSD.n2155 VSSD.t210 100.001
R10079 VSSD.n2158 VSSD.t316 100.001
R10080 VSSD.n1708 VSSD.t1661 100.001
R10081 VSSD.n1689 VSSD.t1655 100.001
R10082 VSSD.n1665 VSSD.t1665 100.001
R10083 VSSD.n1631 VSSD.t265 100.001
R10084 VSSD.n1881 VSSD.t233 100.001
R10085 VSSD.n1578 VSSD.t1649 100.001
R10086 VSSD.n470 VSSD.t239 100.001
R10087 VSSD.n154 VSSD.t257 100.001
R10088 VSSD.n187 VSSD.t898 100.001
R10089 VSSD.n195 VSSD.t1675 100.001
R10090 VSSD.n222 VSSD.t1689 100.001
R10091 VSSD.n240 VSSD.t1679 100.001
R10092 VSSD.n34 VSSD.t481 100.001
R10093 VSSD.n3709 VSSD.t1788 100.001
R10094 VSSD.n3730 VSSD.t1055 100.001
R10095 VSSD.n3176 VSSD.t1873 99.7825
R10096 VSSD.n3023 VSSD.t1887 99.7825
R10097 VSSD.n1381 VSSD.t1945 99.7825
R10098 VSSD.n3783 VSSD.t1935 99.7825
R10099 VSSD.n499 VSSD.t1890 96.5628
R10100 VSSD.n1833 VSSD.t1965 94.8164
R10101 VSSD.n3228 VSSD.t1966 94.8077
R10102 VSSD.n3157 VSSD.t1949 94.8077
R10103 VSSD.t679 VSSD 92.7208
R10104 VSSD.t1122 VSSD.t275 92.7208
R10105 VSSD.t372 VSSD 92.7208
R10106 VSSD VSSD.t656 92.7208
R10107 VSSD.t1806 VSSD.t1419 92.7208
R10108 VSSD VSSD.t103 84.2917
R10109 VSSD.t605 VSSD.t68 84.2917
R10110 VSSD.t837 VSSD.t941 84.2917
R10111 VSSD.t404 VSSD.t1239 84.2917
R10112 VSSD.t16 VSSD.t1476 84.2917
R10113 VSSD.t1732 VSSD.t1502 84.2917
R10114 VSSD.t1384 VSSD.t829 84.2917
R10115 VSSD.t1181 VSSD 75.8626
R10116 VSSD.t1056 VSSD.t1656 75.8626
R10117 VSSD.t162 VSSD.t215 75.8626
R10118 VSSD.t510 VSSD.t1147 75.8626
R10119 VSSD VSSD.t301 75.8626
R10120 VSSD.t667 VSSD.t1697 75.8626
R10121 VSSD.t733 VSSD.t471 75.8626
R10122 VSSD.t693 VSSD.t1746 75.8626
R10123 VSSD.n697 VSSD.t494 72.8576
R10124 VSSD.n846 VSSD.t492 72.8576
R10125 VSSD.n831 VSSD.t169 72.8576
R10126 VSSD.n773 VSSD.t1597 72.8576
R10127 VSSD.n750 VSSD.t509 72.8576
R10128 VSSD.n523 VSSD.t1728 72.8576
R10129 VSSD.n877 VSSD.t1053 72.8576
R10130 VSSD.n880 VSSD.t1784 72.8576
R10131 VSSD.n1185 VSSD.t1780 72.8576
R10132 VSSD.n1186 VSSD.t918 72.8576
R10133 VSSD.n3240 VSSD.t1142 72.8576
R10134 VSSD.n1119 VSSD.t1590 72.8576
R10135 VSSD.n2974 VSSD.t1657 72.8576
R10136 VSSD.n2984 VSSD.t163 72.8576
R10137 VSSD.n1066 VSSD.t1653 72.8576
R10138 VSSD.n1067 VSSD.t251 72.8576
R10139 VSSD.n3067 VSSD.t1731 72.8576
R10140 VSSD.n3068 VSSD.t515 72.8576
R10141 VSSD.n1324 VSSD.t1786 72.8576
R10142 VSSD.n2601 VSSD.t498 72.8576
R10143 VSSD.n2604 VSSD.t165 72.8576
R10144 VSSD.n2631 VSSD.t557 72.8576
R10145 VSSD.n1360 VSSD.t270 72.8576
R10146 VSSD.n2705 VSSD.t1132 72.8576
R10147 VSSD.n2336 VSSD.t1677 72.8576
R10148 VSSD.n2359 VSSD.t892 72.8576
R10149 VSSD.n1398 VSSD.t272 72.8576
R10150 VSSD.n1393 VSSD.t220 72.8576
R10151 VSSD.n1387 VSSD.t318 72.8576
R10152 VSSD.n1502 VSSD.t218 72.8576
R10153 VSSD.n1505 VSSD.t229 72.8576
R10154 VSSD.n2391 VSSD.t1681 72.8576
R10155 VSSD.n2001 VSSD.t1663 72.8576
R10156 VSSD.n1465 VSSD.t1669 72.8576
R10157 VSSD.n2061 VSSD.t561 72.8576
R10158 VSSD.n2113 VSSD.t243 72.8576
R10159 VSSD.n2131 VSSD.t1687 72.8576
R10160 VSSD.n2150 VSSD.t1685 72.8576
R10161 VSSD.n2153 VSSD.t224 72.8576
R10162 VSSD.n1703 VSSD.t237 72.8576
R10163 VSSD.n1791 VSSD.t214 72.8576
R10164 VSSD.n1804 VSSD.t896 72.8576
R10165 VSSD.n1634 VSSD.t259 72.8576
R10166 VSSD.n1630 VSSD.t1673 72.8576
R10167 VSSD.n1582 VSSD.t235 72.8576
R10168 VSSD.n459 VSSD.t249 72.8576
R10169 VSSD.n462 VSSD.t241 72.8576
R10170 VSSD.n191 VSSD.t1659 72.8576
R10171 VSSD.n192 VSSD.t263 72.8576
R10172 VSSD.n217 VSSD.t890 72.8576
R10173 VSSD.n223 VSSD.t894 72.8576
R10174 VSSD.n3690 VSSD.t1730 72.8576
R10175 VSSD.n3711 VSSD.t483 72.8576
R10176 VSSD.n13 VSSD.t513 72.8576
R10177 VSSD.n548 VSSD.t806 70.0005
R10178 VSSD.n858 VSSD.t1715 70.0005
R10179 VSSD.n749 VSSD.t449 70.0005
R10180 VSSD.n813 VSSD.t411 70.0005
R10181 VSSD.n3344 VSSD.t739 70.0005
R10182 VSSD.n518 VSSD.t640 70.0005
R10183 VSSD.n869 VSSD.t207 70.0005
R10184 VSSD.n875 VSSD.t568 70.0005
R10185 VSSD.n1165 VSSD.t1644 70.0005
R10186 VSSD.n1166 VSSD.t981 70.0005
R10187 VSSD.n3244 VSSD.t309 70.0005
R10188 VSSD.n1122 VSSD.t184 70.0005
R10189 VSSD.n2975 VSSD.t966 70.0005
R10190 VSSD.n2983 VSSD.t290 70.0005
R10191 VSSD.n1070 VSSD.t615 70.0005
R10192 VSSD.n1071 VSSD.t7 70.0005
R10193 VSSD.n3071 VSSD.t676 70.0005
R10194 VSSD.n3072 VSSD.t767 70.0005
R10195 VSSD.n2647 VSSD.t348 70.0005
R10196 VSSD.n2542 VSSD.t1080 70.0005
R10197 VSSD.n2593 VSSD.t972 70.0005
R10198 VSSD.n1366 VSSD.t1765 70.0005
R10199 VSSD.n2709 VSSD.t591 70.0005
R10200 VSSD.n2429 VSSD.t1842 70.0005
R10201 VSSD.n2356 VSSD.t40 70.0005
R10202 VSSD.n1420 VSSD.t812 70.0005
R10203 VSSD.n1412 VSSD.t570 70.0005
R10204 VSSD.n2500 VSSD.t886 70.0005
R10205 VSSD.n1497 VSSD.t440 70.0005
R10206 VSSD.n1500 VSSD.t82 70.0005
R10207 VSSD.n1468 VSSD.t997 70.0005
R10208 VSSD.n1469 VSSD.t296 70.0005
R10209 VSSD.n2055 VSSD.t924 70.0005
R10210 VSSD.n2122 VSSD.t836 70.0005
R10211 VSSD.n2135 VSSD.t405 70.0005
R10212 VSSD.n2155 VSSD.t42 70.0005
R10213 VSSD.n2158 VSSD.t932 70.0005
R10214 VSSD.n1708 VSSD.t332 70.0005
R10215 VSSD.n1689 VSSD.t828 70.0005
R10216 VSSD.n1665 VSSD.t914 70.0005
R10217 VSSD.n1631 VSSD.t574 70.0005
R10218 VSSD.n1881 VSSD.t454 70.0005
R10219 VSSD.n1578 VSSD.t670 70.0005
R10220 VSSD.n470 VSSD.t1756 70.0005
R10221 VSSD.n154 VSSD.t353 70.0005
R10222 VSSD.n187 VSSD.t369 70.0005
R10223 VSSD.n195 VSSD.t938 70.0005
R10224 VSSD.n222 VSSD.t696 70.0005
R10225 VSSD.n240 VSSD.t537 70.0005
R10226 VSSD.n34 VSSD.t126 70.0005
R10227 VSSD.n3709 VSSD.t1798 70.0005
R10228 VSSD.n3730 VSSD.t1170 70.0005
R10229 VSSD VSSD.t1181 67.4335
R10230 VSSD.n1099 VSSD.t756 67.4335
R10231 VSSD.t990 VSSD.t965 67.4335
R10232 VSSD.t289 VSSD.t399 67.4335
R10233 VSSD.t20 VSSD.t1569 67.4335
R10234 VSSD.t4 VSSD.t616 67.4335
R10235 VSSD.t1077 VSSD.t949 67.4335
R10236 VSSD.t142 VSSD.t1702 67.4335
R10237 VSSD.t1716 VSSD.t849 67.4335
R10238 VSSD.t533 VSSD.t1691 67.4335
R10239 VSSD.t835 VSSD.t875 67.4335
R10240 VSSD.t1046 VSSD.t354 67.4335
R10241 VSSD.t1766 VSSD.t52 67.4335
R10242 VSSD.t1155 VSSD.t1729 67.4335
R10243 VSSD.t482 VSSD.t434 67.4335
R10244 VSSD.n1280 VSSD.n1233 61.4405
R10245 VSSD.n697 VSSD.t320 60.5809
R10246 VSSD.n846 VSSD.t680 60.5809
R10247 VSSD.n831 VSSD.t11 60.5809
R10248 VSSD.n773 VSSD.t196 60.5809
R10249 VSSD.n750 VSSD.t989 60.5809
R10250 VSSD.n523 VSSD.t1792 60.5809
R10251 VSSD.n877 VSSD.t97 60.5809
R10252 VSSD.n880 VSSD.t158 60.5809
R10253 VSSD.n1185 VSSD.t1812 60.5809
R10254 VSSD.n1186 VSSD.t854 60.5809
R10255 VSSD.n3240 VSSD.t579 60.5809
R10256 VSSD.n1119 VSSD.t1849 60.5809
R10257 VSSD.n2974 VSSD.t991 60.5809
R10258 VSSD.n2984 VSSD.t400 60.5809
R10259 VSSD.n1066 VSSD.t701 60.5809
R10260 VSSD.n1067 VSSD.t1166 60.5809
R10261 VSSD.n3067 VSSD.t294 60.5809
R10262 VSSD.n3068 VSSD.t750 60.5809
R10263 VSSD.n1324 VSSD.t61 60.5809
R10264 VSSD.n2601 VSSD.t904 60.5809
R10265 VSSD.n2604 VSSD.t1790 60.5809
R10266 VSSD.n1360 VSSD.t789 60.5809
R10267 VSSD.n2705 VSSD.t172 60.5809
R10268 VSSD.n2336 VSSD.t1698 60.5809
R10269 VSSD.n2359 VSSD.t850 60.5809
R10270 VSSD.n1398 VSSD.t1039 60.5809
R10271 VSSD.n1393 VSSD.t1616 60.5809
R10272 VSSD.n1502 VSSD.t1701 60.5809
R10273 VSSD.n1505 VSSD.t1809 60.5809
R10274 VSSD.n2391 VSSD.t330 60.5809
R10275 VSSD.n2001 VSSD.t1017 60.5809
R10276 VSSD.n1465 VSSD.t456 60.5809
R10277 VSSD.n2061 VSSD.t1739 60.5809
R10278 VSSD.n2113 VSSD.t116 60.5809
R10279 VSSD.n2131 VSSD.t749 60.5809
R10280 VSSD.n2150 VSSD.t1152 60.5809
R10281 VSSD.n2153 VSSD.t705 60.5809
R10282 VSSD.n1703 VSSD.t772 60.5809
R10283 VSSD.n1791 VSSD.t419 60.5809
R10284 VSSD.n1804 VSSD.t735 60.5809
R10285 VSSD.n1634 VSSD.t612 60.5809
R10286 VSSD.n1630 VSSD.t1724 60.5809
R10287 VSSD.n1582 VSSD.t447 60.5809
R10288 VSSD.n459 VSSD.t1719 60.5809
R10289 VSSD.n462 VSSD.t583 60.5809
R10290 VSSD.n191 VSSD.t118 60.5809
R10291 VSSD.n192 VSSD.t1754 60.5809
R10292 VSSD.n217 VSSD.t63 60.5809
R10293 VSSD.n223 VSSD.t176 60.5809
R10294 VSSD.n3690 VSSD.t1098 60.5809
R10295 VSSD.n3711 VSSD.t1611 60.5809
R10296 VSSD.n13 VSSD.t946 60.5809
R10297 VSSD.t548 VSSD.t1165 59.0043
R10298 VSSD.t432 VSSD.t903 59.0043
R10299 VSSD.t149 VSSD 59.0043
R10300 VSSD.t395 VSSD.t915 59.0043
R10301 VSSD.t604 VSSD.t1640 59.0043
R10302 VSSD.t366 VSSD.t743 59.0043
R10303 VSSD.t264 VSSD.t1723 59.0043
R10304 VSSD.t582 VSSD.t472 59.0043
R10305 VSSD.t871 VSSD.t1029 50.5752
R10306 VSSD.t300 VSSD.t611 50.5752
R10307 VSSD.t132 VSSD.t1112 42.1461
R10308 VSSD VSSD.t1596 42.1461
R10309 VSSD.t266 VSSD.t170 42.1461
R10310 VSSD.t1696 VSSD.t99 42.1461
R10311 VSSD VSSD.t179 42.1461
R10312 VSSD.t634 VSSD 42.1461
R10313 VSSD.n1834 VSSD.n1833 41.022
R10314 VSSD.n1032 VSSD.t661 40.0005
R10315 VSSD.n1032 VSSD.t655 40.0005
R10316 VSSD.n1249 VSSD.t373 40.0005
R10317 VSSD.n1249 VSSD.t375 40.0005
R10318 VSSD.n1034 VSSD.t824 40.0005
R10319 VSSD.n1034 VSSD.t663 40.0005
R10320 VSSD.n1030 VSSD.t89 40.0005
R10321 VSSD.n1030 VSSD.t822 40.0005
R10322 VSSD.n1023 VSSD.t91 40.0005
R10323 VSSD.n1023 VSSD.t371 40.0005
R10324 VSSD.n1026 VSSD.t93 40.0005
R10325 VSSD.n1248 VSSD.t653 40.0005
R10326 VSSD.n1248 VSSD.t820 40.0005
R10327 VSSD.n1246 VSSD.t462 40.0005
R10328 VSSD.n1246 VSSD.t377 40.0005
R10329 VSSD.n1242 VSSD.t906 40.0005
R10330 VSSD.n1242 VSSD.t29 40.0005
R10331 VSSD.n2643 VSSD.t138 40.0005
R10332 VSSD.n2646 VSSD.t1148 40.0005
R10333 VSSD.n2646 VSSD.t978 40.0005
R10334 VSSD.n2648 VSSD.t976 40.0005
R10335 VSSD.n2648 VSSD.t134 40.0005
R10336 VSSD.n1323 VSSD.t1146 40.0005
R10337 VSSD.n1323 VSSD.t802 40.0005
R10338 VSSD.n2642 VSSD.t193 40.0005
R10339 VSSD.n2642 VSSD.t189 40.0005
R10340 VSSD.n2639 VSSD.t187 40.0005
R10341 VSSD.n2639 VSSD.t136 40.0005
R10342 VSSD.n2669 VSSD.t798 40.0005
R10343 VSSD.n2669 VSSD.t191 40.0005
R10344 VSSD.n2636 VSSD.t1076 40.0005
R10345 VSSD.n2636 VSSD.t1072 40.0005
R10346 VSSD.n2674 VSSD.t359 40.0005
R10347 VSSD.n2674 VSSD.t804 40.0005
R10348 VSSD.n2677 VSSD.t597 40.0005
R10349 VSSD.n2677 VSSD.t1070 40.0005
R10350 VSSD.n2679 VSSD.t361 40.0005
R10351 VSSD.n2679 VSSD.t644 40.0005
R10352 VSSD.n2633 VSSD.t593 40.0005
R10353 VSSD.n2633 VSSD.t1074 40.0005
R10354 VSSD.n2685 VSSD.t429 40.0005
R10355 VSSD.n2685 VSSD.t595 40.0005
R10356 VSSD.n1449 VSSD.t485 40.0005
R10357 VSSD.n1449 VSSD.t610 40.0005
R10358 VSSD.n1448 VSSD.t285 40.0005
R10359 VSSD.n1448 VSSD.t281 40.0005
R10360 VSSD.n2047 VSSD.t1607 40.0005
R10361 VSSD.n2047 VSSD.t287 40.0005
R10362 VSSD.n2050 VSSD.t1609 40.0005
R10363 VSSD.n2051 VSSD.t1605 40.0005
R10364 VSSD.n2051 VSSD.t1851 40.0005
R10365 VSSD.n2054 VSSD.t277 40.0005
R10366 VSSD.n2054 VSSD.t487 40.0005
R10367 VSSD.n2058 VSSD.t1603 40.0005
R10368 VSSD.n2058 VSSD.t279 40.0005
R10369 VSSD.n2060 VSSD.t606 40.0005
R10370 VSSD.n2060 VSSD.t27 40.0005
R10371 VSSD.n2064 VSSD.t25 40.0005
R10372 VSSD.n2064 VSSD.t23 40.0005
R10373 VSSD.n3758 VSSD.t944 38.5719
R10374 VSSD.n3758 VSSD.t781 38.5719
R10375 VSSD.n709 VSSD.t519 38.5719
R10376 VSSD.n709 VSSD.t732 38.5719
R10377 VSSD.n885 VSSD.t529 38.5719
R10378 VSSD.n885 VSSD.t599 38.5719
R10379 VSSD.n848 VSSD.t1847 38.5719
R10380 VSSD.n848 VSSD.t383 38.5719
R10381 VSSD.n834 VSSD.t385 38.5719
R10382 VSSD.n834 VSSD.t722 38.5719
R10383 VSSD.n782 VSSD.t1095 38.5719
R10384 VSSD.n782 VSSD.t785 38.5719
R10385 VSSD.n810 VSSD.t141 38.5719
R10386 VSSD.n810 VSSD.t787 38.5719
R10387 VSSD.n758 VSSD.t1113 38.5719
R10388 VSSD.n758 VSSD.t95 38.5719
R10389 VSSD.n906 VSSD.t808 38.5719
R10390 VSSD.n906 VSSD.t852 38.5719
R10391 VSSD.n1026 VSSD.t659 38.5719
R10392 VSSD.n1155 VSSD.t920 38.5719
R10393 VSSD.n1155 VSSD.t146 38.5719
R10394 VSSD.n1156 VSSD.t1022 38.5719
R10395 VSSD.n1156 VSSD.t145 38.5719
R10396 VSSD.n3231 VSSD.t603 38.5719
R10397 VSSD.n3231 VSSD.t521 38.5719
R10398 VSSD.n3017 VSSD.t698 38.5719
R10399 VSSD.n3017 VSSD.t148 38.5719
R10400 VSSD.n2935 VSSD.t1020 38.5719
R10401 VSSD.n2935 VSSD.t1159 38.5719
R10402 VSSD.n1096 VSSD.t711 38.5719
R10403 VSSD.n1096 VSSD.t181 38.5719
R10404 VSSD.n3028 VSSD.t1584 38.5719
R10405 VSSD.n3028 VSSD.t1570 38.5719
R10406 VSSD.n3031 VSSD.t21 38.5719
R10407 VSSD.n3031 VSSD.t1776 38.5719
R10408 VSSD.n3060 VSSD.t1161 38.5719
R10409 VSSD.n3060 VSSD.t681 38.5719
R10410 VSSD.n3062 VSSD.t1838 38.5719
R10411 VSSD.n3062 VSSD.t345 38.5719
R10412 VSSD.n2643 VSSD.t974 38.5719
R10413 VSSD.n2617 VSSD.t638 38.5719
R10414 VSSD.n2617 VSSD.t143 38.5719
R10415 VSSD.n2619 VSSD.t1703 38.5719
R10416 VSSD.n2619 VSSD.t1837 38.5719
R10417 VSSD.n1332 VSSD.t727 38.5719
R10418 VSSD.n1332 VSSD.t1163 38.5719
R10419 VSSD.n1339 VSSD.t630 38.5719
R10420 VSSD.n1339 VSSD.t1744 38.5719
R10421 VSSD.n2696 VSSD.t1835 38.5719
R10422 VSSD.n2696 VSSD.t79 38.5719
R10423 VSSD.n2320 VSSD.t957 38.5719
R10424 VSSD.n2320 VSSD.t178 38.5719
R10425 VSSD.n2315 VSSD.t1622 38.5719
R10426 VSSD.n2315 VSSD.t1049 38.5719
R10427 VSSD.n2384 VSSD.t1637 38.5719
R10428 VSSD.n2384 VSSD.t703 38.5719
R10429 VSSD.n1399 VSSD.t842 38.5719
R10430 VSSD.n1399 VSSD.t389 38.5719
R10431 VSSD.n1390 VSSD.t423 38.5719
R10432 VSSD.n1390 VSSD.t1136 38.5719
R10433 VSSD.n1511 VSSD.t576 38.5719
R10434 VSSD.n1511 VSSD.t465 38.5719
R10435 VSSD.n1512 VSSD.t778 38.5719
R10436 VSSD.n1512 VSSD.t1007 38.5719
R10437 VSSD.n1457 VSSD.t1115 38.5719
R10438 VSSD.n1457 VSSD.t1005 38.5719
R10439 VSSD.n1460 VSSD.t1802 38.5719
R10440 VSSD.n1460 VSSD.t469 38.5719
R10441 VSSD.n2050 VSSD.t283 38.5719
R10442 VSSD.n1439 VSSD.t112 38.5719
R10443 VSSD.n1439 VSSD.t427 38.5719
R10444 VSSD.n1443 VSSD.t878 38.5719
R10445 VSSD.n1443 VSSD.t928 38.5719
R10446 VSSD.n2120 VSSD.t876 38.5719
R10447 VSSD.n2120 VSSD.t1125 38.5719
R10448 VSSD.n2142 VSSD.t324 38.5719
R10449 VSSD.n2142 VSSD.t542 38.5719
R10450 VSSD.n2144 VSSD.t1639 38.5719
R10451 VSSD.n2144 VSSD.t1750 38.5719
R10452 VSSD.n1696 VSSD.t742 38.5719
R10453 VSSD.n1696 VSSD.t1619 38.5719
R10454 VSSD.n1688 VSSD.t397 38.5719
R10455 VSSD.n1688 VSSD.t33 38.5719
R10456 VSSD.n1668 VSSD.t1626 38.5719
R10457 VSSD.n1668 VSSD.t833 38.5719
R10458 VSSD.n1652 VSSD.t444 38.5719
R10459 VSSD.n1652 VSSD.t1130 38.5719
R10460 VSSD.n1637 VSSD.t299 38.5719
R10461 VSSD.n1637 VSSD.t36 38.5719
R10462 VSSD.n1588 VSSD.t1579 38.5719
R10463 VSSD.n1588 VSSD.t467 38.5719
R10464 VSSD.n444 VSSD.t1767 38.5719
R10465 VSSD.n444 VSSD.t59 38.5719
R10466 VSSD.n446 VSSD.t1120 38.5719
R10467 VSSD.n446 VSSD.t53 38.5719
R10468 VSSD.n184 VSSD.t1003 38.5719
R10469 VSSD.n184 VSSD.t414 38.5719
R10470 VSSD.n199 VSSD.t328 38.5719
R10471 VSSD.n199 VSSD.t57 38.5719
R10472 VSSD.n210 VSSD.t55 38.5719
R10473 VSSD.n210 VSSD.t633 38.5719
R10474 VSSD.n216 VSSD.t626 38.5719
R10475 VSSD.n216 VSSD.t564 38.5719
R10476 VSSD.n41 VSSD.t601 38.5719
R10477 VSSD.n41 VSSD.t1033 38.5719
R10478 VSSD.n16 VSSD.t73 38.5719
R10479 VSSD.n16 VSSD.t783 38.5719
R10480 VSSD.n857 VSSD.n856 34.6358
R10481 VSSD.n850 VSSD.n838 34.6358
R10482 VSSD.n970 VSSD.n836 34.6358
R10483 VSSD.n970 VSSD.n969 34.6358
R10484 VSSD.n976 VSSD.n975 34.6358
R10485 VSSD.n819 VSSD.n769 34.6358
R10486 VSSD.n3350 VSSD.n525 34.6358
R10487 VSSD.n3346 VSSD.n525 34.6358
R10488 VSSD.n928 VSSD.n927 34.6358
R10489 VSSD.n927 VSSD.n926 34.6358
R10490 VSSD.n926 VSSD.n873 34.6358
R10491 VSSD.n920 VSSD.n919 34.6358
R10492 VSSD.n919 VSSD.n878 34.6358
R10493 VSSD.n915 VSSD.n878 34.6358
R10494 VSSD.n913 VSSD.n912 34.6358
R10495 VSSD.n3208 VSSD.n1044 34.6358
R10496 VSSD.n1254 VSSD.n1252 34.6358
R10497 VSSD.n1258 VSSD.n1257 34.6358
R10498 VSSD.n1262 VSSD.n1261 34.6358
R10499 VSSD.n1192 VSSD.n1161 34.6358
R10500 VSSD.n1193 VSSD.n1192 34.6358
R10501 VSSD.n1194 VSSD.n1193 34.6358
R10502 VSSD.n1194 VSSD.n1159 34.6358
R10503 VSSD.n1198 VSSD.n1159 34.6358
R10504 VSSD.n1179 VSSD.n1163 34.6358
R10505 VSSD.n1183 VSSD.n1163 34.6358
R10506 VSSD.n1184 VSSD.n1183 34.6358
R10507 VSSD.n1188 VSSD.n1184 34.6358
R10508 VSSD.n1176 VSSD.n1137 34.6358
R10509 VSSD.n1177 VSSD.n1176 34.6358
R10510 VSSD.n2933 VSSD.n2932 34.6358
R10511 VSSD.n2954 VSSD.n2951 34.6358
R10512 VSSD.n2958 VSSD.n1098 34.6358
R10513 VSSD.n2972 VSSD.n1092 34.6358
R10514 VSSD.n2973 VSSD.n2972 34.6358
R10515 VSSD.n2977 VSSD.n1090 34.6358
R10516 VSSD.n2981 VSSD.n1090 34.6358
R10517 VSSD.n2982 VSSD.n2981 34.6358
R10518 VSSD.n2986 VSSD.n2982 34.6358
R10519 VSSD.n2994 VSSD.n1088 34.6358
R10520 VSSD.n2996 VSSD.n2994 34.6358
R10521 VSSD.n3144 VSSD.n1059 34.6358
R10522 VSSD.n3144 VSSD.n3143 34.6358
R10523 VSSD.n3143 VSSD.n1060 34.6358
R10524 VSSD.n3136 VSSD.n1060 34.6358
R10525 VSSD.n3132 VSSD.n1068 34.6358
R10526 VSSD.n3128 VSSD.n1068 34.6358
R10527 VSSD.n3128 VSSD.n3127 34.6358
R10528 VSSD.n3122 VSSD.n3121 34.6358
R10529 VSSD.n3106 VSSD.n3105 34.6358
R10530 VSSD.n3105 VSSD.n3104 34.6358
R10531 VSSD.n3104 VSSD.n3065 34.6358
R10532 VSSD.n3100 VSSD.n3065 34.6358
R10533 VSSD.n3100 VSSD.n3099 34.6358
R10534 VSSD.n3097 VSSD.n3069 34.6358
R10535 VSSD.n3093 VSSD.n3069 34.6358
R10536 VSSD.n3093 VSSD.n3092 34.6358
R10537 VSSD.n3092 VSSD.n3091 34.6358
R10538 VSSD.n3088 VSSD.n3087 34.6358
R10539 VSSD.n3087 VSSD.n3086 34.6358
R10540 VSSD.n2658 VSSD.n2644 34.6358
R10541 VSSD.n2589 VSSD.n2588 34.6358
R10542 VSSD.n2596 VSSD.n2595 34.6358
R10543 VSSD.n2596 VSSD.n2540 34.6358
R10544 VSSD.n2600 VSSD.n2540 34.6358
R10545 VSSD.n2606 VSSD.n2538 34.6358
R10546 VSSD.n2610 VSSD.n2538 34.6358
R10547 VSSD.n2611 VSSD.n2610 34.6358
R10548 VSSD.n2612 VSSD.n2611 34.6358
R10549 VSSD.n2692 VSSD.n1371 34.6358
R10550 VSSD.n2813 VSSD.n2812 34.6358
R10551 VSSD.n2804 VSSD.n2803 34.6358
R10552 VSSD.n2339 VSSD.n2335 34.6358
R10553 VSSD.n2343 VSSD.n2312 34.6358
R10554 VSSD.n2344 VSSD.n2343 34.6358
R10555 VSSD.n2344 VSSD.n1425 34.6358
R10556 VSSD.n2355 VSSD.n1425 34.6358
R10557 VSSD.n2361 VSSD.n1423 34.6358
R10558 VSSD.n1411 VSSD.n1407 34.6358
R10559 VSSD.n2484 VSSD.n1394 34.6358
R10560 VSSD.n2484 VSSD.n2483 34.6358
R10561 VSSD.n2483 VSSD.n2482 34.6358
R10562 VSSD.n2499 VSSD.n1389 34.6358
R10563 VSSD.n2495 VSSD.n1389 34.6358
R10564 VSSD.n2495 VSSD.n2494 34.6358
R10565 VSSD.n2503 VSSD.n2502 34.6358
R10566 VSSD.n1560 VSSD.n1498 34.6358
R10567 VSSD.n1549 VSSD.n1548 34.6358
R10568 VSSD.n1548 VSSD.n1547 34.6358
R10569 VSSD.n1544 VSSD.n1543 34.6358
R10570 VSSD.n1541 VSSD.n1506 34.6358
R10571 VSSD.n1537 VSSD.n1506 34.6358
R10572 VSSD.n1537 VSSD.n1536 34.6358
R10573 VSSD.n2007 VSSD.n1463 34.6358
R10574 VSSD.n2008 VSSD.n2007 34.6358
R10575 VSSD.n2009 VSSD.n2008 34.6358
R10576 VSSD.n2003 VSSD.n2000 34.6358
R10577 VSSD.n1994 VSSD.n1466 34.6358
R10578 VSSD.n1998 VSSD.n1466 34.6358
R10579 VSSD.n1992 VSSD.n1991 34.6358
R10580 VSSD.n1971 VSSD.n1969 34.6358
R10581 VSSD.n2097 VSSD.n2096 34.6358
R10582 VSSD.n2093 VSSD.n2092 34.6358
R10583 VSSD.n2089 VSSD.n2056 34.6358
R10584 VSSD.n2235 VSSD.n2129 34.6358
R10585 VSSD.n2203 VSSD.n2148 34.6358
R10586 VSSD.n2199 VSSD.n2148 34.6358
R10587 VSSD.n2199 VSSD.n2198 34.6358
R10588 VSSD.n2196 VSSD.n2151 34.6358
R10589 VSSD.n2192 VSSD.n2191 34.6358
R10590 VSSD.n2191 VSSD.n2190 34.6358
R10591 VSSD.n2187 VSSD.n2186 34.6358
R10592 VSSD.n1781 VSSD.n1690 34.6358
R10593 VSSD.n1785 VSSD.n1784 34.6358
R10594 VSSD.n1790 VSSD.n1789 34.6358
R10595 VSSD.n1803 VSSD.n1672 34.6358
R10596 VSSD.n1685 VSSD.n1672 34.6358
R10597 VSSD.n1793 VSSD.n1685 34.6358
R10598 VSSD.n1806 VSSD.n1670 34.6358
R10599 VSSD.n1812 VSSD.n1811 34.6358
R10600 VSSD.n1856 VSSD.n1855 34.6358
R10601 VSSD.n1871 VSSD.n1632 34.6358
R10602 VSSD.n1867 VSSD.n1632 34.6358
R10603 VSSD.n1867 VSSD.n1866 34.6358
R10604 VSSD.n1866 VSSD.n1865 34.6358
R10605 VSSD.n1875 VSSD.n1628 34.6358
R10606 VSSD.n1875 VSSD.n1874 34.6358
R10607 VSSD.n1888 VSSD.n1887 34.6358
R10608 VSSD.n1887 VSSD.n1626 34.6358
R10609 VSSD.n458 VSSD.n158 34.6358
R10610 VSSD.n454 VSSD.n158 34.6358
R10611 VSSD.n454 VSSD.n453 34.6358
R10612 VSSD.n453 VSSD.n452 34.6358
R10613 VSSD.n469 VSSD.n468 34.6358
R10614 VSSD.n468 VSSD.n156 34.6358
R10615 VSSD.n464 VSSD.n156 34.6358
R10616 VSSD.n482 VSSD.n142 34.6358
R10617 VSSD.n412 VSSD.n411 34.6358
R10618 VSSD.n408 VSSD.n407 34.6358
R10619 VSSD.n407 VSSD.n406 34.6358
R10620 VSSD.n406 VSSD.n189 34.6358
R10621 VSSD.n402 VSSD.n189 34.6358
R10622 VSSD.n398 VSSD.n193 34.6358
R10623 VSSD.n394 VSSD.n193 34.6358
R10624 VSSD.n394 VSSD.n393 34.6358
R10625 VSSD.n393 VSSD.n392 34.6358
R10626 VSSD.n389 VSSD.n388 34.6358
R10627 VSSD.n355 VSSD.n354 34.6358
R10628 VSSD.n354 VSSD.n220 34.6358
R10629 VSSD.n350 VSSD.n220 34.6358
R10630 VSSD.n348 VSSD.n347 34.6358
R10631 VSSD.n489 VSSD.n133 34.6358
R10632 VSSD.n3689 VSSD.n3688 34.6358
R10633 VSSD.n3696 VSSD.n3695 34.6358
R10634 VSSD.n3696 VSSD.n23 34.6358
R10635 VSSD.n3708 VSSD.n23 34.6358
R10636 VSSD.n3717 VSSD.n21 34.6358
R10637 VSSD.n3732 VSSD.n3729 34.6358
R10638 VSSD.n3736 VSSD.n15 34.6358
R10639 VSSD.n652 VSSD.t1908 34.2973
R10640 VSSD.n781 VSSD.t1914 34.2973
R10641 VSSD.n1277 VSSD.t1892 34.2973
R10642 VSSD.n3312 VSSD.t1882 34.2973
R10643 VSSD.n1127 VSSD.t1947 34.2973
R10644 VSSD.n2222 VSSD.t1854 34.2973
R10645 VSSD.n2117 VSSD.t1929 34.2973
R10646 VSSD.n1822 VSSD.t1901 34.2973
R10647 VSSD.n179 VSSD.t1937 34.2973
R10648 VSSD.n1265 VSSD.n1239 33.8829
R10649 VSSD.n2939 VSSD.n2938 33.8829
R10650 VSSD.n1407 VSSD.n1400 33.8829
R10651 VSSD.n2494 VSSD.n1391 33.8829
R10652 VSSD.n1530 VSSD.n1529 33.8829
R10653 VSSD.n2017 VSSD.n2016 33.8829
R10654 VSSD.n2121 VSSD.n2118 33.8829
R10655 VSSD.n2210 VSSD.n2145 33.8829
R10656 VSSD.t786 VSSD.t1096 33.717
R10657 VSSD.t1576 VSSD.t1818 33.717
R10658 VSSD.t614 VSSD.t1777 33.717
R10659 VSSD.t971 VSSD.t1720 33.717
R10660 VSSD.t431 VSSD.t636 33.717
R10661 VSSD.t197 VSSD.t973 33.717
R10662 VSSD.t133 VSSD.t728 33.717
R10663 VSSD.t832 VSSD.t913 33.717
R10664 VSSD.t827 VSSD.t396 33.717
R10665 VSSD.t1654 VSSD 33.717
R10666 VSSD.t1121 VSSD.t1755 33.717
R10667 VSSD.t1118 VSSD.t473 33.717
R10668 VSSD.n1975 VSSD.n1974 33.1299
R10669 VSSD.n3190 VSSD.n1048 33.1299
R10670 VSSD.n2212 VSSD.n2141 32.7534
R10671 VSSD.n2662 VSSD.n2661 32.377
R10672 VSSD.n2367 VSSD.n2366 32.377
R10673 VSSD.n2508 VSSD.n1384 32.377
R10674 VSSD.n1491 VSSD.n1479 32.377
R10675 VSSD.n1979 VSSD.n1962 32.377
R10676 VSSD.n1974 VSSD.n1963 32.377
R10677 VSSD.n2100 VSSD.n2048 32.377
R10678 VSSD.n2180 VSSD.n2179 32.377
R10679 VSSD.n2085 VSSD.n2084 31.624
R10680 VSSD.n968 VSSD.n838 29.7417
R10681 VSSD.n975 VSSD.n974 29.7417
R10682 VSSD.n3342 VSSD.n527 29.7417
R10683 VSSD.n908 VSSD.n881 29.7417
R10684 VSSD.n1200 VSSD.n1199 29.7417
R10685 VSSD.n3110 VSSD.n3063 29.7417
R10686 VSSD.n2654 VSSD.n2653 29.7417
R10687 VSSD.n2478 VSSD.n1396 29.7417
R10688 VSSD.n2489 VSSD.n2488 29.7417
R10689 VSSD.n1535 VSSD.n1534 29.7417
R10690 VSSD.n2013 VSSD.n1461 29.7417
R10691 VSSD.n2256 VSSD.n2255 29.7417
R10692 VSSD.n2205 VSSD.n2204 29.7417
R10693 VSSD.n1785 VSSD.n1686 29.7417
R10694 VSSD.n1811 VSSD.n1810 29.7417
R10695 VSSD.n1861 VSSD.n1860 29.7417
R10696 VSSD.n3163 VSSD.n1035 28.9887
R10697 VSSD.n2836 VSSD.n2835 28.9887
R10698 VSSD.n2817 VSSD.n2816 28.9887
R10699 VSSD.n2934 VSSD.n2933 27.8593
R10700 VSSD.n2236 VSSD.n2235 27.4829
R10701 VSSD.n1883 VSSD.n1626 27.4829
R10702 VSSD.n239 VSSD.n226 27.4829
R10703 VSSD.n825 VSSD.n752 27.4829
R10704 VSSD.n3213 VSSD.n1042 27.1064
R10705 VSSD.n2929 VSSD.n2928 27.1064
R10706 VSSD.n1534 VSSD.n1509 27.1064
R10707 VSSD.n2014 VSSD.n2013 27.1064
R10708 VSSD.n2277 VSSD.n2108 27.1064
R10709 VSSD.n2206 VSSD.n2205 27.1064
R10710 VSSD.n356 VSSD.n355 27.1064
R10711 VSSD.n2873 VSSD.n2872 26.7039
R10712 VSSD.n956 VSSD.n857 26.6009
R10713 VSSD.n2452 VSSD.n2385 26.6009
R10714 VSSD.n2077 VSSD.n2066 26.6009
R10715 VSSD.n3655 VSSD.n3592 26.6009
R10716 VSSD.n3738 VSSD.n3736 26.6009
R10717 VSSD.n2281 VSSD.n2280 26.314
R10718 VSSD.n3356 VSSD.n3355 26.314
R10719 VSSD.n2929 VSSD.n2927 26.314
R10720 VSSD.n3191 VSSD.n3190 25.977
R10721 VSSD.n2962 VSSD.n2961 25.977
R10722 VSSD.n2808 VSSD.n1345 25.977
R10723 VSSD.n987 VSSD.n828 25.7355
R10724 VSSD.n980 VSSD.n979 25.7355
R10725 VSSD.n806 VSSD.n771 25.7355
R10726 VSSD.n3404 VSSD.n132 25.7355
R10727 VSSD.n2869 VSSD.n2862 25.6926
R10728 VSSD.n2832 VSSD.n2831 25.6926
R10729 VSSD.n2803 VSSD.n1347 25.6926
R10730 VSSD.n2330 VSSD.n2314 25.6926
R10731 VSSD.n2372 VSSD.n2371 25.6926
R10732 VSSD.n2464 VSSD.n1411 25.6926
R10733 VSSD.n2277 VSSD.n2276 25.6926
R10734 VSSD.n1777 VSSD.n1690 25.6926
R10735 VSSD.n1615 VSSD.n1598 25.6926
R10736 VSSD.n3206 VSSD.n3205 25.6005
R10737 VSSD.n2100 VSSD.n2099 25.6005
R10738 VSSD.t1571 VSSD.t338 25.2879
R10739 VSSD.t882 VSSD.t108 25.2879
R10740 VSSD VSSD.t1666 25.2879
R10741 VSSD.t1738 VSSD.t26 25.2879
R10742 VSSD.t30 VSSD.t1768 25.2879
R10743 VSSD.n3118 VSSD.n3117 25.224
R10744 VSSD.n2651 VSSD.n2649 25.224
R10745 VSSD.n2649 VSSD.n1322 25.224
R10746 VSSD.n488 VSSD.n487 25.224
R10747 VSSD.n2216 VSSD.n2215 24.9894
R10748 VSSD.n2262 VSSD.n2118 24.9894
R10749 VSSD.n1816 VSSD.n1815 24.9894
R10750 VSSD.n1043 VSSD.t649 24.9236
R10751 VSSD.n1043 VSSD.t1710 24.9236
R10752 VSSD.n3185 VSSD.t1015 24.9236
R10753 VSSD.n3185 VSSD.t1065 24.9236
R10754 VSSD.n1047 VSSD.t1011 24.9236
R10755 VSSD.n1047 VSSD.t547 24.9236
R10756 VSSD.n1046 VSSD.t1013 24.9236
R10757 VSSD.n1046 VSSD.t1067 24.9236
R10758 VSSD.n1279 VSSD.t566 24.9236
R10759 VSSD.n1279 VSSD.t381 24.9236
R10760 VSSD.n1238 VSSD.t1630 24.9236
R10761 VSSD.n1238 VSSD.t1182 24.9236
R10762 VSSD.n1243 VSSD.t1634 24.9236
R10763 VSSD.n1243 VSSD.t1180 24.9236
R10764 VSSD.n1241 VSSD.t1632 24.9236
R10765 VSSD.n1241 VSSD.t1628 24.9236
R10766 VSSD.n1236 VSSD.t421 24.9236
R10767 VSSD.n1236 VSSD.t1178 24.9236
R10768 VSSD.n1113 VSSD.t1104 24.9236
R10769 VSSD.n1113 VSSD.t1100 24.9236
R10770 VSSD.n1112 VSSD.t1102 24.9236
R10771 VSSD.n1112 VSSD.t846 24.9236
R10772 VSSD.n1100 VSSD.t848 24.9236
R10773 VSSD.n1100 VSSD.t757 24.9236
R10774 VSSD.n2952 VSSD.t1832 24.9236
R10775 VSSD.n2952 VSSD.t759 24.9236
R10776 VSSD.n1097 VSSD.t1828 24.9236
R10777 VSSD.n1097 VSSD.t755 24.9236
R10778 VSSD.n1331 VSSD.t1586 24.9236
R10779 VSSD.n1331 VSSD.t391 24.9236
R10780 VSSD.n1335 VSSD.t393 24.9236
R10781 VSSD.n1335 VSSD.t150 24.9236
R10782 VSSD.n1336 VSSD.t1093 24.9236
R10783 VSSD.n1336 VSSD.t105 24.9236
R10784 VSSD.n1341 VSSD.t910 24.9236
R10785 VSSD.n1341 VSSD.t107 24.9236
R10786 VSSD.n1344 VSSD.t912 24.9236
R10787 VSSD.n1344 VSSD.t152 24.9236
R10788 VSSD.n820 VSSD.n819 24.8476
R10789 VSSD.n3351 VSSD.n3350 24.8476
R10790 VSSD.n931 VSSD.n870 24.8476
R10791 VSSD.n1304 VSSD.n1137 24.8476
R10792 VSSD.n2968 VSSD.n1092 24.8476
R10793 VSSD.n2996 VSSD.n2995 24.8476
R10794 VSSD.n3121 VSSD.n3120 24.8476
R10795 VSSD.n3086 VSSD.n3075 24.8476
R10796 VSSD.n2588 VSSD.n2587 24.8476
R10797 VSSD.n2365 VSSD.n1423 24.8476
R10798 VSSD.n2371 VSSD.n1421 24.8476
R10799 VSSD.n2507 VSSD.n1385 24.8476
R10800 VSSD.n1562 VSSD.n1496 24.8476
R10801 VSSD.n1980 VSSD.n1961 24.8476
R10802 VSSD.n2257 VSSD.n2256 24.8476
R10803 VSSD.n2254 VSSD.n2124 24.8476
R10804 VSSD.n2184 VSSD.n2159 24.8476
R10805 VSSD.n1782 VSSD.n1781 24.8476
R10806 VSSD.n1815 VSSD.n1666 24.8476
R10807 VSSD.n1879 VSSD.n1628 24.8476
R10808 VSSD.n483 VSSD.n482 24.8476
R10809 VSSD.n344 VSSD.n343 24.8476
R10810 VSSD.n3688 VSSD.n37 24.8476
R10811 VSSD.n3718 VSSD.n3717 24.8476
R10812 VSSD.n3732 VSSD.n3731 24.8476
R10813 VSSD.n1625 VSSD.n1624 24.8081
R10814 VSSD.n2518 VSSD.n1382 24.8035
R10815 VSSD.n3217 VSSD.n1042 24.8035
R10816 VSSD.n1205 VSSD.n1204 24.0946
R10817 VSSD.n2960 VSSD.n2959 24.0946
R10818 VSSD.n2177 VSSD.n2176 23.8103
R10819 VSSD.n3116 VSSD.n3059 23.7181
R10820 VSSD.n563 VSSD.n560 23.7181
R10821 VSSD.n670 VSSD.n560 23.7181
R10822 VSSD.n3193 VSSD.n3184 23.7181
R10823 VSSD.n2865 VSSD.n2862 23.7181
R10824 VSSD.n3112 VSSD.n3059 23.7181
R10825 VSSD.n1969 VSSD.n1966 23.7181
R10826 VSSD.n2078 VSSD.n2077 23.7181
R10827 VSSD.n1602 VSSD.n1598 23.7181
R10828 VSSD.n3408 VSSD.n132 23.7181
R10829 VSSD.n3656 VSSD.n3655 23.7181
R10830 VSSD.n440 VSSD.n162 23.7181
R10831 VSSD.n362 VSSD.n214 23.7181
R10832 VSSD.n136 VSSD.n133 23.7181
R10833 VSSD.n3670 VSSD.n3669 23.7181
R10834 VSSD.n746 VSSD.n743 23.2027
R10835 VSSD.n999 VSSD.n743 22.9652
R10836 VSSD.n812 VSSD.n811 22.9652
R10837 VSSD.n821 VSSD.n752 22.9652
R10838 VSSD.n761 VSSD.n527 22.9652
R10839 VSSD.n932 VSSD.n931 22.9652
R10840 VSSD.n908 VSSD.n907 22.9652
R10841 VSSD.n1200 VSSD.n1157 22.9652
R10842 VSSD.n1303 VSSD.n1138 22.9652
R10843 VSSD.n2967 VSSD.n2966 22.9652
R10844 VSSD.n3007 VSSD.n1081 22.9652
R10845 VSSD.n3111 VSSD.n3110 22.9652
R10846 VSSD.n3082 VSSD.n3081 22.9652
R10847 VSSD.n2335 VSSD.n2334 22.9652
R10848 VSSD.n1529 VSSD.n1528 22.9652
R10849 VSSD.n2453 VSSD.n2452 22.9652
R10850 VSSD.n2017 VSSD.n1458 22.9652
R10851 VSSD.n2237 VSSD.n2236 22.9652
R10852 VSSD.n2211 VSSD.n2210 22.9652
R10853 VSSD.n1860 VSSD.n1638 22.9652
R10854 VSSD.n413 VSSD.n412 22.9652
R10855 VSSD.n388 VSSD.n200 22.9652
R10856 VSSD.n361 VSSD.n360 22.9652
R10857 VSSD.n342 VSSD.n226 22.9652
R10858 VSSD.n3684 VSSD.n3683 22.9652
R10859 VSSD.n3719 VSSD.n19 22.9652
R10860 VSSD.n2690 VSSD.n2632 22.5887
R10861 VSSD.n2686 VSSD.n2632 22.5887
R10862 VSSD.n2080 VSSD.n2079 22.5887
R10863 VSSD.n2079 VSSD.n2078 22.5887
R10864 VSSD.n3042 VSSD.n3041 22.5419
R10865 VSSD.n2631 VSSD.t959 22.3257
R10866 VSSD.n1387 VSSD.t1800 22.3257
R10867 VSSD.n1490 VSSD.n1489 22.2123
R10868 VSSD.n2938 VSSD.n1101 21.8358
R10869 VSSD.n2816 VSSD.n1337 21.8358
R10870 VSSD.n1001 VSSD.n742 21.4593
R10871 VSSD.n811 VSSD.n771 21.4593
R10872 VSSD.n821 VSSD.n820 21.4593
R10873 VSSD.n762 VSSD.n761 21.4593
R10874 VSSD.n3352 VSSD.n3351 21.4593
R10875 VSSD.n907 VSSD.n905 21.4593
R10876 VSSD.n1204 VSSD.n1157 21.4593
R10877 VSSD.n1304 VSSD.n1303 21.4593
R10878 VSSD.n2968 VSSD.n2967 21.4593
R10879 VSSD.n2995 VSSD.n1081 21.4593
R10880 VSSD.n3112 VSSD.n3111 21.4593
R10881 VSSD.n3082 VSSD.n3075 21.4593
R10882 VSSD.n2620 VSSD.n1371 21.4593
R10883 VSSD.n2334 VSSD.n2314 21.4593
R10884 VSSD.n2366 VSSD.n2365 21.4593
R10885 VSSD.n2508 VSSD.n2507 21.4593
R10886 VSSD.n1496 VSSD.n1479 21.4593
R10887 VSSD.n1980 VSSD.n1979 21.4593
R10888 VSSD.n2237 VSSD.n2124 21.4593
R10889 VSSD.n2212 VSSD.n2211 21.4593
R10890 VSSD.n2180 VSSD.n2159 21.4593
R10891 VSSD.n1856 VSSD.n1638 21.4593
R10892 VSSD.n1880 VSSD.n1879 21.4593
R10893 VSSD.n445 VSSD.n162 21.4593
R10894 VSSD.n376 VSSD.n209 21.4593
R10895 VSSD.n376 VSSD.n375 21.4593
R10896 VSSD.n362 VSSD.n361 21.4593
R10897 VSSD.n343 VSSD.n342 21.4593
R10898 VSSD.n3670 VSSD.n43 21.4593
R10899 VSSD.n3684 VSSD.n37 21.4593
R10900 VSSD.n3719 VSSD.n3718 21.4593
R10901 VSSD.n3729 VSSD.n17 21.4593
R10902 VSSD.n2836 VSSD.n1322 20.7064
R10903 VSSD.n825 VSSD.n751 20.3299
R10904 VSSD.n3352 VSSD.n524 20.3299
R10905 VSSD.n2478 VSSD.n2477 20.3299
R10906 VSSD.n2490 VSSD.n2489 20.3299
R10907 VSSD.n360 VSSD.n218 20.3299
R10908 VSSD.n3723 VSSD.n19 20.3299
R10909 VSSD.n849 VSSD.n847 19.577
R10910 VSSD.n835 VSSD.n832 19.577
R10911 VSSD.n1256 VSSD.n1255 19.577
R10912 VSSD.n2680 VSSD.n2634 19.577
R10913 VSSD.n2660 VSSD.n2659 19.2005
R10914 VSSD.n2105 VSSD.n2104 19.2005
R10915 VSSD.n3207 VSSD.n3206 18.824
R10916 VSSD.n3212 VSSD.n1044 18.824
R10917 VSSD.n2666 VSSD.n2640 18.824
R10918 VSSD.n2692 VSSD.n2691 18.824
R10919 VSSD.n1299 VSSD.n1138 18.5826
R10920 VSSD.n3683 VSSD.n3682 18.5397
R10921 VSSD.n2804 VSSD.n1345 18.4476
R10922 VSSD.n700 VSSD.n696 18.2791
R10923 VSSD.n3279 VSSD.n3278 18.2791
R10924 VSSD.n2744 VSSD.n2743 18.2791
R10925 VSSD.n1743 VSSD.n1742 18.2791
R10926 VSSD.n1920 VSSD.n1919 18.2791
R10927 VSSD.n3445 VSSD.n3444 18.2791
R10928 VSSD.n3502 VSSD.n3500 18.2791
R10929 VSSD.n3571 VSSD.n3570 18.2791
R10930 VSSD.n3635 VSSD.n3634 18.2791
R10931 VSSD.n1247 VSSD.n1244 18.0711
R10932 VSSD.n3037 VSSD.n3036 18.0711
R10933 VSSD.n2676 VSSD.n2675 18.0711
R10934 VSSD.n2618 VSSD.n2616 18.0711
R10935 VSSD.n2084 VSSD.n2083 18.0711
R10936 VSSD.n448 VSSD.n447 18.0711
R10937 VSSD.n3416 VSSD.n3415 17.7007
R10938 VSSD.n3481 VSSD.n3480 17.7007
R10939 VSSD.n3542 VSSD.n3541 17.7007
R10940 VSSD.n3346 VSSD.n3345 17.6946
R10941 VSSD.n876 VSSD.n873 17.6946
R10942 VSSD.n1178 VSSD.n1177 17.6946
R10943 VSSD.n3126 VSSD.n3125 17.6946
R10944 VSSD.n3122 VSSD.n1072 17.6946
R10945 VSSD.n3088 VSSD.n3073 17.6946
R10946 VSSD.n2589 VSSD.n2543 17.6946
R10947 VSSD.n2594 VSSD.n2592 17.6946
R10948 VSSD.n2358 VSSD.n2357 17.6946
R10949 VSSD.n2502 VSSD.n2501 17.6946
R10950 VSSD.n1562 VSSD.n1561 17.6946
R10951 VSSD.n1501 VSSD.n1498 17.6946
R10952 VSSD.n1993 VSSD.n1992 17.6946
R10953 VSSD.n1961 VSSD.n1470 17.6946
R10954 VSSD.n2187 VSSD.n2156 17.6946
R10955 VSSD.n2185 VSSD.n2184 17.6946
R10956 VSSD.n472 VSSD.n471 17.6946
R10957 VSSD.n155 VSSD.n142 17.6946
R10958 VSSD.n349 VSSD.n348 17.6946
R10959 VSSD.n3692 VSSD.n35 17.6946
R10960 VSSD.n3713 VSSD.n3710 17.6946
R10961 VSSD.n2790 VSSD.n2789 17.6577
R10962 VSSD.n1947 VSSD.n1575 17.6577
R10963 VSSD.n3615 VSSD.n3614 17.4137
R10964 VSSD.n188 VSSD.n185 17.3181
R10965 VSSD.n198 VSSD.n196 17.3181
R10966 VSSD.n3164 VSSD.n3163 17.1605
R10967 VSSD.n2878 VSSD.n2859 16.9936
R10968 VSSD.n2879 VSSD.n2878 16.9936
R10969 VSSD.n1832 VSSD.n1656 16.9936
R10970 VSSD.n1835 VSSD.n1832 16.9936
R10971 VSSD.n2906 VSSD.n2905 16.9545
R10972 VSSD.t157 VSSD.t1752 16.8587
R10973 VSSD.t1542 VSSD.t565 16.8587
R10974 VSSD.t304 VSSD.t1558 16.8587
R10975 VSSD.t1563 VSSD.t1762 16.8587
R10976 VSSD.t1172 VSSD.t1381 16.8587
R10977 VSSD.t986 VSSD 16.8587
R10978 VSSD.t313 VSSD.t1204 16.8587
R10979 VSSD VSSD.t173 16.8587
R10980 VSSD.n800 VSSD.n774 16.7924
R10981 VSSD.n933 VSSD.n932 16.5652
R10982 VSSD.n1264 VSSD.n1263 16.5652
R10983 VSSD.n3081 VSSD.n3080 16.5652
R10984 VSSD.n2820 VSSD.n2819 16.5652
R10985 VSSD.n1485 VSSD.n1480 16.5652
R10986 VSSD.n3725 VSSD.n3724 16.5652
R10987 VSSD.n2654 VSSD.n2644 16.1887
R10988 VSSD.n2686 VSSD.n2684 16.1887
R10989 VSSD.n291 VSSD.n290 16.0722
R10990 VSSD.n989 VSSD.n988 15.9044
R10991 VSSD.n1265 VSSD.n1264 15.8123
R10992 VSSD.n2663 VSSD.n2640 15.8123
R10993 VSSD.n2583 VSSD.n2582 15.8123
R10994 VSSD.n2092 VSSD.n2091 15.8123
R10995 VSSD.n905 VSSD.n883 15.6771
R10996 VSSD.n1855 VSSD.n1639 15.6771
R10997 VSSD.n3669 VSSD.n44 15.3963
R10998 VSSD.n934 VSSD.n933 15.3963
R10999 VSSD.n3473 VSSD.n95 15.3963
R11000 VSSD.n3534 VSSD.n72 15.3963
R11001 VSSD.n3656 VSSD.n47 15.3963
R11002 VSSD.n3213 VSSD.n3212 15.0593
R11003 VSSD.n1144 VSSD.n1143 14.8179
R11004 VSSD.n3409 VSSD.n3408 14.8179
R11005 VSSD.n3474 VSSD.n3473 14.8179
R11006 VSSD.n3535 VSSD.n3534 14.8179
R11007 VSSD.n496 VSSD.n495 14.775
R11008 VSSD.n2824 VSSD.n1329 14.775
R11009 VSSD.n2563 VSSD.n2562 14.775
R11010 VSSD.n2169 VSSD.n2168 14.775
R11011 VSSD.n366 VSSD.n214 14.775
R11012 VSSD.n974 VSSD.n836 14.6829
R11013 VSSD.n969 VSSD.n968 14.6829
R11014 VSSD.n815 VSSD.n769 14.6829
R11015 VSSD.n3343 VSSD.n3342 14.6829
R11016 VSSD.n912 VSSD.n881 14.6829
R11017 VSSD.n1199 VSSD.n1198 14.6829
R11018 VSSD.n3035 VSSD.n1059 14.6829
R11019 VSSD.n3106 VSSD.n3063 14.6829
R11020 VSSD.n2612 VSSD.n2536 14.6829
R11021 VSSD.n2488 VSSD.n1394 14.6829
R11022 VSSD.n2482 VSSD.n1396 14.6829
R11023 VSSD.n1536 VSSD.n1535 14.6829
R11024 VSSD.n2009 VSSD.n1461 14.6829
R11025 VSSD.n2255 VSSD.n2254 14.6829
R11026 VSSD.n2204 VSSD.n2203 14.6829
R11027 VSSD.n1789 VSSD.n1686 14.6829
R11028 VSSD.n1810 VSSD.n1670 14.6829
R11029 VSSD.n1862 VSSD.n1861 14.6829
R11030 VSSD.n452 VSSD.n160 14.6829
R11031 VSSD.n311 VSSD.n310 14.5992
R11032 VSSD.n2321 VSSD.n1416 14.3064
R11033 VSSD.n2453 VSSD.n1417 14.3064
R11034 VSSD.n2477 VSSD.n2476 14.3064
R11035 VSSD.n2491 VSSD.n2490 14.3064
R11036 VSSD.n357 VSSD.n218 14.3064
R11037 VSSD.n856 VSSD.n847 14.3064
R11038 VSSD.n979 VSSD.n832 14.3064
R11039 VSSD.n762 VSSD.n751 14.3064
R11040 VSSD.n2835 VSSD.n1325 14.3064
R11041 VSSD.n2337 VSSD.n2312 14.3064
R11042 VSSD.n1874 VSSD.n1873 14.3064
R11043 VSSD.n271 VSSD.n270 14.2735
R11044 VSSD.n3306 VSSD.n3305 14.0717
R11045 VSSD.n3255 VSSD.n3254 14.0503
R11046 VSSD.n2720 VSSD.n2719 14.0503
R11047 VSSD.n2407 VSSD.n2406 14.0503
R11048 VSSD.n1719 VSSD.n1718 14.0503
R11049 VSSD.n3790 VSSD.n3787 14.0503
R11050 VSSD.n2322 VSSD.n2321 14.022
R11051 VSSD.n2380 VSSD.n1417 14.022
R11052 VSSD.n375 VSSD.n374 14.022
R11053 VSSD.n2661 VSSD.n2660 13.9299
R11054 VSSD.n2962 VSSD.n1094 13.5534
R11055 VSSD.n2671 VSSD.n2670 13.5534
R11056 VSSD.n2085 VSSD.n2059 13.5534
R11057 VSSD.n1326 VSSD.n1325 13.177
R11058 VSSD.n3725 VSSD.n17 13.177
R11059 VSSD.n2767 VSSD.n2766 13.1375
R11060 VSSD.n670 VSSD.n559 12.8005
R11061 VSSD.n893 VSSD.n889 12.8005
R11062 VSSD.n815 VSSD.n814 12.8005
R11063 VSSD.n2951 VSSD.n1101 12.8005
R11064 VSSD.n2338 VSSD.n2337 12.8005
R11065 VSSD.n2105 VSSD.n1451 12.8005
R11066 VSSD.n1269 VSSD.n1268 12.7129
R11067 VSSD.n3020 VSSD.n3019 12.5161
R11068 VSSD.n2021 VSSD.n1458 12.5161
R11069 VSSD.n1766 VSSD.n1765 12.5161
R11070 VSSD.n2809 VSSD.n2808 12.424
R11071 VSSD.n3229 VSSD.n3228 12.1788
R11072 VSSD.n3157 VSSD.n3156 12.1788
R11073 VSSD.n524 VSSD.n521 12.0476
R11074 VSSD.n1340 VSSD.n1337 12.0476
R11075 VSSD.n2810 VSSD.n2809 12.0476
R11076 VSSD.n1489 VSSD.n1480 12.0476
R11077 VSSD.n2456 VSSD.n1416 12.0476
R11078 VSSD.n417 VSSD.n181 11.8129
R11079 VSSD.n3120 VSSD.n3119 11.6711
R11080 VSSD.n2587 VSSD.n2545 11.6711
R11081 VSSD.n2096 VSSD.n2052 11.6711
R11082 VSSD.n483 VSSD.n140 11.6711
R11083 VSSD.n413 VSSD.n181 11.6711
R11084 VSSD.n209 VSSD.n200 11.6711
R11085 VSSD.n1270 VSSD.n1269 11.4892
R11086 VSSD.n1255 VSSD.n1254 11.2946
R11087 VSSD.n2819 VSSD.n2818 11.2946
R11088 VSSD.n1281 VSSD.n1280 10.9719
R11089 VSSD.n3764 VSSD.n7 10.9181
R11090 VSSD.n3040 VSSD.n3039 10.7135
R11091 VSSD.n2582 VSSD.n2547 10.7135
R11092 VSSD.n440 VSSD.n439 10.7135
R11093 VSSD.n512 VSSD.n499 10.6521
R11094 VSSD.n3302 VSSD.n3301 10.5417
R11095 VSSD.n3039 VSSD.n3038 10.5417
R11096 VSSD.n2456 VSSD.n1415 10.5417
R11097 VSSD.n1873 VSSD.n1872 10.5417
R11098 VSSD.n568 VSSD.n559 10.4353
R11099 VSSD.n2430 VSSD.n2428 10.2976
R11100 VSSD.n988 VSSD.n987 9.78874
R11101 VSSD.n3305 VSSD.n1035 9.78874
R11102 VSSD.n1261 VSSD.n1244 9.78874
R11103 VSSD.n2959 VSSD.n2958 9.78874
R11104 VSSD.n3038 VSSD.n3037 9.78874
R11105 VSSD.n3036 VSSD.n3035 9.78874
R11106 VSSD.n3119 VSSD.n3118 9.78874
R11107 VSSD.n2583 VSSD.n2545 9.78874
R11108 VSSD.n2616 VSSD.n2536 9.78874
R11109 VSSD.n2620 VSSD.n2618 9.78874
R11110 VSSD.n2368 VSSD.n1421 9.78874
R11111 VSSD.n2090 VSSD.n2089 9.78874
R11112 VSSD.n2258 VSSD.n2257 9.78874
R11113 VSSD.n1872 VSSD.n1871 9.78874
R11114 VSSD.n447 VSSD.n445 9.78874
R11115 VSSD.n448 VSSD.n160 9.78874
R11116 VSSD.n487 VSSD.n140 9.78874
R11117 VSSD.n408 VSSD.n188 9.78874
R11118 VSSD.n392 VSSD.n196 9.78874
R11119 VSSD.n3731 VSSD.n15 9.78874
R11120 VSSD.n3400 VSSD 9.74003
R11121 VSSD.n3609 VSSD.n3608 9.71789
R11122 VSSD.n332 VSSD.n241 9.65974
R11123 VSSD.n2691 VSSD.n2690 9.41227
R11124 VSSD.n1388 VSSD.n1385 9.41227
R11125 VSSD.n907 VSSD.n882 9.3005
R11126 VSSD.n903 VSSD.n902 9.3005
R11127 VSSD.n900 VSSD.n884 9.3005
R11128 VSSD.n899 VSSD.n898 9.3005
R11129 VSSD.n897 VSSD.n896 9.3005
R11130 VSSD.n905 VSSD.n904 9.3005
R11131 VSSD.n909 VSSD.n908 9.3005
R11132 VSSD.n910 VSSD.n881 9.3005
R11133 VSSD.n912 VSSD.n911 9.3005
R11134 VSSD.n913 VSSD.n879 9.3005
R11135 VSSD.n916 VSSD.n915 9.3005
R11136 VSSD.n917 VSSD.n878 9.3005
R11137 VSSD.n919 VSSD.n918 9.3005
R11138 VSSD.n920 VSSD.n874 9.3005
R11139 VSSD.n923 VSSD.n922 9.3005
R11140 VSSD.n924 VSSD.n873 9.3005
R11141 VSSD.n926 VSSD.n925 9.3005
R11142 VSSD.n927 VSSD.n871 9.3005
R11143 VSSD.n929 VSSD.n928 9.3005
R11144 VSSD.n931 VSSD.n930 9.3005
R11145 VSSD.n932 VSSD.n868 9.3005
R11146 VSSD.n933 VSSD.n867 9.3005
R11147 VSSD.n934 VSSD.n865 9.3005
R11148 VSSD.n938 VSSD.n937 9.3005
R11149 VSSD.n940 VSSD.n939 9.3005
R11150 VSSD.n941 VSSD.n862 9.3005
R11151 VSSD.n945 VSSD.n944 9.3005
R11152 VSSD.n946 VSSD.n861 9.3005
R11153 VSSD.n948 VSSD.n947 9.3005
R11154 VSSD.n949 VSSD.n860 9.3005
R11155 VSSD.n951 VSSD.n950 9.3005
R11156 VSSD.n953 VSSD.n952 9.3005
R11157 VSSD.n954 VSSD.n845 9.3005
R11158 VSSD.n957 VSSD.n956 9.3005
R11159 VSSD.n497 VSSD.n496 9.3005
R11160 VSSD.n3388 VSSD.n498 9.3005
R11161 VSSD.n3386 VSSD.n3385 9.3005
R11162 VSSD.n3376 VSSD.n513 9.3005
R11163 VSSD.n3377 VSSD.n3376 9.3005
R11164 VSSD.n3374 VSSD.n3373 9.3005
R11165 VSSD.n3372 VSSD.n3371 9.3005
R11166 VSSD.n3369 VSSD.n515 9.3005
R11167 VSSD.n3368 VSSD.n3367 9.3005
R11168 VSSD.n3366 VSSD.n516 9.3005
R11169 VSSD.n3365 VSSD.n3364 9.3005
R11170 VSSD.n3361 VSSD.n517 9.3005
R11171 VSSD.n3360 VSSD.n3359 9.3005
R11172 VSSD.n3358 VSSD.n519 9.3005
R11173 VSSD.n3357 VSSD.n3356 9.3005
R11174 VSSD.n3355 VSSD.n3354 9.3005
R11175 VSSD.n3353 VSSD.n3352 9.3005
R11176 VSSD.n3351 VSSD.n522 9.3005
R11177 VSSD.n3350 VSSD.n3349 9.3005
R11178 VSSD.n3348 VSSD.n525 9.3005
R11179 VSSD.n3347 VSSD.n3346 9.3005
R11180 VSSD.n3343 VSSD.n526 9.3005
R11181 VSSD.n3342 VSSD.n3341 9.3005
R11182 VSSD.n528 VSSD.n527 9.3005
R11183 VSSD.n761 VSSD.n760 9.3005
R11184 VSSD.n763 VSSD.n762 9.3005
R11185 VSSD.n825 VSSD.n824 9.3005
R11186 VSSD.n823 VSSD.n752 9.3005
R11187 VSSD.n822 VSSD.n821 9.3005
R11188 VSSD.n820 VSSD.n768 9.3005
R11189 VSSD.n819 VSSD.n818 9.3005
R11190 VSSD.n817 VSSD.n769 9.3005
R11191 VSSD.n816 VSSD.n815 9.3005
R11192 VSSD.n812 VSSD.n770 9.3005
R11193 VSSD.n811 VSSD.n809 9.3005
R11194 VSSD.n808 VSSD.n771 9.3005
R11195 VSSD.n807 VSSD.n806 9.3005
R11196 VSSD.n804 VSSD.n772 9.3005
R11197 VSSD.n800 VSSD.n799 9.3005
R11198 VSSD.n798 VSSD.n774 9.3005
R11199 VSSD.n797 VSSD.n796 9.3005
R11200 VSSD.n795 VSSD.n775 9.3005
R11201 VSSD.n794 VSSD.n793 9.3005
R11202 VSSD.n792 VSSD.n777 9.3005
R11203 VSSD.n791 VSSD.n790 9.3005
R11204 VSSD.n779 VSSD.n739 9.3005
R11205 VSSD.n784 VSSD.n740 9.3005
R11206 VSSD.n1002 VSSD.n1001 9.3005
R11207 VSSD.n999 VSSD.n998 9.3005
R11208 VSSD.n997 VSSD.n743 9.3005
R11209 VSSD.n996 VSSD.n995 9.3005
R11210 VSSD.n993 VSSD.n745 9.3005
R11211 VSSD.n992 VSSD.n991 9.3005
R11212 VSSD.n990 VSSD.n989 9.3005
R11213 VSSD.n987 VSSD.n986 9.3005
R11214 VSSD.n985 VSSD.n828 9.3005
R11215 VSSD.n984 VSSD.n983 9.3005
R11216 VSSD.n980 VSSD.n829 9.3005
R11217 VSSD.n979 VSSD.n978 9.3005
R11218 VSSD.n977 VSSD.n976 9.3005
R11219 VSSD.n975 VSSD.n833 9.3005
R11220 VSSD.n974 VSSD.n973 9.3005
R11221 VSSD.n972 VSSD.n836 9.3005
R11222 VSSD.n971 VSSD.n970 9.3005
R11223 VSSD.n969 VSSD.n837 9.3005
R11224 VSSD.n968 VSSD.n967 9.3005
R11225 VSSD.n966 VSSD.n838 9.3005
R11226 VSSD.n851 VSSD.n850 9.3005
R11227 VSSD.n856 VSSD.n855 9.3005
R11228 VSSD.n857 VSSD.n844 9.3005
R11229 VSSD.n1145 VSSD.n1144 9.3005
R11230 VSSD.n1296 VSSD.n1146 9.3005
R11231 VSSD.n1300 VSSD.n1299 9.3005
R11232 VSSD.n1301 VSSD.n1138 9.3005
R11233 VSSD.n1303 VSSD.n1302 9.3005
R11234 VSSD.n1305 VSSD.n1304 9.3005
R11235 VSSD.n1167 VSSD.n1137 9.3005
R11236 VSSD.n1176 VSSD.n1175 9.3005
R11237 VSSD.n1177 VSSD.n1164 9.3005
R11238 VSSD.n1180 VSSD.n1179 9.3005
R11239 VSSD.n1181 VSSD.n1163 9.3005
R11240 VSSD.n1183 VSSD.n1182 9.3005
R11241 VSSD.n1184 VSSD.n1162 9.3005
R11242 VSSD.n1189 VSSD.n1188 9.3005
R11243 VSSD.n1190 VSSD.n1161 9.3005
R11244 VSSD.n1192 VSSD.n1191 9.3005
R11245 VSSD.n1193 VSSD.n1160 9.3005
R11246 VSSD.n1195 VSSD.n1194 9.3005
R11247 VSSD.n1196 VSSD.n1159 9.3005
R11248 VSSD.n1198 VSSD.n1197 9.3005
R11249 VSSD.n1199 VSSD.n1158 9.3005
R11250 VSSD.n1201 VSSD.n1200 9.3005
R11251 VSSD.n1202 VSSD.n1157 9.3005
R11252 VSSD.n1204 VSSD.n1203 9.3005
R11253 VSSD.n1205 VSSD.n1154 9.3005
R11254 VSSD.n1208 VSSD.n1207 9.3005
R11255 VSSD.n1214 VSSD.n1213 9.3005
R11256 VSSD.n1218 VSSD.n1217 9.3005
R11257 VSSD.n1219 VSSD.n1147 9.3005
R11258 VSSD.n1294 VSSD.n1293 9.3005
R11259 VSSD.n1291 VSSD.n1290 9.3005
R11260 VSSD.n1288 VSSD.n1230 9.3005
R11261 VSSD.n1286 VSSD.n1285 9.3005
R11262 VSSD.n1284 VSSD.n1231 9.3005
R11263 VSSD.n1283 VSSD.n1282 9.3005
R11264 VSSD.n1234 VSSD.n1232 9.3005
R11265 VSSD.n1273 VSSD.n1272 9.3005
R11266 VSSD.n1271 VSSD.n1270 9.3005
R11267 VSSD.n1268 VSSD.n1267 9.3005
R11268 VSSD.n1266 VSSD.n1265 9.3005
R11269 VSSD.n1262 VSSD.n1240 9.3005
R11270 VSSD.n1261 VSSD.n1260 9.3005
R11271 VSSD.n1259 VSSD.n1258 9.3005
R11272 VSSD.n1257 VSSD.n1245 9.3005
R11273 VSSD.n1254 VSSD.n1253 9.3005
R11274 VSSD.n1252 VSSD.n1018 9.3005
R11275 VSSD.n1250 VSSD.n1019 9.3005
R11276 VSSD.n3321 VSSD.n3320 9.3005
R11277 VSSD.n3318 VSSD.n3317 9.3005
R11278 VSSD.n3316 VSSD.n1024 9.3005
R11279 VSSD.n3315 VSSD.n3314 9.3005
R11280 VSSD.n1028 VSSD.n1025 9.3005
R11281 VSSD.n3309 VSSD.n3308 9.3005
R11282 VSSD.n3307 VSSD.n3306 9.3005
R11283 VSSD.n3305 VSSD.n1036 9.3005
R11284 VSSD.n3161 VSSD.n1035 9.3005
R11285 VSSD.n3163 VSSD.n3162 9.3005
R11286 VSSD.n3166 VSSD.n3165 9.3005
R11287 VSSD.n3168 VSSD.n3167 9.3005
R11288 VSSD.n3169 VSSD.n3159 9.3005
R11289 VSSD.n3172 VSSD.n3171 9.3005
R11290 VSSD.n3173 VSSD.n3158 9.3005
R11291 VSSD.n3175 VSSD.n3174 9.3005
R11292 VSSD.n3177 VSSD.n3155 9.3005
R11293 VSSD.n3181 VSSD.n3180 9.3005
R11294 VSSD.n3184 VSSD.n3182 9.3005
R11295 VSSD.n3184 VSSD.n3183 9.3005
R11296 VSSD.n3194 VSSD.n3193 9.3005
R11297 VSSD.n3190 VSSD.n3189 9.3005
R11298 VSSD.n3204 VSSD.n3203 9.3005
R11299 VSSD.n3206 VSSD.n1045 9.3005
R11300 VSSD.n3209 VSSD.n3208 9.3005
R11301 VSSD.n3210 VSSD.n1044 9.3005
R11302 VSSD.n3212 VSSD.n3211 9.3005
R11303 VSSD.n3214 VSSD.n3213 9.3005
R11304 VSSD.n3215 VSSD.n1042 9.3005
R11305 VSSD.n3217 VSSD.n3216 9.3005
R11306 VSSD.n3219 VSSD.n1041 9.3005
R11307 VSSD.n3221 VSSD.n3220 9.3005
R11308 VSSD.n3222 VSSD.n1040 9.3005
R11309 VSSD.n3225 VSSD.n3224 9.3005
R11310 VSSD.n3223 VSSD.n1039 9.3005
R11311 VSSD.n3302 VSSD.n1038 9.3005
R11312 VSSD.n3302 VSSD.n1037 9.3005
R11313 VSSD.n3300 VSSD.n3299 9.3005
R11314 VSSD.n3298 VSSD.n3297 9.3005
R11315 VSSD.n3296 VSSD.n3234 9.3005
R11316 VSSD.n3294 VSSD.n3293 9.3005
R11317 VSSD.n3292 VSSD.n3236 9.3005
R11318 VSSD.n3291 VSSD.n3290 9.3005
R11319 VSSD.n3289 VSSD.n3237 9.3005
R11320 VSSD.n3288 VSSD.n3287 9.3005
R11321 VSSD.n3286 VSSD.n3285 9.3005
R11322 VSSD.n3283 VSSD.n3239 9.3005
R11323 VSSD.n3282 VSSD.n3281 9.3005
R11324 VSSD.n3280 VSSD.n3279 9.3005
R11325 VSSD.n3278 VSSD.n3277 9.3005
R11326 VSSD.n3276 VSSD.n3275 9.3005
R11327 VSSD.n3273 VSSD.n3243 9.3005
R11328 VSSD.n3272 VSSD.n3271 9.3005
R11329 VSSD.n3270 VSSD.n3245 9.3005
R11330 VSSD.n3269 VSSD.n3268 9.3005
R11331 VSSD.n3266 VSSD.n3246 9.3005
R11332 VSSD.n3264 VSSD.n3263 9.3005
R11333 VSSD.n3262 VSSD.n3261 9.3005
R11334 VSSD.n3259 VSSD.n3248 9.3005
R11335 VSSD.n3258 VSSD.n3257 9.3005
R11336 VSSD.n3256 VSSD.n3255 9.3005
R11337 VSSD.n2867 VSSD.n2862 9.3005
R11338 VSSD.n2869 VSSD.n2868 9.3005
R11339 VSSD.n2871 VSSD.n2860 9.3005
R11340 VSSD.n2876 VSSD.n2875 9.3005
R11341 VSSD.n2878 VSSD.n2877 9.3005
R11342 VSSD.n2884 VSSD.n2883 9.3005
R11343 VSSD.n2882 VSSD.n2881 9.3005
R11344 VSSD.n2893 VSSD.n1128 9.3005
R11345 VSSD.n2895 VSSD.n2894 9.3005
R11346 VSSD.n2898 VSSD.n1125 9.3005
R11347 VSSD.n2903 VSSD.n2902 9.3005
R11348 VSSD.n2905 VSSD.n2904 9.3005
R11349 VSSD.n2907 VSSD.n2906 9.3005
R11350 VSSD.n2909 VSSD.n2908 9.3005
R11351 VSSD.n2911 VSSD.n1121 9.3005
R11352 VSSD.n2913 VSSD.n2912 9.3005
R11353 VSSD.n2914 VSSD.n1120 9.3005
R11354 VSSD.n2916 VSSD.n2915 9.3005
R11355 VSSD.n2917 VSSD.n1118 9.3005
R11356 VSSD.n2920 VSSD.n2919 9.3005
R11357 VSSD.n2922 VSSD.n2921 9.3005
R11358 VSSD.n2923 VSSD.n1116 9.3005
R11359 VSSD.n2925 VSSD.n2924 9.3005
R11360 VSSD.n2927 VSSD.n2926 9.3005
R11361 VSSD.n2930 VSSD.n2929 9.3005
R11362 VSSD.n2932 VSSD.n2931 9.3005
R11363 VSSD.n2933 VSSD.n1108 9.3005
R11364 VSSD.n2941 VSSD.n2940 9.3005
R11365 VSSD.n2938 VSSD.n2937 9.3005
R11366 VSSD.n2951 VSSD.n2950 9.3005
R11367 VSSD.n2955 VSSD.n2954 9.3005
R11368 VSSD.n2956 VSSD.n1098 9.3005
R11369 VSSD.n2958 VSSD.n2957 9.3005
R11370 VSSD.n2961 VSSD.n1095 9.3005
R11371 VSSD.n2963 VSSD.n2962 9.3005
R11372 VSSD.n2964 VSSD.n1094 9.3005
R11373 VSSD.n2966 VSSD.n2965 9.3005
R11374 VSSD.n2967 VSSD.n1093 9.3005
R11375 VSSD.n2969 VSSD.n2968 9.3005
R11376 VSSD.n2970 VSSD.n1092 9.3005
R11377 VSSD.n2972 VSSD.n2971 9.3005
R11378 VSSD.n2973 VSSD.n1091 9.3005
R11379 VSSD.n2978 VSSD.n2977 9.3005
R11380 VSSD.n2979 VSSD.n1090 9.3005
R11381 VSSD.n2981 VSSD.n2980 9.3005
R11382 VSSD.n2982 VSSD.n1089 9.3005
R11383 VSSD.n2987 VSSD.n2986 9.3005
R11384 VSSD.n2988 VSSD.n1088 9.3005
R11385 VSSD.n2994 VSSD.n2993 9.3005
R11386 VSSD.n2997 VSSD.n2996 9.3005
R11387 VSSD.n2995 VSSD.n1082 9.3005
R11388 VSSD.n3005 VSSD.n1081 9.3005
R11389 VSSD.n3007 VSSD.n3006 9.3005
R11390 VSSD.n3010 VSSD.n3009 9.3005
R11391 VSSD.n3013 VSSD.n3012 9.3005
R11392 VSSD.n3011 VSSD.n1079 9.3005
R11393 VSSD.n3021 VSSD.n3020 9.3005
R11394 VSSD.n3054 VSSD.n3053 9.3005
R11395 VSSD.n3052 VSSD.n1078 9.3005
R11396 VSSD.n3051 VSSD.n3050 9.3005
R11397 VSSD.n3048 VSSD.n3022 9.3005
R11398 VSSD.n3047 VSSD.n3046 9.3005
R11399 VSSD.n3045 VSSD.n3044 9.3005
R11400 VSSD.n3026 VSSD.n3024 9.3005
R11401 VSSD.n3039 VSSD.n3027 9.3005
R11402 VSSD.n3038 VSSD.n3029 9.3005
R11403 VSSD.n3037 VSSD.n3030 9.3005
R11404 VSSD.n3036 VSSD.n3032 9.3005
R11405 VSSD.n3035 VSSD.n3034 9.3005
R11406 VSSD.n3033 VSSD.n1059 9.3005
R11407 VSSD.n3145 VSSD.n3144 9.3005
R11408 VSSD.n3143 VSSD.n3142 9.3005
R11409 VSSD.n1061 VSSD.n1060 9.3005
R11410 VSSD.n3137 VSSD.n3136 9.3005
R11411 VSSD.n3134 VSSD.n1065 9.3005
R11412 VSSD.n3132 VSSD.n3131 9.3005
R11413 VSSD.n3130 VSSD.n1068 9.3005
R11414 VSSD.n3129 VSSD.n3128 9.3005
R11415 VSSD.n3127 VSSD.n1069 9.3005
R11416 VSSD.n3125 VSSD.n3124 9.3005
R11417 VSSD.n3123 VSSD.n3122 9.3005
R11418 VSSD.n3121 VSSD.n1073 9.3005
R11419 VSSD.n3120 VSSD.n1074 9.3005
R11420 VSSD.n3119 VSSD.n1075 9.3005
R11421 VSSD.n3118 VSSD.n1076 9.3005
R11422 VSSD.n3116 VSSD.n3115 9.3005
R11423 VSSD.n3113 VSSD.n3112 9.3005
R11424 VSSD.n3111 VSSD.n3061 9.3005
R11425 VSSD.n3110 VSSD.n3109 9.3005
R11426 VSSD.n3108 VSSD.n3063 9.3005
R11427 VSSD.n3107 VSSD.n3106 9.3005
R11428 VSSD.n3105 VSSD.n3064 9.3005
R11429 VSSD.n3104 VSSD.n3103 9.3005
R11430 VSSD.n3102 VSSD.n3065 9.3005
R11431 VSSD.n3101 VSSD.n3100 9.3005
R11432 VSSD.n3099 VSSD.n3066 9.3005
R11433 VSSD.n3097 VSSD.n3096 9.3005
R11434 VSSD.n3095 VSSD.n3069 9.3005
R11435 VSSD.n3094 VSSD.n3093 9.3005
R11436 VSSD.n3092 VSSD.n3070 9.3005
R11437 VSSD.n3091 VSSD.n3090 9.3005
R11438 VSSD.n3089 VSSD.n3088 9.3005
R11439 VSSD.n3087 VSSD.n3074 9.3005
R11440 VSSD.n3086 VSSD.n3085 9.3005
R11441 VSSD.n3084 VSSD.n3075 9.3005
R11442 VSSD.n3083 VSSD.n3082 9.3005
R11443 VSSD.n3081 VSSD.n3076 9.3005
R11444 VSSD.n2564 VSSD.n2563 9.3005
R11445 VSSD.n2567 VSSD.n2565 9.3005
R11446 VSSD.n2569 VSSD.n2568 9.3005
R11447 VSSD.n2572 VSSD.n2551 9.3005
R11448 VSSD.n2573 VSSD.n2572 9.3005
R11449 VSSD.n2582 VSSD.n2581 9.3005
R11450 VSSD.n2584 VSSD.n2583 9.3005
R11451 VSSD.n2585 VSSD.n2545 9.3005
R11452 VSSD.n2587 VSSD.n2586 9.3005
R11453 VSSD.n2588 VSSD.n2544 9.3005
R11454 VSSD.n2590 VSSD.n2589 9.3005
R11455 VSSD.n2592 VSSD.n2591 9.3005
R11456 VSSD.n2595 VSSD.n2541 9.3005
R11457 VSSD.n2597 VSSD.n2596 9.3005
R11458 VSSD.n2598 VSSD.n2540 9.3005
R11459 VSSD.n2600 VSSD.n2599 9.3005
R11460 VSSD.n2603 VSSD.n2539 9.3005
R11461 VSSD.n2607 VSSD.n2606 9.3005
R11462 VSSD.n2608 VSSD.n2538 9.3005
R11463 VSSD.n2610 VSSD.n2609 9.3005
R11464 VSSD.n2611 VSSD.n2537 9.3005
R11465 VSSD.n2613 VSSD.n2612 9.3005
R11466 VSSD.n2614 VSSD.n2536 9.3005
R11467 VSSD.n2616 VSSD.n2615 9.3005
R11468 VSSD.n2618 VSSD.n2530 9.3005
R11469 VSSD.n2621 VSSD.n2620 9.3005
R11470 VSSD.n2531 VSSD.n1371 9.3005
R11471 VSSD.n2692 VSSD.n2630 9.3005
R11472 VSSD.n2690 VSSD.n2689 9.3005
R11473 VSSD.n2688 VSSD.n2632 9.3005
R11474 VSSD.n2687 VSSD.n2686 9.3005
R11475 VSSD.n2684 VSSD.n2683 9.3005
R11476 VSSD.n2682 VSSD.n2634 9.3005
R11477 VSSD.n2681 VSSD.n2680 9.3005
R11478 VSSD.n2676 VSSD.n2635 9.3005
R11479 VSSD.n2675 VSSD.n2673 9.3005
R11480 VSSD.n2672 VSSD.n2671 9.3005
R11481 VSSD.n2668 VSSD.n2638 9.3005
R11482 VSSD.n2666 VSSD.n2665 9.3005
R11483 VSSD.n2664 VSSD.n2663 9.3005
R11484 VSSD.n2661 VSSD.n2641 9.3005
R11485 VSSD.n2658 VSSD.n2657 9.3005
R11486 VSSD.n2656 VSSD.n2644 9.3005
R11487 VSSD.n2655 VSSD.n2654 9.3005
R11488 VSSD.n2653 VSSD.n2645 9.3005
R11489 VSSD.n2651 VSSD.n2650 9.3005
R11490 VSSD.n2649 VSSD.n1318 9.3005
R11491 VSSD.n1322 VSSD.n1319 9.3005
R11492 VSSD.n2837 VSSD.n2836 9.3005
R11493 VSSD.n2835 VSSD.n2834 9.3005
R11494 VSSD.n2833 VSSD.n2832 9.3005
R11495 VSSD.n2831 VSSD.n2830 9.3005
R11496 VSSD.n2829 VSSD.n2828 9.3005
R11497 VSSD.n2827 VSSD.n1328 9.3005
R11498 VSSD.n2824 VSSD.n2823 9.3005
R11499 VSSD.n2822 VSSD.n1329 9.3005
R11500 VSSD.n2821 VSSD.n2820 9.3005
R11501 VSSD.n2819 VSSD.n1330 9.3005
R11502 VSSD.n2818 VSSD.n1333 9.3005
R11503 VSSD.n2817 VSSD.n1334 9.3005
R11504 VSSD.n2816 VSSD.n2815 9.3005
R11505 VSSD.n2814 VSSD.n2813 9.3005
R11506 VSSD.n2812 VSSD.n1338 9.3005
R11507 VSSD.n2810 VSSD.n1342 9.3005
R11508 VSSD.n2809 VSSD.n1343 9.3005
R11509 VSSD.n2808 VSSD.n2807 9.3005
R11510 VSSD.n2806 VSSD.n1345 9.3005
R11511 VSSD.n2805 VSSD.n2804 9.3005
R11512 VSSD.n2803 VSSD.n2802 9.3005
R11513 VSSD.n1349 VSSD.n1347 9.3005
R11514 VSSD.n1363 VSSD.n1358 9.3005
R11515 VSSD.n2794 VSSD.n2793 9.3005
R11516 VSSD.n2790 VSSD.n1359 9.3005
R11517 VSSD.n2789 VSSD.n2788 9.3005
R11518 VSSD.n2787 VSSD.n2786 9.3005
R11519 VSSD.n2784 VSSD.n1365 9.3005
R11520 VSSD.n2783 VSSD.n2782 9.3005
R11521 VSSD.n2781 VSSD.n1367 9.3005
R11522 VSSD.n2780 VSSD.n2779 9.3005
R11523 VSSD.n2777 VSSD.n1368 9.3005
R11524 VSSD.n2775 VSSD.n2774 9.3005
R11525 VSSD.n2773 VSSD.n2772 9.3005
R11526 VSSD.n2771 VSSD.n1370 9.3005
R11527 VSSD.n2770 VSSD.n2769 9.3005
R11528 VSSD.n2768 VSSD.n2767 9.3005
R11529 VSSD.n2765 VSSD.n2764 9.3005
R11530 VSSD.n2763 VSSD.n2762 9.3005
R11531 VSSD.n2761 VSSD.n2699 9.3005
R11532 VSSD.n2759 VSSD.n2758 9.3005
R11533 VSSD.n2757 VSSD.n2701 9.3005
R11534 VSSD.n2756 VSSD.n2755 9.3005
R11535 VSSD.n2754 VSSD.n2702 9.3005
R11536 VSSD.n2753 VSSD.n2752 9.3005
R11537 VSSD.n2751 VSSD.n2750 9.3005
R11538 VSSD.n2748 VSSD.n2704 9.3005
R11539 VSSD.n2747 VSSD.n2746 9.3005
R11540 VSSD.n2745 VSSD.n2744 9.3005
R11541 VSSD.n2743 VSSD.n2742 9.3005
R11542 VSSD.n2741 VSSD.n2740 9.3005
R11543 VSSD.n2738 VSSD.n2708 9.3005
R11544 VSSD.n2737 VSSD.n2736 9.3005
R11545 VSSD.n2735 VSSD.n2710 9.3005
R11546 VSSD.n2734 VSSD.n2733 9.3005
R11547 VSSD.n2731 VSSD.n2711 9.3005
R11548 VSSD.n2729 VSSD.n2728 9.3005
R11549 VSSD.n2727 VSSD.n2726 9.3005
R11550 VSSD.n2724 VSSD.n2713 9.3005
R11551 VSSD.n2723 VSSD.n2722 9.3005
R11552 VSSD.n2721 VSSD.n2720 9.3005
R11553 VSSD.n2408 VSSD.n2407 9.3005
R11554 VSSD.n2409 VSSD.n2401 9.3005
R11555 VSSD.n2411 VSSD.n2410 9.3005
R11556 VSSD.n2412 VSSD.n2400 9.3005
R11557 VSSD.n2415 VSSD.n2414 9.3005
R11558 VSSD.n2417 VSSD.n2416 9.3005
R11559 VSSD.n2418 VSSD.n2398 9.3005
R11560 VSSD.n2421 VSSD.n2420 9.3005
R11561 VSSD.n2423 VSSD.n2422 9.3005
R11562 VSSD.n2424 VSSD.n2396 9.3005
R11563 VSSD.n2426 VSSD.n2425 9.3005
R11564 VSSD.n2428 VSSD.n2427 9.3005
R11565 VSSD.n1487 VSSD.n1480 9.3005
R11566 VSSD.n1489 VSSD.n1488 9.3005
R11567 VSSD.n1493 VSSD.n1492 9.3005
R11568 VSSD.n1494 VSSD.n1479 9.3005
R11569 VSSD.n1496 VSSD.n1495 9.3005
R11570 VSSD.n1563 VSSD.n1562 9.3005
R11571 VSSD.n1560 VSSD.n1559 9.3005
R11572 VSSD.n1551 VSSD.n1498 9.3005
R11573 VSSD.n1550 VSSD.n1549 9.3005
R11574 VSSD.n1548 VSSD.n1499 9.3005
R11575 VSSD.n1547 VSSD.n1546 9.3005
R11576 VSSD.n1545 VSSD.n1544 9.3005
R11577 VSSD.n1543 VSSD.n1504 9.3005
R11578 VSSD.n1541 VSSD.n1540 9.3005
R11579 VSSD.n1539 VSSD.n1506 9.3005
R11580 VSSD.n1538 VSSD.n1537 9.3005
R11581 VSSD.n1536 VSSD.n1507 9.3005
R11582 VSSD.n1535 VSSD.n1508 9.3005
R11583 VSSD.n1534 VSSD.n1533 9.3005
R11584 VSSD.n1532 VSSD.n1531 9.3005
R11585 VSSD.n1529 VSSD.n1510 9.3005
R11586 VSSD.n1527 VSSD.n1526 9.3005
R11587 VSSD.n1525 VSSD.n1524 9.3005
R11588 VSSD.n1523 VSSD.n1522 9.3005
R11589 VSSD.n1521 VSSD.n1520 9.3005
R11590 VSSD.n1519 VSSD.n1517 9.3005
R11591 VSSD.n1518 VSSD.n1379 9.3005
R11592 VSSD.n2521 VSSD.n2520 9.3005
R11593 VSSD.n2518 VSSD.n2517 9.3005
R11594 VSSD.n2510 VSSD.n1382 9.3005
R11595 VSSD.n2509 VSSD.n2508 9.3005
R11596 VSSD.n2507 VSSD.n2506 9.3005
R11597 VSSD.n2505 VSSD.n1385 9.3005
R11598 VSSD.n2504 VSSD.n2503 9.3005
R11599 VSSD.n2502 VSSD.n1386 9.3005
R11600 VSSD.n2499 VSSD.n2498 9.3005
R11601 VSSD.n2497 VSSD.n1389 9.3005
R11602 VSSD.n2496 VSSD.n2495 9.3005
R11603 VSSD.n2494 VSSD.n2493 9.3005
R11604 VSSD.n2492 VSSD.n2491 9.3005
R11605 VSSD.n2489 VSSD.n1392 9.3005
R11606 VSSD.n2488 VSSD.n2487 9.3005
R11607 VSSD.n2486 VSSD.n1394 9.3005
R11608 VSSD.n2485 VSSD.n2484 9.3005
R11609 VSSD.n2483 VSSD.n1395 9.3005
R11610 VSSD.n2482 VSSD.n2481 9.3005
R11611 VSSD.n2480 VSSD.n1396 9.3005
R11612 VSSD.n2479 VSSD.n2478 9.3005
R11613 VSSD.n2476 VSSD.n2475 9.3005
R11614 VSSD.n1408 VSSD.n1407 9.3005
R11615 VSSD.n1411 VSSD.n1410 9.3005
R11616 VSSD.n2465 VSSD.n2464 9.3005
R11617 VSSD.n2462 VSSD.n1406 9.3005
R11618 VSSD.n2460 VSSD.n2459 9.3005
R11619 VSSD.n2457 VSSD.n2456 9.3005
R11620 VSSD.n2318 VSSD.n1416 9.3005
R11621 VSSD.n2321 VSSD.n2319 9.3005
R11622 VSSD.n2323 VSSD.n2322 9.3005
R11623 VSSD.n2325 VSSD.n2324 9.3005
R11624 VSSD.n2327 VSSD.n2316 9.3005
R11625 VSSD.n2331 VSSD.n2330 9.3005
R11626 VSSD.n2332 VSSD.n2314 9.3005
R11627 VSSD.n2334 VSSD.n2333 9.3005
R11628 VSSD.n2335 VSSD.n2313 9.3005
R11629 VSSD.n2340 VSSD.n2339 9.3005
R11630 VSSD.n2341 VSSD.n2312 9.3005
R11631 VSSD.n2343 VSSD.n2342 9.3005
R11632 VSSD.n2345 VSSD.n2344 9.3005
R11633 VSSD.n2308 VSSD.n1425 9.3005
R11634 VSSD.n2355 VSSD.n2354 9.3005
R11635 VSSD.n2358 VSSD.n1424 9.3005
R11636 VSSD.n2362 VSSD.n2361 9.3005
R11637 VSSD.n2363 VSSD.n1423 9.3005
R11638 VSSD.n2365 VSSD.n2364 9.3005
R11639 VSSD.n2366 VSSD.n1422 9.3005
R11640 VSSD.n2369 VSSD.n2368 9.3005
R11641 VSSD.n2371 VSSD.n2370 9.3005
R11642 VSSD.n2373 VSSD.n2372 9.3005
R11643 VSSD.n2375 VSSD.n2374 9.3005
R11644 VSSD.n2376 VSSD.n1418 9.3005
R11645 VSSD.n2381 VSSD.n2380 9.3005
R11646 VSSD.n2382 VSSD.n1417 9.3005
R11647 VSSD.n2453 VSSD.n2383 9.3005
R11648 VSSD.n2452 VSSD.n2451 9.3005
R11649 VSSD.n2450 VSSD.n2385 9.3005
R11650 VSSD.n2449 VSSD.n2448 9.3005
R11651 VSSD.n2447 VSSD.n2386 9.3005
R11652 VSSD.n2446 VSSD.n2445 9.3005
R11653 VSSD.n2444 VSSD.n2389 9.3005
R11654 VSSD.n2443 VSSD.n2442 9.3005
R11655 VSSD.n2441 VSSD.n2390 9.3005
R11656 VSSD.n2439 VSSD.n2438 9.3005
R11657 VSSD.n2437 VSSD.n2436 9.3005
R11658 VSSD.n2435 VSSD.n2393 9.3005
R11659 VSSD.n2434 VSSD.n2433 9.3005
R11660 VSSD.n2432 VSSD.n2431 9.3005
R11661 VSSD.n1969 VSSD.n1968 9.3005
R11662 VSSD.n1972 VSSD.n1971 9.3005
R11663 VSSD.n1974 VSSD.n1973 9.3005
R11664 VSSD.n1977 VSSD.n1976 9.3005
R11665 VSSD.n1979 VSSD.n1978 9.3005
R11666 VSSD.n1981 VSSD.n1980 9.3005
R11667 VSSD.n1961 VSSD.n1960 9.3005
R11668 VSSD.n1991 VSSD.n1990 9.3005
R11669 VSSD.n1992 VSSD.n1467 9.3005
R11670 VSSD.n1995 VSSD.n1994 9.3005
R11671 VSSD.n1996 VSSD.n1466 9.3005
R11672 VSSD.n1998 VSSD.n1997 9.3005
R11673 VSSD.n2000 VSSD.n1464 9.3005
R11674 VSSD.n2004 VSSD.n2003 9.3005
R11675 VSSD.n2005 VSSD.n1463 9.3005
R11676 VSSD.n2007 VSSD.n2006 9.3005
R11677 VSSD.n2008 VSSD.n1462 9.3005
R11678 VSSD.n2010 VSSD.n2009 9.3005
R11679 VSSD.n2011 VSSD.n1461 9.3005
R11680 VSSD.n2013 VSSD.n2012 9.3005
R11681 VSSD.n2015 VSSD.n1459 9.3005
R11682 VSSD.n2018 VSSD.n2017 9.3005
R11683 VSSD.n2019 VSSD.n1458 9.3005
R11684 VSSD.n2021 VSSD.n2020 9.3005
R11685 VSSD.n2023 VSSD.n1456 9.3005
R11686 VSSD.n2028 VSSD.n2027 9.3005
R11687 VSSD.n2031 VSSD.n1451 9.3005
R11688 VSSD.n2037 VSSD.n1451 9.3005
R11689 VSSD.n2032 VSSD.n1451 9.3005
R11690 VSSD.n2105 VSSD.n2046 9.3005
R11691 VSSD.n2103 VSSD.n2102 9.3005
R11692 VSSD.n2101 VSSD.n2100 9.3005
R11693 VSSD.n2097 VSSD.n2049 9.3005
R11694 VSSD.n2096 VSSD.n2095 9.3005
R11695 VSSD.n2094 VSSD.n2093 9.3005
R11696 VSSD.n2092 VSSD.n2053 9.3005
R11697 VSSD.n2089 VSSD.n2088 9.3005
R11698 VSSD.n2087 VSSD.n2056 9.3005
R11699 VSSD.n2086 VSSD.n2085 9.3005
R11700 VSSD.n2084 VSSD.n2057 9.3005
R11701 VSSD.n2083 VSSD.n2082 9.3005
R11702 VSSD.n2081 VSSD.n2080 9.3005
R11703 VSSD.n2079 VSSD.n2063 9.3005
R11704 VSSD.n2078 VSSD.n2065 9.3005
R11705 VSSD.n2077 VSSD.n2076 9.3005
R11706 VSSD.n2075 VSSD.n2066 9.3005
R11707 VSSD.n2074 VSSD.n2073 9.3005
R11708 VSSD.n2071 VSSD.n2067 9.3005
R11709 VSSD.n2070 VSSD.n1436 9.3005
R11710 VSSD.n2069 VSSD.n1437 9.3005
R11711 VSSD.n2289 VSSD.n2288 9.3005
R11712 VSSD.n2286 VSSD.n2285 9.3005
R11713 VSSD.n2284 VSSD.n2283 9.3005
R11714 VSSD.n2281 VSSD.n1447 9.3005
R11715 VSSD.n2280 VSSD.n2279 9.3005
R11716 VSSD.n2278 VSSD.n2277 9.3005
R11717 VSSD.n2276 VSSD.n2275 9.3005
R11718 VSSD.n2274 VSSD.n2273 9.3005
R11719 VSSD.n2272 VSSD.n2110 9.3005
R11720 VSSD.n2271 VSSD.n2270 9.3005
R11721 VSSD.n2269 VSSD.n2111 9.3005
R11722 VSSD.n2268 VSSD.n2267 9.3005
R11723 VSSD.n2115 VSSD.n2112 9.3005
R11724 VSSD.n2262 VSSD.n2261 9.3005
R11725 VSSD.n2260 VSSD.n2118 9.3005
R11726 VSSD.n2259 VSSD.n2258 9.3005
R11727 VSSD.n2256 VSSD.n2119 9.3005
R11728 VSSD.n2255 VSSD.n2123 9.3005
R11729 VSSD.n2254 VSSD.n2253 9.3005
R11730 VSSD.n2126 VSSD.n2124 9.3005
R11731 VSSD.n2238 VSSD.n2237 9.3005
R11732 VSSD.n2236 VSSD.n2128 9.3005
R11733 VSSD.n2235 VSSD.n2234 9.3005
R11734 VSSD.n2233 VSSD.n2129 9.3005
R11735 VSSD.n2232 VSSD.n2231 9.3005
R11736 VSSD.n2229 VSSD.n2130 9.3005
R11737 VSSD.n2228 VSSD.n2227 9.3005
R11738 VSSD.n2226 VSSD.n2133 9.3005
R11739 VSSD.n2225 VSSD.n2224 9.3005
R11740 VSSD.n2138 VSSD.n2134 9.3005
R11741 VSSD.n2219 VSSD.n2218 9.3005
R11742 VSSD.n2217 VSSD.n2216 9.3005
R11743 VSSD.n2215 VSSD.n2214 9.3005
R11744 VSSD.n2213 VSSD.n2212 9.3005
R11745 VSSD.n2211 VSSD.n2143 9.3005
R11746 VSSD.n2210 VSSD.n2209 9.3005
R11747 VSSD.n2208 VSSD.n2207 9.3005
R11748 VSSD.n2205 VSSD.n2146 9.3005
R11749 VSSD.n2204 VSSD.n2147 9.3005
R11750 VSSD.n2203 VSSD.n2202 9.3005
R11751 VSSD.n2201 VSSD.n2148 9.3005
R11752 VSSD.n2200 VSSD.n2199 9.3005
R11753 VSSD.n2198 VSSD.n2149 9.3005
R11754 VSSD.n2196 VSSD.n2195 9.3005
R11755 VSSD.n2194 VSSD.n2151 9.3005
R11756 VSSD.n2193 VSSD.n2192 9.3005
R11757 VSSD.n2191 VSSD.n2152 9.3005
R11758 VSSD.n2190 VSSD.n2189 9.3005
R11759 VSSD.n2188 VSSD.n2187 9.3005
R11760 VSSD.n2186 VSSD.n2157 9.3005
R11761 VSSD.n2184 VSSD.n2183 9.3005
R11762 VSSD.n2182 VSSD.n2159 9.3005
R11763 VSSD.n2181 VSSD.n2180 9.3005
R11764 VSSD.n2178 VSSD.n2160 9.3005
R11765 VSSD.n2176 VSSD.n2175 9.3005
R11766 VSSD.n2174 VSSD.n2173 9.3005
R11767 VSSD.n2172 VSSD.n2171 9.3005
R11768 VSSD.n2170 VSSD.n2169 9.3005
R11769 VSSD.n1889 VSSD.n1888 9.3005
R11770 VSSD.n1858 VSSD.n1638 9.3005
R11771 VSSD.n1649 VSSD.n1648 9.3005
R11772 VSSD.n1651 VSSD.n1644 9.3005
R11773 VSSD.n1844 VSSD.n1843 9.3005
R11774 VSSD.n1841 VSSD.n1645 9.3005
R11775 VSSD.n1840 VSSD.n1839 9.3005
R11776 VSSD.n1838 VSSD.n1654 9.3005
R11777 VSSD.n1837 VSSD.n1836 9.3005
R11778 VSSD.n1832 VSSD.n1831 9.3005
R11779 VSSD.n1830 VSSD.n1829 9.3005
R11780 VSSD.n1826 VSSD.n1658 9.3005
R11781 VSSD.n1663 VSSD.n1659 9.3005
R11782 VSSD.n1784 VSSD.n1687 9.3005
R11783 VSSD.n1778 VSSD.n1777 9.3005
R11784 VSSD.n1775 VSSD.n1691 9.3005
R11785 VSSD.n1773 VSSD.n1772 9.3005
R11786 VSSD.n1771 VSSD.n1770 9.3005
R11787 VSSD.n1769 VSSD.n1768 9.3005
R11788 VSSD.n1767 VSSD.n1766 9.3005
R11789 VSSD.n1698 VSSD.n1695 9.3005
R11790 VSSD.n1761 VSSD.n1760 9.3005
R11791 VSSD.n1759 VSSD.n1697 9.3005
R11792 VSSD.n1758 VSSD.n1757 9.3005
R11793 VSSD.n1756 VSSD.n1699 9.3005
R11794 VSSD.n1755 VSSD.n1754 9.3005
R11795 VSSD.n1753 VSSD.n1701 9.3005
R11796 VSSD.n1752 VSSD.n1751 9.3005
R11797 VSSD.n1749 VSSD.n1702 9.3005
R11798 VSSD.n1747 VSSD.n1746 9.3005
R11799 VSSD.n1745 VSSD.n1704 9.3005
R11800 VSSD.n1744 VSSD.n1743 9.3005
R11801 VSSD.n1742 VSSD.n1741 9.3005
R11802 VSSD.n1740 VSSD.n1739 9.3005
R11803 VSSD.n1737 VSSD.n1707 9.3005
R11804 VSSD.n1736 VSSD.n1735 9.3005
R11805 VSSD.n1734 VSSD.n1709 9.3005
R11806 VSSD.n1733 VSSD.n1732 9.3005
R11807 VSSD.n1730 VSSD.n1710 9.3005
R11808 VSSD.n1728 VSSD.n1727 9.3005
R11809 VSSD.n1726 VSSD.n1725 9.3005
R11810 VSSD.n1723 VSSD.n1712 9.3005
R11811 VSSD.n1722 VSSD.n1721 9.3005
R11812 VSSD.n1720 VSSD.n1719 9.3005
R11813 VSSD.n1779 VSSD.n1690 9.3005
R11814 VSSD.n1781 VSSD.n1780 9.3005
R11815 VSSD.n1786 VSSD.n1785 9.3005
R11816 VSSD.n1787 VSSD.n1686 9.3005
R11817 VSSD.n1789 VSSD.n1788 9.3005
R11818 VSSD.n1790 VSSD.n1684 9.3005
R11819 VSSD.n1794 VSSD.n1793 9.3005
R11820 VSSD.n1685 VSSD.n1683 9.3005
R11821 VSSD.n1674 VSSD.n1672 9.3005
R11822 VSSD.n1803 VSSD.n1802 9.3005
R11823 VSSD.n1807 VSSD.n1806 9.3005
R11824 VSSD.n1808 VSSD.n1670 9.3005
R11825 VSSD.n1810 VSSD.n1809 9.3005
R11826 VSSD.n1811 VSSD.n1667 9.3005
R11827 VSSD.n1813 VSSD.n1812 9.3005
R11828 VSSD.n1815 VSSD.n1814 9.3005
R11829 VSSD.n1817 VSSD.n1816 9.3005
R11830 VSSD.n1819 VSSD.n1818 9.3005
R11831 VSSD.n1825 VSSD.n1824 9.3005
R11832 VSSD.n1828 VSSD.n1827 9.3005
R11833 VSSD.n1855 VSSD.n1854 9.3005
R11834 VSSD.n1857 VSSD.n1856 9.3005
R11835 VSSD.n1860 VSSD.n1859 9.3005
R11836 VSSD.n1861 VSSD.n1636 9.3005
R11837 VSSD.n1863 VSSD.n1862 9.3005
R11838 VSSD.n1865 VSSD.n1864 9.3005
R11839 VSSD.n1866 VSSD.n1633 9.3005
R11840 VSSD.n1868 VSSD.n1867 9.3005
R11841 VSSD.n1869 VSSD.n1632 9.3005
R11842 VSSD.n1871 VSSD.n1870 9.3005
R11843 VSSD.n1874 VSSD.n1629 9.3005
R11844 VSSD.n1876 VSSD.n1875 9.3005
R11845 VSSD.n1877 VSSD.n1628 9.3005
R11846 VSSD.n1879 VSSD.n1878 9.3005
R11847 VSSD.n1880 VSSD.n1627 9.3005
R11848 VSSD.n1884 VSSD.n1883 9.3005
R11849 VSSD.n1885 VSSD.n1626 9.3005
R11850 VSSD.n1887 VSSD.n1886 9.3005
R11851 VSSD.n1624 VSSD.n1623 9.3005
R11852 VSSD.n1620 VSSD.n1592 9.3005
R11853 VSSD.n1900 VSSD.n1899 9.3005
R11854 VSSD.n1903 VSSD.n1591 9.3005
R11855 VSSD.n1906 VSSD.n1905 9.3005
R11856 VSSD.n1908 VSSD.n1907 9.3005
R11857 VSSD.n1910 VSSD.n1909 9.3005
R11858 VSSD.n1911 VSSD.n1587 9.3005
R11859 VSSD.n1913 VSSD.n1912 9.3005
R11860 VSSD.n1914 VSSD.n1586 9.3005
R11861 VSSD.n1917 VSSD.n1916 9.3005
R11862 VSSD.n1919 VSSD.n1918 9.3005
R11863 VSSD.n1604 VSSD.n1598 9.3005
R11864 VSSD.n1615 VSSD.n1614 9.3005
R11865 VSSD.n1613 VSSD.n1612 9.3005
R11866 VSSD.n1610 VSSD.n1606 9.3005
R11867 VSSD.n1605 VSSD.n1575 9.3005
R11868 VSSD.n1948 VSSD.n1947 9.3005
R11869 VSSD.n1945 VSSD.n1944 9.3005
R11870 VSSD.n1936 VSSD.n1576 9.3005
R11871 VSSD.n1935 VSSD.n1934 9.3005
R11872 VSSD.n1933 VSSD.n1577 9.3005
R11873 VSSD.n1932 VSSD.n1931 9.3005
R11874 VSSD.n1930 VSSD.n1580 9.3005
R11875 VSSD.n1929 VSSD.n1928 9.3005
R11876 VSSD.n1925 VSSD.n1581 9.3005
R11877 VSSD.n1924 VSSD.n1923 9.3005
R11878 VSSD.n1922 VSSD.n1583 9.3005
R11879 VSSD.n1921 VSSD.n1920 9.3005
R11880 VSSD.n3612 VSSD.n3611 9.3005
R11881 VSSD.n3614 VSSD.n3613 9.3005
R11882 VSSD.n3616 VSSD.n3615 9.3005
R11883 VSSD.n3618 VSSD.n3617 9.3005
R11884 VSSD.n3619 VSSD.n3605 9.3005
R11885 VSSD.n3621 VSSD.n3620 9.3005
R11886 VSSD.n3623 VSSD.n3622 9.3005
R11887 VSSD.n3624 VSSD.n3603 9.3005
R11888 VSSD.n3626 VSSD.n3625 9.3005
R11889 VSSD.n3627 VSSD.n3602 9.3005
R11890 VSSD.n3629 VSSD.n3628 9.3005
R11891 VSSD.n3630 VSSD.n3601 9.3005
R11892 VSSD.n3632 VSSD.n3631 9.3005
R11893 VSSD.n3634 VSSD.n3633 9.3005
R11894 VSSD.n3402 VSSD.n3399 9.3005
R11895 VSSD.n3405 VSSD.n3404 9.3005
R11896 VSSD.n3406 VSSD.n132 9.3005
R11897 VSSD.n3408 VSSD.n3407 9.3005
R11898 VSSD.n3409 VSSD.n131 9.3005
R11899 VSSD.n3413 VSSD.n3412 9.3005
R11900 VSSD.n3415 VSSD.n3414 9.3005
R11901 VSSD.n3417 VSSD.n3416 9.3005
R11902 VSSD.n3428 VSSD.n3427 9.3005
R11903 VSSD.n3429 VSSD.n119 9.3005
R11904 VSSD.n3431 VSSD.n3430 9.3005
R11905 VSSD.n3432 VSSD.n118 9.3005
R11906 VSSD.n3434 VSSD.n3433 9.3005
R11907 VSSD.n3435 VSSD.n117 9.3005
R11908 VSSD.n3437 VSSD.n3436 9.3005
R11909 VSSD.n3439 VSSD.n3438 9.3005
R11910 VSSD.n3440 VSSD.n115 9.3005
R11911 VSSD.n3442 VSSD.n3441 9.3005
R11912 VSSD.n3444 VSSD.n3443 9.3005
R11913 VSSD.n3446 VSSD.n3445 9.3005
R11914 VSSD.n3448 VSSD.n3447 9.3005
R11915 VSSD.n3449 VSSD.n112 9.3005
R11916 VSSD.n3451 VSSD.n3450 9.3005
R11917 VSSD.n3452 VSSD.n111 9.3005
R11918 VSSD.n3454 VSSD.n3453 9.3005
R11919 VSSD.n3455 VSSD.n110 9.3005
R11920 VSSD.n3457 VSSD.n3456 9.3005
R11921 VSSD.n3459 VSSD.n3458 9.3005
R11922 VSSD.n3460 VSSD.n103 9.3005
R11923 VSSD.n3463 VSSD.n3462 9.3005
R11924 VSSD.n104 VSSD.n95 9.3005
R11925 VSSD.n3473 VSSD.n3472 9.3005
R11926 VSSD.n3474 VSSD.n94 9.3005
R11927 VSSD.n3478 VSSD.n3477 9.3005
R11928 VSSD.n3480 VSSD.n3479 9.3005
R11929 VSSD.n3482 VSSD.n3481 9.3005
R11930 VSSD.n3484 VSSD.n3483 9.3005
R11931 VSSD.n3485 VSSD.n91 9.3005
R11932 VSSD.n3487 VSSD.n3486 9.3005
R11933 VSSD.n3488 VSSD.n90 9.3005
R11934 VSSD.n3490 VSSD.n3489 9.3005
R11935 VSSD.n3491 VSSD.n89 9.3005
R11936 VSSD.n3493 VSSD.n3492 9.3005
R11937 VSSD.n3495 VSSD.n3494 9.3005
R11938 VSSD.n3496 VSSD.n87 9.3005
R11939 VSSD.n3498 VSSD.n3497 9.3005
R11940 VSSD.n3500 VSSD.n3499 9.3005
R11941 VSSD.n3503 VSSD.n3502 9.3005
R11942 VSSD.n3504 VSSD.n85 9.3005
R11943 VSSD.n3506 VSSD.n3505 9.3005
R11944 VSSD.n3508 VSSD.n3507 9.3005
R11945 VSSD.n3509 VSSD.n77 9.3005
R11946 VSSD.n3522 VSSD.n3521 9.3005
R11947 VSSD.n3523 VSSD.n76 9.3005
R11948 VSSD.n3525 VSSD.n3524 9.3005
R11949 VSSD.n3527 VSSD.n3526 9.3005
R11950 VSSD.n3528 VSSD.n74 9.3005
R11951 VSSD.n3531 VSSD.n3530 9.3005
R11952 VSSD.n3532 VSSD.n72 9.3005
R11953 VSSD.n3534 VSSD.n3533 9.3005
R11954 VSSD.n3535 VSSD.n71 9.3005
R11955 VSSD.n3539 VSSD.n3538 9.3005
R11956 VSSD.n3541 VSSD.n3540 9.3005
R11957 VSSD.n3543 VSSD.n3542 9.3005
R11958 VSSD.n3545 VSSD.n3544 9.3005
R11959 VSSD.n3546 VSSD.n68 9.3005
R11960 VSSD.n3548 VSSD.n3547 9.3005
R11961 VSSD.n3549 VSSD.n67 9.3005
R11962 VSSD.n3551 VSSD.n3550 9.3005
R11963 VSSD.n3552 VSSD.n66 9.3005
R11964 VSSD.n3554 VSSD.n3553 9.3005
R11965 VSSD.n3556 VSSD.n3555 9.3005
R11966 VSSD.n3560 VSSD.n3559 9.3005
R11967 VSSD.n3558 VSSD.n3557 9.3005
R11968 VSSD.n3570 VSSD.n3569 9.3005
R11969 VSSD.n3572 VSSD.n3571 9.3005
R11970 VSSD.n3574 VSSD.n3573 9.3005
R11971 VSSD.n3575 VSSD.n52 9.3005
R11972 VSSD.n3577 VSSD.n3576 9.3005
R11973 VSSD.n3578 VSSD.n51 9.3005
R11974 VSSD.n3580 VSSD.n3579 9.3005
R11975 VSSD.n3581 VSSD.n50 9.3005
R11976 VSSD.n3583 VSSD.n3582 9.3005
R11977 VSSD.n3585 VSSD.n3584 9.3005
R11978 VSSD.n3586 VSSD.n48 9.3005
R11979 VSSD.n3589 VSSD.n3588 9.3005
R11980 VSSD.n3590 VSSD.n47 9.3005
R11981 VSSD.n3656 VSSD.n3591 9.3005
R11982 VSSD.n3655 VSSD.n3654 9.3005
R11983 VSSD.n3653 VSSD.n3592 9.3005
R11984 VSSD.n3652 VSSD.n3651 9.3005
R11985 VSSD.n3650 VSSD.n3593 9.3005
R11986 VSSD.n3649 VSSD.n3648 9.3005
R11987 VSSD.n3647 VSSD.n3595 9.3005
R11988 VSSD.n3646 VSSD.n3645 9.3005
R11989 VSSD.n3644 VSSD.n3596 9.3005
R11990 VSSD.n3643 VSSD.n3642 9.3005
R11991 VSSD.n3641 VSSD.n3640 9.3005
R11992 VSSD.n3639 VSSD.n3598 9.3005
R11993 VSSD.n3638 VSSD.n3637 9.3005
R11994 VSSD.n3636 VSSD.n3635 9.3005
R11995 VSSD.n272 VSSD.n271 9.3005
R11996 VSSD.n274 VSSD.n273 9.3005
R11997 VSSD.n275 VSSD.n265 9.3005
R11998 VSSD.n277 VSSD.n276 9.3005
R11999 VSSD.n279 VSSD.n278 9.3005
R12000 VSSD.n280 VSSD.n263 9.3005
R12001 VSSD.n282 VSSD.n281 9.3005
R12002 VSSD.n283 VSSD.n262 9.3005
R12003 VSSD.n285 VSSD.n284 9.3005
R12004 VSSD.n286 VSSD.n261 9.3005
R12005 VSSD.n288 VSSD.n287 9.3005
R12006 VSSD.n290 VSSD.n289 9.3005
R12007 VSSD.n487 VSSD.n486 9.3005
R12008 VSSD.n485 VSSD.n140 9.3005
R12009 VSSD.n484 VSSD.n483 9.3005
R12010 VSSD.n482 VSSD.n481 9.3005
R12011 VSSD.n144 VSSD.n142 9.3005
R12012 VSSD.n473 VSSD.n472 9.3005
R12013 VSSD.n469 VSSD.n153 9.3005
R12014 VSSD.n468 VSSD.n467 9.3005
R12015 VSSD.n466 VSSD.n156 9.3005
R12016 VSSD.n465 VSSD.n464 9.3005
R12017 VSSD.n461 VSSD.n157 9.3005
R12018 VSSD.n458 VSSD.n457 9.3005
R12019 VSSD.n456 VSSD.n158 9.3005
R12020 VSSD.n455 VSSD.n454 9.3005
R12021 VSSD.n453 VSSD.n159 9.3005
R12022 VSSD.n452 VSSD.n451 9.3005
R12023 VSSD.n450 VSSD.n160 9.3005
R12024 VSSD.n449 VSSD.n448 9.3005
R12025 VSSD.n447 VSSD.n161 9.3005
R12026 VSSD.n445 VSSD.n443 9.3005
R12027 VSSD.n442 VSSD.n162 9.3005
R12028 VSSD.n441 VSSD.n440 9.3005
R12029 VSSD.n438 VSSD.n437 9.3005
R12030 VSSD.n436 VSSD.n435 9.3005
R12031 VSSD.n434 VSSD.n433 9.3005
R12032 VSSD.n166 VSSD.n165 9.3005
R12033 VSSD.n176 VSSD.n175 9.3005
R12034 VSSD.n423 VSSD.n422 9.3005
R12035 VSSD.n182 VSSD.n178 9.3005
R12036 VSSD.n417 VSSD.n416 9.3005
R12037 VSSD.n415 VSSD.n181 9.3005
R12038 VSSD.n414 VSSD.n413 9.3005
R12039 VSSD.n412 VSSD.n183 9.3005
R12040 VSSD.n411 VSSD.n410 9.3005
R12041 VSSD.n409 VSSD.n408 9.3005
R12042 VSSD.n407 VSSD.n186 9.3005
R12043 VSSD.n406 VSSD.n405 9.3005
R12044 VSSD.n404 VSSD.n189 9.3005
R12045 VSSD.n403 VSSD.n402 9.3005
R12046 VSSD.n400 VSSD.n190 9.3005
R12047 VSSD.n398 VSSD.n397 9.3005
R12048 VSSD.n396 VSSD.n193 9.3005
R12049 VSSD.n395 VSSD.n394 9.3005
R12050 VSSD.n393 VSSD.n194 9.3005
R12051 VSSD.n392 VSSD.n391 9.3005
R12052 VSSD.n390 VSSD.n389 9.3005
R12053 VSSD.n388 VSSD.n387 9.3005
R12054 VSSD.n206 VSSD.n200 9.3005
R12055 VSSD.n209 VSSD.n208 9.3005
R12056 VSSD.n377 VSSD.n376 9.3005
R12057 VSSD.n375 VSSD.n211 9.3005
R12058 VSSD.n374 VSSD.n373 9.3005
R12059 VSSD.n372 VSSD.n371 9.3005
R12060 VSSD.n369 VSSD.n213 9.3005
R12061 VSSD.n366 VSSD.n365 9.3005
R12062 VSSD.n364 VSSD.n214 9.3005
R12063 VSSD.n363 VSSD.n362 9.3005
R12064 VSSD.n361 VSSD.n215 9.3005
R12065 VSSD.n360 VSSD.n359 9.3005
R12066 VSSD.n358 VSSD.n357 9.3005
R12067 VSSD.n355 VSSD.n219 9.3005
R12068 VSSD.n354 VSSD.n353 9.3005
R12069 VSSD.n352 VSSD.n220 9.3005
R12070 VSSD.n351 VSSD.n350 9.3005
R12071 VSSD.n348 VSSD.n221 9.3005
R12072 VSSD.n347 VSSD.n346 9.3005
R12073 VSSD.n345 VSSD.n344 9.3005
R12074 VSSD.n343 VSSD.n225 9.3005
R12075 VSSD.n342 VSSD.n341 9.3005
R12076 VSSD.n228 VSSD.n226 9.3005
R12077 VSSD.n239 VSSD.n237 9.3005
R12078 VSSD.n333 VSSD.n332 9.3005
R12079 VSSD.n330 VSSD.n238 9.3005
R12080 VSSD.n329 VSSD.n328 9.3005
R12081 VSSD.n327 VSSD.n242 9.3005
R12082 VSSD.n326 VSSD.n325 9.3005
R12083 VSSD.n323 VSSD.n243 9.3005
R12084 VSSD.n322 VSSD.n321 9.3005
R12085 VSSD.n320 VSSD.n319 9.3005
R12086 VSSD.n317 VSSD.n246 9.3005
R12087 VSSD.n316 VSSD.n315 9.3005
R12088 VSSD.n312 VSSD.n311 9.3005
R12089 VSSD.n311 VSSD.n250 9.3005
R12090 VSSD.n310 VSSD.n309 9.3005
R12091 VSSD.n308 VSSD.n307 9.3005
R12092 VSSD.n306 VSSD.n254 9.3005
R12093 VSSD.n305 VSSD.n304 9.3005
R12094 VSSD.n303 VSSD.n255 9.3005
R12095 VSSD.n302 VSSD.n301 9.3005
R12096 VSSD.n300 VSSD.n256 9.3005
R12097 VSSD.n299 VSSD.n298 9.3005
R12098 VSSD.n297 VSSD.n296 9.3005
R12099 VSSD.n295 VSSD.n258 9.3005
R12100 VSSD.n294 VSSD.n293 9.3005
R12101 VSSD.n292 VSSD.n291 9.3005
R12102 VSSD.n138 VSSD.n133 9.3005
R12103 VSSD.n489 VSSD.n139 9.3005
R12104 VSSD.n3787 VSSD.n3786 9.3005
R12105 VSSD.n3785 VSSD.n3784 9.3005
R12106 VSSD.n3782 VSSD.n1 9.3005
R12107 VSSD.n3781 VSSD.n3780 9.3005
R12108 VSSD.n3779 VSSD.n3778 9.3005
R12109 VSSD.n3777 VSSD.n3 9.3005
R12110 VSSD.n3776 VSSD.n3775 9.3005
R12111 VSSD.n3774 VSSD.n3773 9.3005
R12112 VSSD.n3772 VSSD.n3771 9.3005
R12113 VSSD.n3770 VSSD.n3769 9.3005
R12114 VSSD.n3766 VSSD.n6 9.3005
R12115 VSSD.n3764 VSSD.n3763 9.3005
R12116 VSSD.n565 VSSD.n560 9.3005
R12117 VSSD.n670 VSSD.n669 9.3005
R12118 VSSD.n668 VSSD.n559 9.3005
R12119 VSSD.n664 VSSD.n663 9.3005
R12120 VSSD.n582 VSSD.n571 9.3005
R12121 VSSD.n655 VSSD.n654 9.3005
R12122 VSSD.n583 VSSD.n581 9.3005
R12123 VSSD.n649 VSSD.n648 9.3005
R12124 VSSD.n647 VSSD.n646 9.3005
R12125 VSSD.n645 VSSD.n644 9.3005
R12126 VSSD.n643 VSSD.n642 9.3005
R12127 VSSD.n640 VSSD.n587 9.3005
R12128 VSSD.n639 VSSD.n638 9.3005
R12129 VSSD.n637 VSSD.n588 9.3005
R12130 VSSD.n636 VSSD.n635 9.3005
R12131 VSSD.n634 VSSD.n633 9.3005
R12132 VSSD.n632 VSSD.n631 9.3005
R12133 VSSD.n629 VSSD.n591 9.3005
R12134 VSSD.n628 VSSD.n627 9.3005
R12135 VSSD.n626 VSSD.n592 9.3005
R12136 VSSD.n625 VSSD.n624 9.3005
R12137 VSSD.n623 VSSD.n622 9.3005
R12138 VSSD.n621 VSSD.n620 9.3005
R12139 VSSD.n618 VSSD.n595 9.3005
R12140 VSSD.n617 VSSD.n616 9.3005
R12141 VSSD.n599 VSSD.n597 9.3005
R12142 VSSD.n606 VSSD.n556 9.3005
R12143 VSSD.n673 VSSD.n558 9.3005
R12144 VSSD.n678 VSSD.n552 9.3005
R12145 VSSD.n682 VSSD.n681 9.3005
R12146 VSSD.n683 VSSD.n551 9.3005
R12147 VSSD.n685 VSSD.n684 9.3005
R12148 VSSD.n686 VSSD.n550 9.3005
R12149 VSSD.n689 VSSD.n688 9.3005
R12150 VSSD.n691 VSSD.n690 9.3005
R12151 VSSD.n692 VSSD.n547 9.3005
R12152 VSSD.n694 VSSD.n693 9.3005
R12153 VSSD.n696 VSSD.n695 9.3005
R12154 VSSD.n701 VSSD.n700 9.3005
R12155 VSSD.n702 VSSD.n545 9.3005
R12156 VSSD.n704 VSSD.n703 9.3005
R12157 VSSD.n705 VSSD.n541 9.3005
R12158 VSSD.n706 VSSD.n542 9.3005
R12159 VSSD.n723 VSSD.n722 9.3005
R12160 VSSD.n721 VSSD.n720 9.3005
R12161 VSSD.n719 VSSD.n718 9.3005
R12162 VSSD.n716 VSSD.n708 9.3005
R12163 VSSD.n715 VSSD.n714 9.3005
R12164 VSSD VSSD.n712 9.3005
R12165 VSSD.n713 VSSD.n44 9.3005
R12166 VSSD.n3669 VSSD.n45 9.3005
R12167 VSSD.n3671 VSSD.n3670 9.3005
R12168 VSSD.n3673 VSSD.n3672 9.3005
R12169 VSSD.n3676 VSSD.n40 9.3005
R12170 VSSD.n3680 VSSD.n3679 9.3005
R12171 VSSD.n3682 VSSD.n3681 9.3005
R12172 VSSD.n3683 VSSD.n38 9.3005
R12173 VSSD.n3685 VSSD.n3684 9.3005
R12174 VSSD.n3686 VSSD.n37 9.3005
R12175 VSSD.n3688 VSSD.n3687 9.3005
R12176 VSSD.n3689 VSSD.n36 9.3005
R12177 VSSD.n3693 VSSD.n3692 9.3005
R12178 VSSD.n3695 VSSD.n3694 9.3005
R12179 VSSD.n3697 VSSD.n3696 9.3005
R12180 VSSD.n24 VSSD.n23 9.3005
R12181 VSSD.n3708 VSSD.n3707 9.3005
R12182 VSSD.n3714 VSSD.n3713 9.3005
R12183 VSSD.n3715 VSSD.n21 9.3005
R12184 VSSD.n3717 VSSD.n3716 9.3005
R12185 VSSD.n3718 VSSD.n20 9.3005
R12186 VSSD.n3720 VSSD.n3719 9.3005
R12187 VSSD.n3721 VSSD.n19 9.3005
R12188 VSSD.n3723 VSSD.n3722 9.3005
R12189 VSSD.n3724 VSSD.n18 9.3005
R12190 VSSD.n3726 VSSD.n3725 9.3005
R12191 VSSD.n3727 VSSD.n17 9.3005
R12192 VSSD.n3729 VSSD.n3728 9.3005
R12193 VSSD.n3733 VSSD.n3732 9.3005
R12194 VSSD.n3734 VSSD.n15 9.3005
R12195 VSSD.n3736 VSSD.n3735 9.3005
R12196 VSSD.n3739 VSSD.n3738 9.3005
R12197 VSSD.n3740 VSSD.n14 9.3005
R12198 VSSD.n3742 VSSD.n3741 9.3005
R12199 VSSD.n3744 VSSD.n12 9.3005
R12200 VSSD.n3746 VSSD.n3745 9.3005
R12201 VSSD.n3747 VSSD.n11 9.3005
R12202 VSSD.n3749 VSSD.n3748 9.3005
R12203 VSSD.n3750 VSSD.n10 9.3005
R12204 VSSD.n3753 VSSD.n3752 9.3005
R12205 VSSD.n3755 VSSD.n3754 9.3005
R12206 VSSD.n3756 VSSD.n8 9.3005
R12207 VSSD.n3762 VSSD.n3761 9.3005
R12208 VSSD.n251 VSSD.n247 9.29365
R12209 VSSD.n1252 VSSD.n1251 9.18349
R12210 VSSD.n2091 VSSD.n2090 9.03579
R12211 VSSD.n1783 VSSD.n1782 9.03579
R12212 VSSD.n1669 VSSD.n1666 9.03579
R12213 VSSD.n3008 VSSD.n3007 8.54503
R12214 VSSD.t495 VSSD.t1150 8.42962
R12215 VSSD.t530 VSSD.t475 8.42962
R12216 VSSD.t1629 VSSD 8.42962
R12217 VSSD.t847 VSSD 8.42962
R12218 VSSD.t260 VSSD.t987 8.42962
R12219 VSSD.t1137 VSSD.t288 8.42962
R12220 VSSD VSSD.t556 8.42962
R12221 VSSD VSSD.t1092 8.42962
R12222 VSSD.t1108 VSSD 8.42962
R12223 VSSD.t67 VSSD.t256 8.42962
R12224 VSSD.t64 VSSD.t125 8.42962
R12225 VSSD.t1797 VSSD.t476 8.42962
R12226 VSSD.n872 VSSD.n870 8.28285
R12227 VSSD.n2132 VSSD.n2129 8.259
R12228 VSSD.n3233 VSSD.n3232 8.24457
R12229 VSSD.n2698 VSSD.n2697 8.24457
R12230 VSSD.n1764 VSSD.n1763 8.24457
R12231 VSSD.n704 VSSD.n545 8.23546
R12232 VSSD.n705 VSSD.n704 8.23546
R12233 VSSD.n706 VSSD.n705 8.23546
R12234 VSSD.n722 VSSD.n706 8.23546
R12235 VSSD.n722 VSSD.n721 8.23546
R12236 VSSD.n716 VSSD.n715 8.23546
R12237 VSSD.n685 VSSD.n551 8.23546
R12238 VSSD.n686 VSSD.n685 8.23546
R12239 VSSD.n688 VSSD.n686 8.23546
R12240 VSSD.n692 VSSD.n691 8.23546
R12241 VSSD.n693 VSSD.n692 8.23546
R12242 VSSD.n954 VSSD.n953 8.23546
R12243 VSSD.n950 VSSD.n949 8.23546
R12244 VSSD.n949 VSSD.n948 8.23546
R12245 VSSD.n948 VSSD.n861 8.23546
R12246 VSSD.n941 VSSD.n940 8.23546
R12247 VSSD.n3369 VSSD.n3368 8.23546
R12248 VSSD.n3368 VSSD.n516 8.23546
R12249 VSSD.n3364 VSSD.n516 8.23546
R12250 VSSD.n3361 VSSD.n3360 8.23546
R12251 VSSD.n3360 VSSD.n519 8.23546
R12252 VSSD.n3297 VSSD.n3296 8.23546
R12253 VSSD.n3294 VSSD.n3236 8.23546
R12254 VSSD.n3290 VSSD.n3236 8.23546
R12255 VSSD.n3290 VSSD.n3289 8.23546
R12256 VSSD.n3289 VSSD.n3288 8.23546
R12257 VSSD.n3283 VSSD.n3282 8.23546
R12258 VSSD.n3273 VSSD.n3272 8.23546
R12259 VSSD.n3272 VSSD.n3245 8.23546
R12260 VSSD.n3268 VSSD.n3245 8.23546
R12261 VSSD.n2912 VSSD.n2911 8.23546
R12262 VSSD.n2912 VSSD.n1120 8.23546
R12263 VSSD.n2916 VSSD.n1120 8.23546
R12264 VSSD.n2917 VSSD.n2916 8.23546
R12265 VSSD.n2923 VSSD.n2922 8.23546
R12266 VSSD.n2924 VSSD.n2923 8.23546
R12267 VSSD.n2784 VSSD.n2783 8.23546
R12268 VSSD.n2783 VSSD.n1367 8.23546
R12269 VSSD.n2779 VSSD.n1367 8.23546
R12270 VSSD.n2772 VSSD.n2771 8.23546
R12271 VSSD.n2771 VSSD.n2770 8.23546
R12272 VSSD.n2762 VSSD.n2761 8.23546
R12273 VSSD.n2759 VSSD.n2701 8.23546
R12274 VSSD.n2755 VSSD.n2701 8.23546
R12275 VSSD.n2755 VSSD.n2754 8.23546
R12276 VSSD.n2754 VSSD.n2753 8.23546
R12277 VSSD.n2748 VSSD.n2747 8.23546
R12278 VSSD.n2738 VSSD.n2737 8.23546
R12279 VSSD.n2737 VSSD.n2710 8.23546
R12280 VSSD.n2733 VSSD.n2710 8.23546
R12281 VSSD.n2448 VSSD.n2447 8.23546
R12282 VSSD.n2447 VSSD.n2446 8.23546
R12283 VSSD.n2446 VSSD.n2389 8.23546
R12284 VSSD.n2442 VSSD.n2389 8.23546
R12285 VSSD.n2442 VSSD.n2441 8.23546
R12286 VSSD.n2436 VSSD.n2435 8.23546
R12287 VSSD.n2435 VSSD.n2434 8.23546
R12288 VSSD.n2425 VSSD.n2424 8.23546
R12289 VSSD.n2424 VSSD.n2423 8.23546
R12290 VSSD.n2071 VSSD.n2070 8.23546
R12291 VSSD.n2070 VSSD.n2069 8.23546
R12292 VSSD.n1737 VSSD.n1736 8.23546
R12293 VSSD.n1736 VSSD.n1709 8.23546
R12294 VSSD.n1732 VSSD.n1709 8.23546
R12295 VSSD.n1761 VSSD.n1697 8.23546
R12296 VSSD.n1757 VSSD.n1756 8.23546
R12297 VSSD.n1756 VSSD.n1755 8.23546
R12298 VSSD.n1755 VSSD.n1701 8.23546
R12299 VSSD.n1751 VSSD.n1701 8.23546
R12300 VSSD.n1747 VSSD.n1704 8.23546
R12301 VSSD.n1945 VSSD.n1576 8.23546
R12302 VSSD.n1934 VSSD.n1933 8.23546
R12303 VSSD.n1933 VSSD.n1932 8.23546
R12304 VSSD.n1932 VSSD.n1580 8.23546
R12305 VSSD.n1928 VSSD.n1580 8.23546
R12306 VSSD.n1925 VSSD.n1924 8.23546
R12307 VSSD.n1924 VSSD.n1583 8.23546
R12308 VSSD.n1914 VSSD.n1913 8.23546
R12309 VSSD.n1913 VSSD.n1587 8.23546
R12310 VSSD.n3429 VSSD.n3428 8.23546
R12311 VSSD.n3430 VSSD.n3429 8.23546
R12312 VSSD.n3430 VSSD.n118 8.23546
R12313 VSSD.n3434 VSSD.n118 8.23546
R12314 VSSD.n3435 VSSD.n3434 8.23546
R12315 VSSD.n3436 VSSD.n3435 8.23546
R12316 VSSD.n3440 VSSD.n3439 8.23546
R12317 VSSD.n3441 VSSD.n3440 8.23546
R12318 VSSD.n3449 VSSD.n3448 8.23546
R12319 VSSD.n3450 VSSD.n3449 8.23546
R12320 VSSD.n3450 VSSD.n111 8.23546
R12321 VSSD.n3454 VSSD.n111 8.23546
R12322 VSSD.n3455 VSSD.n3454 8.23546
R12323 VSSD.n3456 VSSD.n3455 8.23546
R12324 VSSD.n3460 VSSD.n3459 8.23546
R12325 VSSD.n3462 VSSD.n3460 8.23546
R12326 VSSD.n3485 VSSD.n3484 8.23546
R12327 VSSD.n3486 VSSD.n3485 8.23546
R12328 VSSD.n3486 VSSD.n90 8.23546
R12329 VSSD.n3490 VSSD.n90 8.23546
R12330 VSSD.n3491 VSSD.n3490 8.23546
R12331 VSSD.n3492 VSSD.n3491 8.23546
R12332 VSSD.n3496 VSSD.n3495 8.23546
R12333 VSSD.n3497 VSSD.n3496 8.23546
R12334 VSSD.n3506 VSSD.n85 8.23546
R12335 VSSD.n3507 VSSD.n3506 8.23546
R12336 VSSD.n3507 VSSD.n77 8.23546
R12337 VSSD.n3522 VSSD.n77 8.23546
R12338 VSSD.n3523 VSSD.n3522 8.23546
R12339 VSSD.n3524 VSSD.n3523 8.23546
R12340 VSSD.n3528 VSSD.n3527 8.23546
R12341 VSSD.n3530 VSSD.n3528 8.23546
R12342 VSSD.n3546 VSSD.n3545 8.23546
R12343 VSSD.n3547 VSSD.n3546 8.23546
R12344 VSSD.n3547 VSSD.n67 8.23546
R12345 VSSD.n3551 VSSD.n67 8.23546
R12346 VSSD.n3552 VSSD.n3551 8.23546
R12347 VSSD.n3553 VSSD.n3552 8.23546
R12348 VSSD.n3559 VSSD.n3556 8.23546
R12349 VSSD.n3559 VSSD.n3558 8.23546
R12350 VSSD.n3575 VSSD.n3574 8.23546
R12351 VSSD.n3576 VSSD.n3575 8.23546
R12352 VSSD.n3576 VSSD.n51 8.23546
R12353 VSSD.n3580 VSSD.n51 8.23546
R12354 VSSD.n3581 VSSD.n3580 8.23546
R12355 VSSD.n3582 VSSD.n3581 8.23546
R12356 VSSD.n3586 VSSD.n3585 8.23546
R12357 VSSD.n3588 VSSD.n3586 8.23546
R12358 VSSD.n3651 VSSD.n3650 8.23546
R12359 VSSD.n3650 VSSD.n3649 8.23546
R12360 VSSD.n3649 VSSD.n3595 8.23546
R12361 VSSD.n3645 VSSD.n3595 8.23546
R12362 VSSD.n3645 VSSD.n3644 8.23546
R12363 VSSD.n3644 VSSD.n3643 8.23546
R12364 VSSD.n3640 VSSD.n3639 8.23546
R12365 VSSD.n3639 VSSD.n3638 8.23546
R12366 VSSD.n3631 VSSD.n3630 8.23546
R12367 VSSD.n3630 VSSD.n3629 8.23546
R12368 VSSD.n3629 VSSD.n3602 8.23546
R12369 VSSD.n3625 VSSD.n3602 8.23546
R12370 VSSD.n3625 VSSD.n3624 8.23546
R12371 VSSD.n3624 VSSD.n3623 8.23546
R12372 VSSD.n3620 VSSD.n3619 8.23546
R12373 VSSD.n3619 VSSD.n3618 8.23546
R12374 VSSD.n330 VSSD.n329 8.23546
R12375 VSSD.n329 VSSD.n242 8.23546
R12376 VSSD.n3742 VSSD.n14 8.23546
R12377 VSSD.n3745 VSSD.n3744 8.23546
R12378 VSSD.n3745 VSSD.n11 8.23546
R12379 VSSD.n3749 VSSD.n11 8.23546
R12380 VSSD.n3750 VSSD.n3749 8.23546
R12381 VSSD.n3756 VSSD.n3755 8.23546
R12382 VSSD.n3376 VSSD.n512 8.16157
R12383 VSSD.n785 VSSD.n783 8.10717
R12384 VSSD.n3018 VSSD.n3016 8.10717
R12385 VSSD.n3674 VSSD.n42 8.10717
R12386 VSSD.n3760 VSSD.n3759 8.10717
R12387 VSSD.n712 VSSD.n710 8.05644
R12388 VSSD.n2288 VSSD.n1440 8.05644
R12389 VSSD.n2286 VSSD.n1444 8.05644
R12390 VSSD.n1909 VSSD.n1589 8.05644
R12391 VSSD.n921 VSSD.n920 7.90638
R12392 VSSD.n914 VSSD.n913 7.90638
R12393 VSSD.n3192 VSSD.n3191 7.90638
R12394 VSSD.n1187 VSSD.n1161 7.90638
R12395 VSSD.n2976 VSSD.n2973 7.90638
R12396 VSSD.n2985 VSSD.n1088 7.90638
R12397 VSSD.n3136 VSSD.n3135 7.90638
R12398 VSSD.n3134 VSSD.n3133 7.90638
R12399 VSSD.n3099 VSSD.n3098 7.90638
R12400 VSSD.n2603 VSSD.n2602 7.90638
R12401 VSSD.n2606 VSSD.n2605 7.90638
R12402 VSSD.n2360 VSSD.n2358 7.90638
R12403 VSSD.n1544 VSSD.n1503 7.90638
R12404 VSSD.n1542 VSSD.n1541 7.90638
R12405 VSSD.n2002 VSSD.n1463 7.90638
R12406 VSSD.n2000 VSSD.n1999 7.90638
R12407 VSSD.n2198 VSSD.n2197 7.90638
R12408 VSSD.n2154 VSSD.n2151 7.90638
R12409 VSSD.n1805 VSSD.n1803 7.90638
R12410 VSSD.n1793 VSSD.n1792 7.90638
R12411 VSSD.n1862 VSSD.n1635 7.90638
R12412 VSSD.n460 VSSD.n458 7.90638
R12413 VSSD.n463 VSSD.n461 7.90638
R12414 VSSD.n401 VSSD.n400 7.90638
R12415 VSSD.n400 VSSD.n399 7.90638
R12416 VSSD.n347 VSSD.n224 7.90638
R12417 VSSD.n3691 VSSD.n3689 7.90638
R12418 VSSD.n3712 VSSD.n21 7.90638
R12419 VSSD.n681 VSSD.n680 7.87742
R12420 VSSD.n3371 VSSD.n3370 7.87742
R12421 VSSD.n944 VSSD.n863 7.78791
R12422 VSSD.n3267 VSSD.n3266 7.78791
R12423 VSSD.n2778 VSSD.n2777 7.78791
R12424 VSSD.n2732 VSSD.n2731 7.78791
R12425 VSSD.n2420 VSSD.n2397 7.78791
R12426 VSSD.n1731 VSSD.n1730 7.78791
R12427 VSSD.n325 VSSD.n244 7.78791
R12428 VSSD.n1206 VSSD.n1205 7.73676
R12429 VSSD.n712 VSSD.n711 7.6984
R12430 VSSD.n681 VSSD.n679 7.6984
R12431 VSSD.n693 VSSD.n546 7.6984
R12432 VSSD.n955 VSSD.n954 7.6984
R12433 VSSD.n937 VSSD.n864 7.6984
R12434 VSSD.n937 VSSD.n936 7.6984
R12435 VSSD.n3371 VSSD.n514 7.6984
R12436 VSSD.n520 VSSD.n519 7.6984
R12437 VSSD.n3297 VSSD.n3235 7.6984
R12438 VSSD.n3282 VSSD.n3241 7.6984
R12439 VSSD.n3275 VSSD.n3242 7.6984
R12440 VSSD.n3266 VSSD.n3265 7.6984
R12441 VSSD.n2909 VSSD.n1123 7.6984
R12442 VSSD.n2924 VSSD.n1115 7.6984
R12443 VSSD.n2786 VSSD.n1364 7.6984
R12444 VSSD.n2777 VSSD.n2776 7.6984
R12445 VSSD.n2770 VSSD.n2695 7.6984
R12446 VSSD.n2762 VSSD.n2700 7.6984
R12447 VSSD.n2747 VSSD.n2706 7.6984
R12448 VSSD.n2740 VSSD.n2707 7.6984
R12449 VSSD.n2731 VSSD.n2730 7.6984
R12450 VSSD.n2434 VSSD.n2394 7.6984
R12451 VSSD.n2425 VSSD.n2395 7.6984
R12452 VSSD.n2420 VSSD.n2419 7.6984
R12453 VSSD.n2073 VSSD.n2068 7.6984
R12454 VSSD.n2283 VSSD.n2282 7.6984
R12455 VSSD.n1739 VSSD.n1706 7.6984
R12456 VSSD.n1730 VSSD.n1729 7.6984
R12457 VSSD.n1762 VSSD.n1761 7.6984
R12458 VSSD.n1705 VSSD.n1704 7.6984
R12459 VSSD.n1946 VSSD.n1945 7.6984
R12460 VSSD.n1584 VSSD.n1583 7.6984
R12461 VSSD.n1916 VSSD.n1585 7.6984
R12462 VSSD.n3428 VSSD.n120 7.6984
R12463 VSSD.n3441 VSSD.n114 7.6984
R12464 VSSD.n3448 VSSD.n113 7.6984
R12465 VSSD.n3462 VSSD.n3461 7.6984
R12466 VSSD.n3484 VSSD.n92 7.6984
R12467 VSSD.n3497 VSSD.n86 7.6984
R12468 VSSD.n3501 VSSD.n85 7.6984
R12469 VSSD.n3530 VSSD.n3529 7.6984
R12470 VSSD.n3545 VSSD.n69 7.6984
R12471 VSSD.n3558 VSSD.n54 7.6984
R12472 VSSD.n3574 VSSD.n53 7.6984
R12473 VSSD.n3588 VSSD.n3587 7.6984
R12474 VSSD.n3651 VSSD.n3594 7.6984
R12475 VSSD.n3638 VSSD.n3599 7.6984
R12476 VSSD.n3631 VSSD.n3600 7.6984
R12477 VSSD.n3618 VSSD.n3606 7.6984
R12478 VSSD.n331 VSSD.n330 7.6984
R12479 VSSD.n325 VSSD.n324 7.6984
R12480 VSSD.n3737 VSSD.n14 7.6984
R12481 VSSD.n3757 VSSD.n3756 7.6984
R12482 VSSD.n1514 VSSD.n1513 7.6005
R12483 VSSD.n3765 VSSD.n3764 7.5961
R12484 VSSD.n2966 VSSD.n1094 7.52991
R12485 VSSD.n2667 VSSD.n2666 7.52991
R12486 VSSD.n2339 VSSD.n2338 7.52991
R12487 VSSD.n1531 VSSD.n1509 7.52991
R12488 VSSD.n2015 VSSD.n2014 7.52991
R12489 VSSD.n2099 VSSD.n2098 7.52991
R12490 VSSD.n2280 VSSD.n2108 7.52991
R12491 VSSD.n2207 VSSD.n2206 7.52991
R12492 VSSD.n411 VSSD.n185 7.52991
R12493 VSSD.n389 VSSD.n198 7.52991
R12494 VSSD.n357 VSSD.n356 7.52991
R12495 VSSD.n2874 VSSD.n2873 7.23528
R12496 VSSD.n1619 VSSD.n1618 7.16134
R12497 VSSD.n2832 VSSD.n1326 7.15344
R12498 VSSD.n673 VSSD.n556 7.11268
R12499 VSSD.n1294 VSSD.n1147 6.88949
R12500 VSSD.n2418 VSSD.n2417 6.88949
R12501 VSSD.n1909 VSSD.n1908 6.88949
R12502 VSSD.n1900 VSSD.n1592 6.88949
R12503 VSSD.n323 VSSD.n322 6.88949
R12504 VSSD.n1001 VSSD.n1000 6.77697
R12505 VSSD.n1258 VSSD.n1247 6.77697
R12506 VSSD.n2928 VSSD.n1114 6.77697
R12507 VSSD.n2940 VSSD.n2934 6.77697
R12508 VSSD.n311 VSSD.n252 6.6092
R12509 VSSD.n666 VSSD.n665 6.57117
R12510 VSSD.n721 VSSD.n707 6.44526
R12511 VSSD.n3295 VSSD.n3294 6.44526
R12512 VSSD.n2760 VSSD.n2759 6.44526
R12513 VSSD.n2448 VSSD.n2388 6.44526
R12514 VSSD.n2073 VSSD.n2072 6.44526
R12515 VSSD.n1757 VSSD.n1700 6.44526
R12516 VSSD.n1916 VSSD.n1915 6.44526
R12517 VSSD.n3752 VSSD.n9 6.44526
R12518 VSSD.n666 VSSD.n568 6.4005
R12519 VSSD.n2953 VSSD.n1098 6.4005
R12520 VSSD.n2503 VSSD.n1388 6.4005
R12521 VSSD.n1841 VSSD.n1840 6.26433
R12522 VSSD.n900 VSSD.n899 6.26433
R12523 VSSD.n993 VSSD.n992 6.26433
R12524 VSSD.n796 VSSD.n795 6.26433
R12525 VSSD.n795 VSSD.n794 6.26433
R12526 VSSD.n3318 VSSD.n1024 6.26433
R12527 VSSD.n2875 VSSD.n2871 6.26433
R12528 VSSD.n2883 VSSD.n2882 6.26433
R12529 VSSD.n3054 VSSD.n1078 6.26433
R12530 VSSD.n2828 VSSD.n2827 6.26433
R12531 VSSD.n2568 VSSD.n2567 6.26433
R12532 VSSD.n2793 VSSD.n1363 6.26433
R12533 VSSD.n2376 VSSD.n2375 6.26433
R12534 VSSD.n2273 VSSD.n2272 6.26433
R12535 VSSD.n2272 VSSD.n2271 6.26433
R12536 VSSD.n2229 VSSD.n2228 6.26433
R12537 VSSD.n2228 VSSD.n2133 6.26433
R12538 VSSD.n2173 VSSD.n2172 6.26433
R12539 VSSD.n1770 VSSD.n1769 6.26433
R12540 VSSD.n1829 VSSD.n1828 6.26433
R12541 VSSD.n1828 VSSD.n1658 6.26433
R12542 VSSD.n1840 VSSD.n1654 6.26433
R12543 VSSD.n1843 VSSD.n1651 6.26433
R12544 VSSD.n3679 VSSD.n3676 6.26433
R12545 VSSD.n896 VSSD.n886 6.12816
R12546 VSSD.n1842 VSSD.n1841 6.12816
R12547 VSSD.n635 VSSD.n634 6.02861
R12548 VSSD.n624 VSSD.n623 6.02861
R12549 VSSD.n2671 VSSD.n2637 6.02403
R12550 VSSD.n2675 VSSD.n2637 6.02403
R12551 VSSD.n2680 VSSD.n2678 6.02403
R12552 VSSD.n2684 VSSD.n2634 6.02403
R12553 VSSD.n1883 VSSD.n1882 6.02403
R12554 VSSD.n983 VSSD.n830 5.98311
R12555 VSSD.n805 VSSD.n804 5.98311
R12556 VSSD.n1296 VSSD.n1139 5.98311
R12557 VSSD.n3013 VSSD.n1080 5.98311
R12558 VSSD.n3403 VSSD.n3402 5.98311
R12559 VSSD.n3412 VSSD.n3410 5.98311
R12560 VSSD.n3477 VSSD.n3475 5.98311
R12561 VSSD.n3538 VSSD.n3536 5.98311
R12562 VSSD.n3611 VSSD.n3607 5.98311
R12563 VSSD.n1774 VSSD.n1773 5.9239
R12564 VSSD.n950 VSSD.n859 5.90819
R12565 VSSD.n3274 VSSD.n3273 5.90819
R12566 VSSD.n2910 VSSD.n2909 5.90819
R12567 VSSD.n2785 VSSD.n2784 5.90819
R12568 VSSD.n2739 VSSD.n2738 5.90819
R12569 VSSD.n1738 VSSD.n1737 5.90819
R12570 VSSD.n1579 VSSD.n1576 5.90819
R12571 VSSD.n1654 VSSD.n1653 5.8885
R12572 VSSD.n901 VSSD.n900 5.85582
R12573 VSSD.n994 VSSD.n993 5.85582
R12574 VSSD.n796 VSSD.n776 5.85582
R12575 VSSD.n3388 VSSD.n491 5.85582
R12576 VSSD.n3168 VSSD.n3160 5.85582
R12577 VSSD.n3320 VSSD.n1022 5.85582
R12578 VSSD.n2871 VSSD.n2870 5.85582
R12579 VSSD.n3054 VSSD.n1077 5.85582
R12580 VSSD.n2828 VSSD.n1327 5.85582
R12581 VSSD.n2567 VSSD.n2558 5.85582
R12582 VSSD.n2325 VSSD.n2317 5.85582
R12583 VSSD.n2375 VSSD.n1419 5.85582
R12584 VSSD.n2463 VSSD.n2462 5.85582
R12585 VSSD.n1524 VSSD.n1515 5.85582
R12586 VSSD.n2023 VSSD.n2022 5.85582
R12587 VSSD.n2273 VSSD.n2109 5.85582
R12588 VSSD.n2230 VSSD.n2229 5.85582
R12589 VSSD.n1776 VSSD.n1775 5.85582
R12590 VSSD.n1773 VSSD.n1692 5.85582
R12591 VSSD.n1769 VSSD.n1694 5.85582
R12592 VSSD.n1651 VSSD.n1650 5.85582
R12593 VSSD.n1612 VSSD.n1599 5.85582
R12594 VSSD.n1611 VSSD.n1610 5.85582
R12595 VSSD.n371 VSSD.n212 5.85582
R12596 VSSD.n3676 VSSD.n3675 5.85582
R12597 VSSD.n794 VSSD.n777 5.65809
R12598 VSSD.n2895 VSSD.n1128 5.65809
R12599 VSSD.n2271 VSSD.n2111 5.65809
R12600 VSSD.n2224 VSSD.n2133 5.65809
R12601 VSSD.n678 VSSD.n677 5.63966
R12602 VSSD.n674 VSSD.n673 5.63966
R12603 VSSD.n3375 VSSD.n3374 5.63966
R12604 VSSD.n1294 VSSD.n1148 5.63966
R12605 VSSD.n2288 VSSD.n2287 5.63966
R12606 VSSD.n2287 VSSD.n2286 5.63966
R12607 VSSD.n3773 VSSD.n3772 5.56058
R12608 VSSD.n1286 VSSD.n1231 5.53969
R12609 VSSD.n2872 VSSD.n2859 5.51774
R12610 VSSD.n646 VSSD.n645 5.48128
R12611 VSSD.n3228 VSSD.n3227 5.47626
R12612 VSSD.n3178 VSSD.n3157 5.47626
R12613 VSSD.n2162 VSSD.n2161 5.44731
R12614 VSSD.n3387 VSSD.n499 5.38843
R12615 VSSD.n3169 VSSD.n3168 5.37524
R12616 VSSD.n3050 VSSD.n1078 5.37524
R12617 VSSD.n1524 VSSD.n1523 5.37524
R12618 VSSD.n3184 VSSD.n3154 5.35702
R12619 VSSD.n3302 VSSD.n3230 5.35702
R12620 VSSD.n1824 VSSD.n1660 5.24958
R12621 VSSD.n563 VSSD.n561 5.13108
R12622 VSSD.n563 VSSD.n562 5.13108
R12623 VSSD.n555 VSSD.n554 5.13108
R12624 VSSD.n889 VSSD.n887 5.13108
R12625 VSSD.n889 VSSD.n888 5.13108
R12626 VSSD.n495 VSSD.n492 5.13108
R12627 VSSD.n495 VSSD.n494 5.13108
R12628 VSSD.n1229 VSSD.n1228 5.13108
R12629 VSSD.n1143 VSSD.n1140 5.13108
R12630 VSSD.n1143 VSSD.n1142 5.13108
R12631 VSSD.n3254 VSSD.n3251 5.13108
R12632 VSSD.n3254 VSSD.n3252 5.13108
R12633 VSSD.n2865 VSSD.n2863 5.13108
R12634 VSSD.n2865 VSSD.n2864 5.13108
R12635 VSSD.n3080 VSSD.n3077 5.13108
R12636 VSSD.n3080 VSSD.n3078 5.13108
R12637 VSSD.n2562 VSSD.n2559 5.13108
R12638 VSSD.n2562 VSSD.n2561 5.13108
R12639 VSSD.n2719 VSSD.n2716 5.13108
R12640 VSSD.n2719 VSSD.n2717 5.13108
R12641 VSSD.n1485 VSSD.n1483 5.13108
R12642 VSSD.n1485 VSSD.n1484 5.13108
R12643 VSSD.n2406 VSSD.n2403 5.13108
R12644 VSSD.n2406 VSSD.n2404 5.13108
R12645 VSSD.n1966 VSSD.n1964 5.13108
R12646 VSSD.n1966 VSSD.n1965 5.13108
R12647 VSSD.n1442 VSSD.n1441 5.13108
R12648 VSSD.n2168 VSSD.n2165 5.13108
R12649 VSSD.n2168 VSSD.n2166 5.13108
R12650 VSSD.n1718 VSSD.n1715 5.13108
R12651 VSSD.n1718 VSSD.n1717 5.13108
R12652 VSSD.n1602 VSSD.n1600 5.13108
R12653 VSSD.n1602 VSSD.n1601 5.13108
R12654 VSSD.n270 VSSD.n267 5.13108
R12655 VSSD.n270 VSSD.n268 5.13108
R12656 VSSD.n136 VSSD.n134 5.13108
R12657 VSSD.n136 VSSD.n135 5.13108
R12658 VSSD.n3790 VSSD.n3788 5.13108
R12659 VSSD.n3790 VSSD.n3789 5.13108
R12660 VSSD.n2027 VSSD.n2024 4.97071
R12661 VSSD.n1836 VSSD.n1655 4.97071
R12662 VSSD.n2327 VSSD.n2326 4.90263
R12663 VSSD.n370 VSSD.n369 4.90263
R12664 VSSD.n652 VSSD.n651 4.85762
R12665 VSSD.n788 VSSD.n781 4.85762
R12666 VSSD.n1277 VSSD.n1276 4.85762
R12667 VSSD.n3312 VSSD.n3311 4.85762
R12668 VSSD.n2900 VSSD.n1127 4.85762
R12669 VSSD.n2222 VSSD.n2221 4.85762
R12670 VSSD.n2265 VSSD.n2117 4.85762
R12671 VSSD.n1822 VSSD.n1821 4.85762
R12672 VSSD.n420 VSSD.n179 4.85762
R12673 VSSD.n698 VSSD.n545 4.83407
R12674 VSSD.n3285 VSSD.n3284 4.83407
R12675 VSSD.n2919 VSSD.n2918 4.83407
R12676 VSSD.n2750 VSSD.n2749 4.83407
R12677 VSSD.n2441 VSSD.n2440 4.83407
R12678 VSSD.n1749 VSSD.n1748 4.83407
R12679 VSSD.n3744 VSSD.n3743 4.83407
R12680 VSSD.n983 VSSD.n982 4.8005
R12681 VSSD.n1297 VSSD.n1296 4.8005
R12682 VSSD.n3014 VSSD.n3013 4.8005
R12683 VSSD.n3402 VSSD.n3401 4.8005
R12684 VSSD.n3412 VSSD.n3411 4.8005
R12685 VSSD.n3477 VSSD.n3476 4.8005
R12686 VSSD.n3538 VSSD.n3537 4.8005
R12687 VSSD.n3611 VSSD.n3610 4.8005
R12688 VSSD.n676 VSSD.n675 4.72533
R12689 VSSD.n3376 VSSD.n3375 4.72533
R12690 VSSD.n640 VSSD.n639 4.67352
R12691 VSSD.n639 VSSD.n588 4.67352
R12692 VSSD.n629 VSSD.n628 4.67352
R12693 VSSD.n628 VSSD.n592 4.67352
R12694 VSSD.n618 VSSD.n617 4.67352
R12695 VSSD.n617 VSSD.n597 4.67352
R12696 VSSD.n307 VSSD.n306 4.67352
R12697 VSSD.n306 VSSD.n305 4.67352
R12698 VSSD.n305 VSSD.n255 4.67352
R12699 VSSD.n301 VSSD.n255 4.67352
R12700 VSSD.n301 VSSD.n300 4.67352
R12701 VSSD.n300 VSSD.n299 4.67352
R12702 VSSD.n296 VSSD.n295 4.67352
R12703 VSSD.n295 VSSD.n294 4.67352
R12704 VSSD.n287 VSSD.n286 4.67352
R12705 VSSD.n286 VSSD.n285 4.67352
R12706 VSSD.n285 VSSD.n262 4.67352
R12707 VSSD.n281 VSSD.n262 4.67352
R12708 VSSD.n281 VSSD.n280 4.67352
R12709 VSSD.n280 VSSD.n279 4.67352
R12710 VSSD.n276 VSSD.n275 4.67352
R12711 VSSD.n275 VSSD.n274 4.67352
R12712 VSSD.n677 VSSD.n676 4.63943
R12713 VSSD.n2572 VSSD.n2570 4.62124
R12714 VSSD.n314 VSSD.n313 4.62124
R12715 VSSD.n667 VSSD.n666 4.62124
R12716 VSSD.n676 VSSD.n553 4.62124
R12717 VSSD.n2668 VSSD.n2667 4.51815
R12718 VSSD.n2104 VSSD.n2103 4.51815
R12719 VSSD.n2093 VSSD.n2052 4.51815
R12720 VSSD.n577 VSSD.n566 4.51401
R12721 VSSD.n657 VSSD.n656 4.51401
R12722 VSSD.n600 VSSD.n598 4.51401
R12723 VSSD.n608 VSSD.n607 4.51401
R12724 VSSD.n167 VSSD.n164 4.51401
R12725 VSSD.n425 VSSD.n424 4.51401
R12726 VSSD.n732 VSSD.n539 4.51401
R12727 VSSD.n544 VSSD.n543 4.51401
R12728 VSSD.n202 VSSD.n197 4.51401
R12729 VSSD.n379 VSSD.n378 4.51401
R12730 VSSD.n3700 VSSD.n30 4.51401
R12731 VSSD.n3704 VSSD.n22 4.51401
R12732 VSSD.n1011 VSSD.n737 4.51401
R12733 VSSD.n744 VSSD.n741 4.51401
R12734 VSSD.n3340 VSSD.n3339 4.51401
R12735 VSSD.n767 VSSD.n766 4.51401
R12736 VSSD.n508 VSSD.n506 4.51401
R12737 VSSD.n3379 VSSD.n3378 4.51401
R12738 VSSD.n965 VSSD.n964 4.51401
R12739 VSSD.n959 VSSD.n958 4.51401
R12740 VSSD.n3330 VSSD 4.51401
R12741 VSSD.n1021 VSSD.n1020 4.51401
R12742 VSSD.n1212 VSSD.n1211 4.51401
R12743 VSSD.n1227 VSSD.n1226 4.51401
R12744 VSSD.n1308 VSSD.n1134 4.51401
R12745 VSSD.n1174 VSSD.n1173 4.51401
R12746 VSSD.n3197 VSSD.n3152 4.51401
R12747 VSSD.n3202 VSSD.n3201 4.51401
R12748 VSSD.n2992 VSSD.n2991 4.51401
R12749 VSSD.n3004 VSSD.n3003 4.51401
R12750 VSSD.n2944 VSSD.n1106 4.51401
R12751 VSSD.n2949 VSSD.n2948 4.51401
R12752 VSSD.n2887 VSSD.n2854 4.51401
R12753 VSSD.n2892 VSSD.n2891 4.51401
R12754 VSSD.n3148 VSSD.n1056 4.51401
R12755 VSSD.n3139 VSSD.n3138 4.51401
R12756 VSSD.n2846 VSSD.n1316 4.51401
R12757 VSSD.n1321 VSSD.n1320 4.51401
R12758 VSSD.n2624 VSSD.n2528 4.51401
R12759 VSSD.n2629 VSSD.n2628 4.51401
R12760 VSSD.n2557 VSSD.n2556 4.51401
R12761 VSSD.n2580 VSSD.n2579 4.51401
R12762 VSSD.n1354 VSSD.n1346 4.51401
R12763 VSSD.n2796 VSSD.n2795 4.51401
R12764 VSSD.n1402 VSSD.n1397 4.51401
R12765 VSSD.n2467 VSSD.n2466 4.51401
R12766 VSSD.n2524 VSSD.n1377 4.51401
R12767 VSSD.n2516 VSSD.n2515 4.51401
R12768 VSSD.n1566 VSSD.n1476 4.51401
R12769 VSSD.n1556 VSSD.n1552 4.51401
R12770 VSSD.n2348 VSSD.n2306 4.51401
R12771 VSSD.n2353 VSSD.n2352 4.51401
R12772 VSSD.n2298 VSSD.n1434 4.51401
R12773 VSSD.n1445 VSSD.n1438 4.51401
R12774 VSSD.n2040 VSSD.n2029 4.51401
R12775 VSSD.n2045 VSSD.n2044 4.51401
R12776 VSSD.n1984 VSSD.n1955 4.51401
R12777 VSSD.n1989 VSSD.n1988 4.51401
R12778 VSSD.n2245 VSSD.n2242 4.51401
R12779 VSSD.n2250 VSSD.n2239 4.51401
R12780 VSSD.n1640 VSSD 4.51401
R12781 VSSD.n1846 VSSD.n1845 4.51401
R12782 VSSD.n1594 VSSD.n1593 4.51401
R12783 VSSD.n1891 VSSD.n1890 4.51401
R12784 VSSD.n1951 VSSD.n1572 4.51401
R12785 VSSD.n1941 VSSD.n1937 4.51401
R12786 VSSD.n1679 VSSD.n1671 4.51401
R12787 VSSD.n1796 VSSD.n1795 4.51401
R12788 VSSD.n233 VSSD.n231 4.51401
R12789 VSSD.n335 VSSD.n334 4.51401
R12790 VSSD.n3515 VSSD.n83 4.51401
R12791 VSSD.n3520 VSSD.n3519 4.51401
R12792 VSSD.n3466 VSSD.n101 4.51401
R12793 VSSD.n3471 VSSD.n3470 4.51401
R12794 VSSD.n3420 VSSD.n127 4.51401
R12795 VSSD.n3424 VSSD.n122 4.51401
R12796 VSSD.n3563 VSSD.n60 4.51401
R12797 VSSD.n3568 VSSD.n3567 4.51401
R12798 VSSD.n148 VSSD.n141 4.51401
R12799 VSSD.n475 VSSD.n474 4.51401
R12800 VSSD.n507 VSSD.n502 4.5005
R12801 VSSD.n3384 VSSD.n3383 4.5005
R12802 VSSD.n511 VSSD.n504 4.5005
R12803 VSSD.n759 VSSD.n529 4.5005
R12804 VSSD.n757 VSSD.n756 4.5005
R12805 VSSD.n765 VSSD.n764 4.5005
R12806 VSSD.n1010 VSSD.n1009 4.5005
R12807 VSSD.n1008 VSSD.n1007 4.5005
R12808 VSSD.n1004 VSSD.n1003 4.5005
R12809 VSSD.n840 VSSD.n839 4.5005
R12810 VSSD.n853 VSSD.n852 4.5005
R12811 VSSD.n854 VSSD.n843 4.5005
R12812 VSSD.n1307 VSSD.n1306 4.5005
R12813 VSSD.n1169 VSSD.n1136 4.5005
R12814 VSSD.n1172 VSSD.n1168 4.5005
R12815 VSSD.n1209 VSSD.n1152 4.5005
R12816 VSSD.n1222 VSSD.n1221 4.5005
R12817 VSSD.n1220 VSSD.n1149 4.5005
R12818 VSSD.n3329 VSSD.n3328 4.5005
R12819 VSSD.n3327 VSSD.n3326 4.5005
R12820 VSSD.n3323 VSSD.n3322 4.5005
R12821 VSSD.n3196 VSSD.n3195 4.5005
R12822 VSSD.n3188 VSSD.n3187 4.5005
R12823 VSSD.n1050 VSSD.n1049 4.5005
R12824 VSSD.n2886 VSSD.n2885 4.5005
R12825 VSSD.n2858 VSSD.n2857 4.5005
R12826 VSSD.n1130 VSSD.n1129 4.5005
R12827 VSSD.n2943 VSSD.n2942 4.5005
R12828 VSSD.n1111 VSSD.n1110 4.5005
R12829 VSSD.n2936 VSSD.n1102 4.5005
R12830 VSSD.n2989 VSSD.n1086 4.5005
R12831 VSSD.n2999 VSSD.n2998 4.5005
R12832 VSSD.n1087 VSSD.n1083 4.5005
R12833 VSSD.n3147 VSSD.n3146 4.5005
R12834 VSSD.n1062 VSSD.n1058 4.5005
R12835 VSSD.n3141 VSSD.n3140 4.5005
R12836 VSSD.n2554 VSSD.n2553 4.5005
R12837 VSSD.n2575 VSSD.n2574 4.5005
R12838 VSSD.n2552 VSSD.n2548 4.5005
R12839 VSSD.n2623 VSSD.n2622 4.5005
R12840 VSSD.n2535 VSSD.n2534 4.5005
R12841 VSSD.n2532 VSSD.n1372 4.5005
R12842 VSSD.n2845 VSSD.n2844 4.5005
R12843 VSSD.n2843 VSSD.n2842 4.5005
R12844 VSSD.n2839 VSSD.n2838 4.5005
R12845 VSSD.n1353 VSSD.n1348 4.5005
R12846 VSSD.n2801 VSSD.n2800 4.5005
R12847 VSSD.n1357 VSSD.n1351 4.5005
R12848 VSSD.n1565 VSSD.n1564 4.5005
R12849 VSSD.n1553 VSSD.n1478 4.5005
R12850 VSSD.n1558 VSSD.n1557 4.5005
R12851 VSSD.n2523 VSSD.n2522 4.5005
R12852 VSSD.n2511 VSSD.n1380 4.5005
R12853 VSSD.n2514 VSSD.n1383 4.5005
R12854 VSSD.n2474 VSSD.n2473 4.5005
R12855 VSSD.n1403 VSSD.n1401 4.5005
R12856 VSSD.n1409 VSSD.n1405 4.5005
R12857 VSSD.n2347 VSSD.n2346 4.5005
R12858 VSSD.n2311 VSSD.n2310 4.5005
R12859 VSSD.n1427 VSSD.n1426 4.5005
R12860 VSSD.n1983 VSSD.n1982 4.5005
R12861 VSSD.n1959 VSSD.n1958 4.5005
R12862 VSSD.n1472 VSSD.n1471 4.5005
R12863 VSSD.n2039 VSSD.n2038 4.5005
R12864 VSSD.n2036 VSSD.n2035 4.5005
R12865 VSSD.n2033 VSSD.n1452 4.5005
R12866 VSSD.n2297 VSSD.n2296 4.5005
R12867 VSSD.n2295 VSSD.n2294 4.5005
R12868 VSSD.n2291 VSSD.n2290 4.5005
R12869 VSSD.n2244 VSSD.n2243 4.5005
R12870 VSSD.n2240 VSSD.n2125 4.5005
R12871 VSSD.n2252 VSSD.n2251 4.5005
R12872 VSSD.n1898 VSSD.n1897 4.5005
R12873 VSSD.n1621 VSSD.n1595 4.5005
R12874 VSSD.n1622 VSSD.n1597 4.5005
R12875 VSSD.n1853 VSSD.n1852 4.5005
R12876 VSSD.n1646 VSSD.n1641 4.5005
R12877 VSSD.n1647 VSSD.n1643 4.5005
R12878 VSSD.n1950 VSSD.n1949 4.5005
R12879 VSSD.n1938 VSSD.n1574 4.5005
R12880 VSSD.n1943 VSSD.n1942 4.5005
R12881 VSSD.n1678 VSSD.n1673 4.5005
R12882 VSSD.n1801 VSSD.n1800 4.5005
R12883 VSSD.n1682 VSSD.n1676 4.5005
R12884 VSSD.n3419 VSSD.n3418 4.5005
R12885 VSSD.n128 VSSD.n121 4.5005
R12886 VSSD.n3426 VSSD.n3425 4.5005
R12887 VSSD.n3465 VSSD.n3464 4.5005
R12888 VSSD.n108 VSSD.n107 4.5005
R12889 VSSD.n105 VSSD.n97 4.5005
R12890 VSSD.n3514 VSSD.n3513 4.5005
R12891 VSSD.n3512 VSSD.n3511 4.5005
R12892 VSSD.n79 VSSD.n78 4.5005
R12893 VSSD.n3562 VSSD.n3561 4.5005
R12894 VSSD.n64 VSSD.n63 4.5005
R12895 VSSD.n56 VSSD.n55 4.5005
R12896 VSSD.n147 VSSD.n143 4.5005
R12897 VSSD.n480 VSSD.n479 4.5005
R12898 VSSD.n152 VSSD.n146 4.5005
R12899 VSSD.n432 VSSD.n431 4.5005
R12900 VSSD.n173 VSSD.n168 4.5005
R12901 VSSD.n174 VSSD.n170 4.5005
R12902 VSSD.n386 VSSD.n385 4.5005
R12903 VSSD.n203 VSSD.n201 4.5005
R12904 VSSD.n207 VSSD.n205 4.5005
R12905 VSSD.n232 VSSD.n227 4.5005
R12906 VSSD.n340 VSSD.n339 4.5005
R12907 VSSD.n236 VSSD.n230 4.5005
R12908 VSSD.n576 VSSD.n570 4.5005
R12909 VSSD.n662 VSSD.n661 4.5005
R12910 VSSD.n580 VSSD.n573 4.5005
R12911 VSSD.n615 VSSD.n614 4.5005
R12912 VSSD.n604 VSSD.n601 4.5005
R12913 VSSD.n605 VSSD.n603 4.5005
R12914 VSSD.n731 VSSD.n730 4.5005
R12915 VSSD.n729 VSSD.n728 4.5005
R12916 VSSD.n725 VSSD.n724 4.5005
R12917 VSSD.n3699 VSSD.n3698 4.5005
R12918 VSSD.n33 VSSD.n32 4.5005
R12919 VSSD.n3706 VSSD.n3705 4.5005
R12920 VSSD.n2461 VSSD.n2460 4.49412
R12921 VSSD.n642 VSSD.n586 4.36875
R12922 VSSD.n589 VSSD.n588 4.36875
R12923 VSSD.n631 VSSD.n590 4.36875
R12924 VSSD.n593 VSSD.n592 4.36875
R12925 VSSD.n620 VSSD.n594 4.36875
R12926 VSSD.n597 VSSD.n596 4.36875
R12927 VSSD.n307 VSSD.n253 4.36875
R12928 VSSD.n294 VSSD.n259 4.36875
R12929 VSSD.n287 VSSD.n260 4.36875
R12930 VSSD.n274 VSSD.n266 4.36875
R12931 VSSD.n1290 VSSD.n1148 4.29369
R12932 VSSD.n896 VSSD.n895 4.28986
R12933 VSSD.n3388 VSSD.n3387 4.28986
R12934 VSSD.n2883 VSSD.n2879 4.28986
R12935 VSSD.n2568 VSSD.n2547 4.28986
R12936 VSSD.n2460 VSSD.n1414 4.28986
R12937 VSSD.n2027 VSSD.n2026 4.28986
R12938 VSSD.n1829 VSSD.n1656 4.28986
R12939 VSSD.n1836 VSSD.n1835 4.28986
R12940 VSSD.n3043 VSSD.n3042 4.2869
R12941 VSSD.n1233 VSSD.n1231 4.22178
R12942 VSSD.n718 VSSD.n717 4.11798
R12943 VSSD.n717 VSSD.n716 4.11798
R12944 VSSD.n688 VSSD.n687 4.11798
R12945 VSSD.n944 VSSD.n943 4.11798
R12946 VSSD.n3364 VSSD.n3363 4.11798
R12947 VSSD.n3288 VSSD.n3238 4.11798
R12948 VSSD.n3285 VSSD.n3238 4.11798
R12949 VSSD.n2919 VSSD.n1117 4.11798
R12950 VSSD.n2922 VSSD.n1117 4.11798
R12951 VSSD.n2775 VSSD.n1369 4.11798
R12952 VSSD.n2772 VSSD.n1369 4.11798
R12953 VSSD.n2753 VSSD.n2703 4.11798
R12954 VSSD.n2750 VSSD.n2703 4.11798
R12955 VSSD.n2439 VSSD.n2392 4.11798
R12956 VSSD.n2436 VSSD.n2392 4.11798
R12957 VSSD.n1751 VSSD.n1750 4.11798
R12958 VSSD.n1750 VSSD.n1749 4.11798
R12959 VSSD.n1926 VSSD.n1925 4.11798
R12960 VSSD.n3436 VSSD.n116 4.11798
R12961 VSSD.n3439 VSSD.n116 4.11798
R12962 VSSD.n3456 VSSD.n109 4.11798
R12963 VSSD.n3459 VSSD.n109 4.11798
R12964 VSSD.n3492 VSSD.n88 4.11798
R12965 VSSD.n3495 VSSD.n88 4.11798
R12966 VSSD.n3524 VSSD.n75 4.11798
R12967 VSSD.n3527 VSSD.n75 4.11798
R12968 VSSD.n3553 VSSD.n65 4.11798
R12969 VSSD.n3556 VSSD.n65 4.11798
R12970 VSSD.n3582 VSSD.n49 4.11798
R12971 VSSD.n3585 VSSD.n49 4.11798
R12972 VSSD.n3643 VSSD.n3597 4.11798
R12973 VSSD.n3640 VSSD.n3597 4.11798
R12974 VSSD.n3623 VSSD.n3604 4.11798
R12975 VSSD.n3620 VSSD.n3604 4.11798
R12976 VSSD.n3751 VSSD.n3750 4.11798
R12977 VSSD.n3752 VSSD.n3751 4.11798
R12978 VSSD.n1415 VSSD.n1414 4.07323
R12979 VSSD.n2026 VSSD.n1451 4.07323
R12980 VSSD.n3264 VSSD.n3247 4.03876
R12981 VSSD.n2729 VSSD.n2712 4.03876
R12982 VSSD.n1728 VSSD.n1711 4.03876
R12983 VSSD.n1835 VSSD.n1834 3.97291
R12984 VSSD.n1217 VSSD.n1214 3.96548
R12985 VSSD.n3259 VSSD.n3258 3.96548
R12986 VSSD.n2724 VSSD.n2723 3.96548
R12987 VSSD.n2412 VSSD.n2411 3.96548
R12988 VSSD.n2411 VSSD.n2401 3.96548
R12989 VSSD.n1723 VSSD.n1722 3.96548
R12990 VSSD.n317 VSSD.n316 3.96548
R12991 VSSD.n3777 VSSD.n3776 3.96548
R12992 VSSD.n3778 VSSD.n3777 3.96548
R12993 VSSD.n3782 VSSD.n3781 3.96548
R12994 VSSD.n3314 VSSD.n1027 3.95596
R12995 VSSD.n893 VSSD.n890 3.90948
R12996 VSSD.n3386 VSSD.n501 3.90948
R12997 VSSD.n3059 VSSD.n3057 3.90948
R12998 VSSD.n3059 VSSD.n3058 3.90948
R12999 VSSD.n2572 VSSD.n2571 3.90948
R13000 VSSD.n1257 VSSD.n1256 3.76521
R13001 VSSD.n2653 VSSD.n2652 3.76521
R13002 VSSD.n2820 VSSD.n1329 3.76521
R13003 VSSD.n3769 VSSD.n3767 3.7575
R13004 VSSD.n3319 VSSD.n3318 3.74518
R13005 VSSD.n582 VSSD.n569 3.7069
R13006 VSSD.n1289 VSSD.n1288 3.7069
R13007 VSSD.n1288 VSSD.n1287 3.7069
R13008 VSSD.n1214 VSSD.n1153 3.7069
R13009 VSSD.n3260 VSSD.n3259 3.7069
R13010 VSSD.n2725 VSSD.n2724 3.7069
R13011 VSSD.n2414 VSSD.n2399 3.7069
R13012 VSSD.n2402 VSSD.n2401 3.7069
R13013 VSSD.n1724 VSSD.n1723 3.7069
R13014 VSSD.n1905 VSSD.n1590 3.7069
R13015 VSSD.n319 VSSD.n245 3.7069
R13016 VSSD.n3776 VSSD.n4 3.7069
R13017 VSSD.n3784 VSSD.n0 3.7069
R13018 VSSD.n654 VSSD.n582 3.68605
R13019 VSSD.n665 VSSD.n664 3.59021
R13020 VSSD.n943 VSSD.n942 3.58092
R13021 VSSD.n3313 VSSD.n1028 3.50735
R13022 VSSD.n1278 VSSD.n1234 3.50735
R13023 VSSD.n2898 VSSD.n2897 3.50735
R13024 VSSD.n1833 VSSD.n1655 3.47385
R13025 VSSD.n2882 VSSD.n2880 3.47284
R13026 VSSD.n3220 VSSD.n3219 3.44377
R13027 VSSD.n3220 VSSD.n1040 3.44377
R13028 VSSD.n3225 VSSD.n1040 3.44377
R13029 VSSD.n3171 VSSD.n3158 3.44377
R13030 VSSD.n3175 VSSD.n3158 3.44377
R13031 VSSD.n3048 VSSD.n3047 3.44377
R13032 VSSD.n1520 VSSD.n1519 3.44377
R13033 VSSD.n1519 VSSD.n1518 3.44377
R13034 VSSD.n435 VSSD.n434 3.44377
R13035 VSSD.n434 VSSD.n165 3.44377
R13036 VSSD.n658 VSSD.n657 3.43925
R13037 VSSD.n578 VSSD.n577 3.43925
R13038 VSSD.n609 VSSD.n608 3.43925
R13039 VSSD.n611 VSSD.n600 3.43925
R13040 VSSD.n426 VSSD.n425 3.43925
R13041 VSSD.n428 VSSD.n167 3.43925
R13042 VSSD.n543 VSSD.n537 3.43925
R13043 VSSD.n733 VSSD.n732 3.43925
R13044 VSSD.n380 VSSD.n379 3.43925
R13045 VSSD.n382 VSSD.n202 3.43925
R13046 VSSD.n3704 VSSD.n3703 3.43925
R13047 VSSD.n3701 VSSD.n3700 3.43925
R13048 VSSD.n741 VSSD.n735 3.43925
R13049 VSSD.n1012 VSSD.n1011 3.43925
R13050 VSSD.n766 VSSD.n532 3.43925
R13051 VSSD.n3339 VSSD.n3338 3.43925
R13052 VSSD.n3380 VSSD.n3379 3.43925
R13053 VSSD.n509 VSSD.n508 3.43925
R13054 VSSD.n960 VSSD.n959 3.43925
R13055 VSSD.n964 VSSD.n963 3.43925
R13056 VSSD.n1020 VSSD.n1014 3.43925
R13057 VSSD.n3331 VSSD.n3330 3.43925
R13058 VSSD.n1226 VSSD.n1225 3.43925
R13059 VSSD.n1211 VSSD.n1210 3.43925
R13060 VSSD.n1173 VSSD.n1132 3.43925
R13061 VSSD.n1309 VSSD.n1308 3.43925
R13062 VSSD.n3201 VSSD.n3200 3.43925
R13063 VSSD.n3198 VSSD.n3197 3.43925
R13064 VSSD.n3003 VSSD.n3002 3.43925
R13065 VSSD.n2991 VSSD.n2990 3.43925
R13066 VSSD.n2948 VSSD.n2947 3.43925
R13067 VSSD.n2945 VSSD.n2944 3.43925
R13068 VSSD.n2891 VSSD.n2890 3.43925
R13069 VSSD.n2888 VSSD.n2887 3.43925
R13070 VSSD.n3139 VSSD.n1053 3.43925
R13071 VSSD.n3149 VSSD.n3148 3.43925
R13072 VSSD.n1320 VSSD.n1313 3.43925
R13073 VSSD.n2847 VSSD.n2846 3.43925
R13074 VSSD.n2628 VSSD.n2627 3.43925
R13075 VSSD.n2625 VSSD.n2624 3.43925
R13076 VSSD.n2579 VSSD.n2578 3.43925
R13077 VSSD.n2556 VSSD.n2555 3.43925
R13078 VSSD.n2797 VSSD.n2796 3.43925
R13079 VSSD.n1355 VSSD.n1354 3.43925
R13080 VSSD.n2468 VSSD.n2467 3.43925
R13081 VSSD.n2470 VSSD.n1402 3.43925
R13082 VSSD.n2515 VSSD.n1374 3.43925
R13083 VSSD.n2525 VSSD.n2524 3.43925
R13084 VSSD.n1556 VSSD.n1474 3.43925
R13085 VSSD.n1567 VSSD.n1566 3.43925
R13086 VSSD.n2352 VSSD.n2351 3.43925
R13087 VSSD.n2349 VSSD.n2348 3.43925
R13088 VSSD.n1438 VSSD.n1431 3.43925
R13089 VSSD.n2299 VSSD.n2298 3.43925
R13090 VSSD.n2044 VSSD.n2043 3.43925
R13091 VSSD.n2041 VSSD.n2040 3.43925
R13092 VSSD.n1988 VSSD.n1987 3.43925
R13093 VSSD.n1985 VSSD.n1984 3.43925
R13094 VSSD.n2250 VSSD.n2249 3.43925
R13095 VSSD.n2246 VSSD.n2245 3.43925
R13096 VSSD.n1847 VSSD.n1846 3.43925
R13097 VSSD.n1849 VSSD.n1640 3.43925
R13098 VSSD.n1892 VSSD.n1891 3.43925
R13099 VSSD.n1894 VSSD.n1594 3.43925
R13100 VSSD.n1941 VSSD.n1570 3.43925
R13101 VSSD.n1952 VSSD.n1951 3.43925
R13102 VSSD.n1797 VSSD.n1796 3.43925
R13103 VSSD.n1680 VSSD.n1679 3.43925
R13104 VSSD.n336 VSSD.n335 3.43925
R13105 VSSD.n234 VSSD.n233 3.43925
R13106 VSSD.n3519 VSSD.n3518 3.43925
R13107 VSSD.n3516 VSSD.n3515 3.43925
R13108 VSSD.n3470 VSSD.n3469 3.43925
R13109 VSSD.n3467 VSSD.n3466 3.43925
R13110 VSSD.n3424 VSSD.n3423 3.43925
R13111 VSSD.n3421 VSSD.n3420 3.43925
R13112 VSSD.n3567 VSSD.n3566 3.43925
R13113 VSSD.n3564 VSSD.n3563 3.43925
R13114 VSSD.n574 VSSD.n572 3.4105
R13115 VSSD.n660 VSSD.n659 3.4105
R13116 VSSD.n613 VSSD.n612 3.4105
R13117 VSSD.n610 VSSD.n602 3.4105
R13118 VSSD.n430 VSSD.n429 3.4105
R13119 VSSD.n427 VSSD.n169 3.4105
R13120 VSSD.n540 VSSD.n538 3.4105
R13121 VSSD.n727 VSSD.n726 3.4105
R13122 VSSD.n384 VSSD.n383 3.4105
R13123 VSSD.n381 VSSD.n204 3.4105
R13124 VSSD.n31 VSSD.n29 3.4105
R13125 VSSD.n26 VSSD.n25 3.4105
R13126 VSSD.n738 VSSD.n736 3.4105
R13127 VSSD.n1006 VSSD.n1005 3.4105
R13128 VSSD.n755 VSSD.n530 3.4105
R13129 VSSD.n754 VSSD.n753 3.4105
R13130 VSSD.n505 VSSD.n503 3.4105
R13131 VSSD.n3382 VSSD.n3381 3.4105
R13132 VSSD.n962 VSSD.n841 3.4105
R13133 VSSD.n961 VSSD.n842 3.4105
R13134 VSSD.n1017 VSSD.n1016 3.4105
R13135 VSSD.n3325 VSSD.n3324 3.4105
R13136 VSSD.n1151 VSSD.n1150 3.4105
R13137 VSSD.n1224 VSSD.n1223 3.4105
R13138 VSSD.n1135 VSSD.n1133 3.4105
R13139 VSSD.n1171 VSSD.n1170 3.4105
R13140 VSSD.n3153 VSSD.n3151 3.4105
R13141 VSSD.n3186 VSSD.n1051 3.4105
R13142 VSSD.n1085 VSSD.n1084 3.4105
R13143 VSSD.n3001 VSSD.n3000 3.4105
R13144 VSSD.n1107 VSSD.n1105 3.4105
R13145 VSSD.n1109 VSSD.n1103 3.4105
R13146 VSSD.n2855 VSSD.n2853 3.4105
R13147 VSSD.n2856 VSSD.n1131 3.4105
R13148 VSSD.n1057 VSSD.n1055 3.4105
R13149 VSSD.n1064 VSSD.n1063 3.4105
R13150 VSSD.n1317 VSSD.n1315 3.4105
R13151 VSSD.n2841 VSSD.n2840 3.4105
R13152 VSSD.n2529 VSSD.n2527 3.4105
R13153 VSSD.n2533 VSSD.n1373 3.4105
R13154 VSSD.n2550 VSSD.n2549 3.4105
R13155 VSSD.n2577 VSSD.n2576 3.4105
R13156 VSSD.n1352 VSSD.n1350 3.4105
R13157 VSSD.n2799 VSSD.n2798 3.4105
R13158 VSSD.n2472 VSSD.n2471 3.4105
R13159 VSSD.n2469 VSSD.n1404 3.4105
R13160 VSSD.n1378 VSSD.n1376 3.4105
R13161 VSSD.n2513 VSSD.n2512 3.4105
R13162 VSSD.n1477 VSSD.n1475 3.4105
R13163 VSSD.n1555 VSSD.n1554 3.4105
R13164 VSSD.n2307 VSSD.n2305 3.4105
R13165 VSSD.n2309 VSSD.n1428 3.4105
R13166 VSSD.n1435 VSSD.n1433 3.4105
R13167 VSSD.n2293 VSSD.n2292 3.4105
R13168 VSSD.n2030 VSSD.n1455 3.4105
R13169 VSSD.n2034 VSSD.n1453 3.4105
R13170 VSSD.n1956 VSSD.n1954 3.4105
R13171 VSSD.n1957 VSSD.n1473 3.4105
R13172 VSSD.n2247 VSSD.n2241 3.4105
R13173 VSSD.n2248 VSSD.n2127 3.4105
R13174 VSSD.n1851 VSSD.n1850 3.4105
R13175 VSSD.n1848 VSSD.n1642 3.4105
R13176 VSSD.n1896 VSSD.n1895 3.4105
R13177 VSSD.n1893 VSSD.n1596 3.4105
R13178 VSSD.n1573 VSSD.n1571 3.4105
R13179 VSSD.n1940 VSSD.n1939 3.4105
R13180 VSSD.n1677 VSSD.n1675 3.4105
R13181 VSSD.n1799 VSSD.n1798 3.4105
R13182 VSSD.n235 VSSD.n229 3.4105
R13183 VSSD.n338 VSSD.n337 3.4105
R13184 VSSD.n84 VSSD.n82 3.4105
R13185 VSSD.n3510 VSSD.n80 3.4105
R13186 VSSD.n102 VSSD.n100 3.4105
R13187 VSSD.n106 VSSD.n98 3.4105
R13188 VSSD.n129 VSSD.n126 3.4105
R13189 VSSD.n124 VSSD.n123 3.4105
R13190 VSSD.n61 VSSD.n59 3.4105
R13191 VSSD.n62 VSSD.n57 3.4105
R13192 VSSD.n476 VSSD.n125 3.4105
R13193 VSSD.n149 VSSD.n125 3.4105
R13194 VSSD.n476 VSSD.n475 3.4105
R13195 VSSD.n149 VSSD.n148 3.4105
R13196 VSSD.n150 VSSD.n145 3.4105
R13197 VSSD.n478 VSSD.n477 3.4105
R13198 VSSD.n3284 VSSD.n3283 3.4019
R13199 VSSD.n2918 VSSD.n2917 3.4019
R13200 VSSD.n2749 VSSD.n2748 3.4019
R13201 VSSD.n2440 VSSD.n2439 3.4019
R13202 VSSD.n1748 VSSD.n1747 3.4019
R13203 VSSD.n1928 VSSD.n1927 3.4019
R13204 VSSD.n3743 VSSD.n3742 3.4019
R13205 VSSD.n1000 VSSD.n999 3.38874
R13206 VSSD.n3208 VSSD.n3207 3.38874
R13207 VSSD.n2954 VSSD.n2953 3.38874
R13208 VSSD.n2812 VSSD.n2811 3.38874
R13209 VSSD.n1823 VSSD.n1661 3.33201
R13210 VSSD.n1362 VSSD.n1361 3.26859
R13211 VSSD.n3219 VSSD.n3218 3.21921
R13212 VSSD.n3171 VSSD.n3170 3.21921
R13213 VSSD.n3049 VSSD.n3048 3.21921
R13214 VSSD.n1520 VSSD.n1516 3.21921
R13215 VSSD.n2520 VSSD.n2519 3.21921
R13216 VSSD.n435 VSSD.n163 3.21921
R13217 VSSD.n172 VSSD.n165 3.21921
R13218 VSSD.n789 VSSD.n779 3.2005
R13219 VSSD.n3310 VSSD.n3309 3.2005
R13220 VSSD.n2266 VSSD.n2115 3.2005
R13221 VSSD.n2220 VSSD.n2219 3.2005
R13222 VSSD.n1820 VSSD.n1819 3.2005
R13223 VSSD.n421 VSSD.n178 3.2005
R13224 VSSD.n675 VSSD.n674 3.13337
R13225 VSSD.n992 VSSD.n747 3.13241
R13226 VSSD.n2874 VSSD.n2859 3.13241
R13227 VSSD.n2827 VSSD.n2826 3.13241
R13228 VSSD.n2793 VSSD.n2792 3.13241
R13229 VSSD.n2328 VSSD.n2327 3.13241
R13230 VSSD.n2172 VSSD.n2163 3.13241
R13231 VSSD.n1610 VSSD.n1609 3.13241
R13232 VSSD.n369 VSSD.n368 3.13241
R13233 VSSD.n495 VSSD.n493 3.05586
R13234 VSSD.n1143 VSSD.n1141 3.05586
R13235 VSSD.n2866 VSSD.n2865 3.05586
R13236 VSSD.n2562 VSSD.n2560 3.05586
R13237 VSSD.n1486 VSSD.n1485 3.05586
R13238 VSSD.n1967 VSSD.n1966 3.05586
R13239 VSSD.n1603 VSSD.n1602 3.05586
R13240 VSSD.n564 VSSD.n563 3.05586
R13241 VSSD.n137 VSSD.n136 3.05586
R13242 VSSD.n891 VSSD.n889 3.04861
R13243 VSSD.n3254 VSSD.n3253 3.04861
R13244 VSSD.n3080 VSSD.n3079 3.04861
R13245 VSSD.n2719 VSSD.n2718 3.04861
R13246 VSSD.n2406 VSSD.n2405 3.04861
R13247 VSSD.n2168 VSSD.n2167 3.04861
R13248 VSSD.n1718 VSSD.n1716 3.04861
R13249 VSSD.n270 VSSD.n269 3.04861
R13250 VSSD.n3791 VSSD.n3790 3.04861
R13251 VSSD.n3386 VSSD.n500 3.04861
R13252 VSSD.n1292 VSSD.n1229 3.04861
R13253 VSSD.n2458 VSSD.n1415 3.04861
R13254 VSSD.n1446 VSSD.n1442 3.04861
R13255 VSSD.n557 VSSD.n555 3.04861
R13256 VSSD.n2899 VSSD.n1126 3.02516
R13257 VSSD.n3769 VSSD.n3768 3.01483
R13258 VSSD.n3724 VSSD.n3723 3.01226
R13259 VSSD.n895 VSSD.n893 2.9514
R13260 VSSD.n3387 VSSD.n3386 2.9514
R13261 VSSD.n2572 VSSD.n2547 2.9514
R13262 VSSD.n674 VSSD.n555 2.90959
R13263 VSSD.n1229 VSSD.n1148 2.90959
R13264 VSSD.n2287 VSSD.n1442 2.90959
R13265 VSSD.n2138 VSSD.n2136 2.89365
R13266 VSSD.n316 VSSD.n247 2.88804
R13267 VSSD.n699 VSSD.n698 2.86484
R13268 VSSD.n2880 VSSD.n1128 2.79199
R13269 VSSD.n2378 VSSD.n2377 2.79199
R13270 VSSD.n3261 VSSD.n3247 2.77203
R13271 VSSD.n2726 VSSD.n2712 2.77203
R13272 VSSD.n1725 VSSD.n1711 2.77203
R13273 VSSD.n422 VSSD.n177 2.76214
R13274 VSSD.n748 VSSD.n747 2.7239
R13275 VSSD.n2826 VSSD.n2825 2.7239
R13276 VSSD.n2792 VSSD.n2791 2.7239
R13277 VSSD.n2329 VSSD.n2328 2.7239
R13278 VSSD.n2379 VSSD.n2378 2.7239
R13279 VSSD.n2164 VSSD.n2163 2.7239
R13280 VSSD.n1609 VSSD.n1608 2.7239
R13281 VSSD.n368 VSSD.n367 2.7239
R13282 VSSD.n3677 VSSD.n39 2.7239
R13283 VSSD.n804 VSSD.n803 2.64398
R13284 VSSD.n814 VSSD.n812 2.63579
R13285 VSSD.n3345 VSSD.n3343 2.63579
R13286 VSSD.n922 VSSD.n876 2.63579
R13287 VSSD.n3205 VSSD.n3204 2.63579
R13288 VSSD.n1179 VSSD.n1178 2.63579
R13289 VSSD.n3127 VSSD.n3126 2.63579
R13290 VSSD.n3125 VSSD.n1072 2.63579
R13291 VSSD.n3091 VSSD.n3073 2.63579
R13292 VSSD.n2652 VSSD.n2651 2.63579
R13293 VSSD.n2592 VSSD.n2543 2.63579
R13294 VSSD.n2595 VSSD.n2594 2.63579
R13295 VSSD.n2357 VSSD.n2355 2.63579
R13296 VSSD.n2501 VSSD.n2499 2.63579
R13297 VSSD.n1561 VSSD.n1560 2.63579
R13298 VSSD.n1549 VSSD.n1501 2.63579
R13299 VSSD.n1994 VSSD.n1993 2.63579
R13300 VSSD.n1991 VSSD.n1470 2.63579
R13301 VSSD.n2190 VSSD.n2156 2.63579
R13302 VSSD.n2186 VSSD.n2185 2.63579
R13303 VSSD.n1882 VSSD.n1880 2.63579
R13304 VSSD.n471 VSSD.n469 2.63579
R13305 VSSD.n472 VSSD.n155 2.63579
R13306 VSSD.n350 VSSD.n349 2.63579
R13307 VSSD.n241 VSSD.n239 2.63579
R13308 VSSD.n3695 VSSD.n35 2.63579
R13309 VSSD.n3710 VSSD.n3708 2.63579
R13310 VSSD.n780 VSSD.n778 2.63064
R13311 VSSD.n787 VSSD.n786 2.63064
R13312 VSSD.n1033 VSSD.n1029 2.63064
R13313 VSSD.n1237 VSSD.n1235 2.63064
R13314 VSSD.n2901 VSSD.n1124 2.63064
R13315 VSSD.n2264 VSSD.n2263 2.63064
R13316 VSSD.n2139 VSSD.n2137 2.63064
R13317 VSSD.n1664 VSSD.n1662 2.63064
R13318 VSSD.n419 VSSD.n418 2.63064
R13319 VSSD.n3761 VSSD.n7 2.5963
R13320 VSSD.n1363 VSSD.n1362 2.58773
R13321 VSSD.n653 VSSD.n583 2.55412
R13322 VSSD.n3320 VSSD.n3319 2.51965
R13323 VSSD.n3301 VSSD.n3300 2.50679
R13324 VSSD.n2766 VSSD.n2765 2.50679
R13325 VSSD.n1765 VSSD.n1695 2.50679
R13326 VSSD.n3041 VSSD.n3040 2.50485
R13327 VSSD.n1275 VSSD.n1274 2.41146
R13328 VSSD.n252 VSSD.n251 2.36572
R13329 VSSD.n642 VSSD.n641 2.33701
R13330 VSSD.n641 VSSD.n640 2.33701
R13331 VSSD.n631 VSSD.n630 2.33701
R13332 VSSD.n630 VSSD.n629 2.33701
R13333 VSSD.n620 VSSD.n619 2.33701
R13334 VSSD.n619 VSSD.n618 2.33701
R13335 VSSD.n299 VSSD.n257 2.33701
R13336 VSSD.n296 VSSD.n257 2.33701
R13337 VSSD.n279 VSSD.n264 2.33701
R13338 VSSD.n276 VSSD.n264 2.33701
R13339 VSSD.n650 VSSD.n649 2.33067
R13340 VSSD.n691 VSSD.n549 2.32777
R13341 VSSD.n953 VSSD.n859 2.32777
R13342 VSSD.n3362 VSSD.n3361 2.32777
R13343 VSSD.n3275 VSSD.n3274 2.32777
R13344 VSSD.n2911 VSSD.n2910 2.32777
R13345 VSSD.n2786 VSSD.n2785 2.32777
R13346 VSSD.n2740 VSSD.n2739 2.32777
R13347 VSSD.n1739 VSSD.n1738 2.32777
R13348 VSSD.n1934 VSSD.n1579 2.32777
R13349 VSSD.n3355 VSSD.n521 2.25932
R13350 VSSD.n1263 VSSD.n1262 2.25932
R13351 VSSD.n3117 VSSD.n3116 2.25932
R13352 VSSD.n2663 VSSD.n2662 2.25932
R13353 VSSD.n2818 VSSD.n2817 2.25932
R13354 VSSD.n2368 VSSD.n2367 2.25932
R13355 VSSD.n1492 VSSD.n1491 2.25932
R13356 VSSD.n1384 VSSD.n1382 2.25932
R13357 VSSD.n1976 VSSD.n1962 2.25932
R13358 VSSD.n1971 VSSD.n1963 2.25932
R13359 VSSD.n2103 VSSD.n2048 2.25932
R13360 VSSD.n2179 VSSD.n2178 2.25932
R13361 VSSD.n489 VSSD.n488 2.25932
R13362 VSSD.n893 VSSD.n892 2.25312
R13363 VSSD.n3114 VSSD.n3059 2.25293
R13364 VSSD.n803 VSSD.n802 2.15702
R13365 VSSD.n3783 VSSD.n3782 2.06919
R13366 VSSD.n3019 VSSD.n1079 2.01789
R13367 VSSD.n313 VSSD.n247 2.01694
R13368 VSSD.n1217 VSSD.n1216 1.98299
R13369 VSSD.n3258 VSSD.n3249 1.98299
R13370 VSSD.n2723 VSSD.n2714 1.98299
R13371 VSSD.n2414 VSSD.n2413 1.98299
R13372 VSSD.n2413 VSSD.n2412 1.98299
R13373 VSSD.n1722 VSSD.n1713 1.98299
R13374 VSSD.n1905 VSSD.n1904 1.98299
R13375 VSSD.n1904 VSSD.n1903 1.98299
R13376 VSSD.n1903 VSSD.n1902 1.98299
R13377 VSSD.n319 VSSD.n318 1.98299
R13378 VSSD.n318 VSSD.n317 1.98299
R13379 VSSD.n3778 VSSD.n2 1.98299
R13380 VSSD.n3781 VSSD.n2 1.98299
R13381 VSSD.n1528 VSSD.n1527 1.97497
R13382 VSSD.n3673 VSSD.n43 1.97497
R13383 VSSD.n2431 VSSD.n2430 1.94656
R13384 VSSD.n585 VSSD.n584 1.91571
R13385 VSSD.n3784 VSSD.n3783 1.8968
R13386 VSSD.n922 VSSD.n921 1.88285
R13387 VSSD.n915 VSSD.n914 1.88285
R13388 VSSD.n1188 VSSD.n1187 1.88285
R13389 VSSD.n2977 VSSD.n2976 1.88285
R13390 VSSD.n2986 VSSD.n2985 1.88285
R13391 VSSD.n3135 VSSD.n3134 1.88285
R13392 VSSD.n3133 VSSD.n3132 1.88285
R13393 VSSD.n3098 VSSD.n3097 1.88285
R13394 VSSD.n2602 VSSD.n2600 1.88285
R13395 VSSD.n2605 VSSD.n2603 1.88285
R13396 VSSD.n2361 VSSD.n2360 1.88285
R13397 VSSD.n1547 VSSD.n1503 1.88285
R13398 VSSD.n1543 VSSD.n1542 1.88285
R13399 VSSD.n2003 VSSD.n2002 1.88285
R13400 VSSD.n1999 VSSD.n1998 1.88285
R13401 VSSD.n2083 VSSD.n2062 1.88285
R13402 VSSD.n2215 VSSD.n2141 1.88285
R13403 VSSD.n2197 VSSD.n2196 1.88285
R13404 VSSD.n2192 VSSD.n2154 1.88285
R13405 VSSD.n2178 VSSD.n2177 1.88285
R13406 VSSD.n1792 VSSD.n1790 1.88285
R13407 VSSD.n1806 VSSD.n1805 1.88285
R13408 VSSD.n1865 VSSD.n1635 1.88285
R13409 VSSD.n461 VSSD.n460 1.88285
R13410 VSSD.n464 VSSD.n463 1.88285
R13411 VSSD.n402 VSSD.n401 1.88285
R13412 VSSD.n399 VSSD.n398 1.88285
R13413 VSSD.n344 VSSD.n224 1.88285
R13414 VSSD.n3692 VSSD.n3691 1.88285
R13415 VSSD.n3713 VSSD.n3712 1.88285
R13416 VSSD.n568 VSSD.n567 1.87783
R13417 VSSD.n2116 VSSD.n2114 1.8416
R13418 VSSD.n1251 VSSD.n1250 1.82498
R13419 VSSD.n3227 VSSD.n3225 1.79699
R13420 VSSD.n3176 VSSD.n3175 1.79699
R13421 VSSD.n3178 VSSD.n3177 1.79699
R13422 VSSD.n3047 VSSD.n3023 1.79699
R13423 VSSD.n1518 VSSD.n1381 1.79699
R13424 VSSD.n718 VSSD.n707 1.79071
R13425 VSSD.n687 VSSD.n549 1.79071
R13426 VSSD.n3363 VSSD.n3362 1.79071
R13427 VSSD.n3296 VSSD.n3295 1.79071
R13428 VSSD.n2761 VSSD.n2760 1.79071
R13429 VSSD.n2072 VSSD.n2071 1.79071
R13430 VSSD.n1700 VSSD.n1697 1.79071
R13431 VSSD.n1915 VSSD.n1914 1.79071
R13432 VSSD.n3755 VSSD.n9 1.79071
R13433 VSSD.n2462 VSSD.n2461 1.77071
R13434 VSSD.n3678 VSSD.n3677 1.77071
R13435 VSSD.n1216 VSSD.n1215 1.72441
R13436 VSSD.n3250 VSSD.n3249 1.72441
R13437 VSSD.n2715 VSSD.n2714 1.72441
R13438 VSSD.n1714 VSSD.n1713 1.72441
R13439 VSSD.n1902 VSSD.n1901 1.72441
R13440 VSSD.n3044 VSSD.n3043 1.72214
R13441 VSSD.n1027 VSSD.n1024 1.70263
R13442 VSSD.n3566 VSSD.n3565 1.69188
R13443 VSSD.n3565 VSSD.n3564 1.69188
R13444 VSSD.n336 VSSD.n58 1.69188
R13445 VSSD.n234 VSSD.n58 1.69188
R13446 VSSD.n1797 VSSD.n1681 1.69188
R13447 VSSD.n1681 VSSD.n1680 1.69188
R13448 VSSD.n2249 VSSD.n1429 1.69188
R13449 VSSD.n2246 VSSD.n1429 1.69188
R13450 VSSD.n2351 VSSD.n2350 1.69188
R13451 VSSD.n2350 VSSD.n2349 1.69188
R13452 VSSD.n2797 VSSD.n1356 1.69188
R13453 VSSD.n1356 VSSD.n1355 1.69188
R13454 VSSD.n3150 VSSD.n1053 1.69188
R13455 VSSD.n3150 VSSD.n3149 1.69188
R13456 VSSD.n3200 VSSD.n3199 1.69188
R13457 VSSD.n3199 VSSD.n3198 1.69188
R13458 VSSD.n960 VSSD.n28 1.69188
R13459 VSSD.n963 VSSD.n28 1.69188
R13460 VSSD.n3703 VSSD.n3702 1.69188
R13461 VSSD.n3702 VSSD.n3701 1.69188
R13462 VSSD.n3518 VSSD.n3517 1.69188
R13463 VSSD.n3517 VSSD.n3516 1.69188
R13464 VSSD.n380 VSSD.n81 1.69188
R13465 VSSD.n382 VSSD.n81 1.69188
R13466 VSSD.n1847 VSSD.n1432 1.69188
R13467 VSSD.n1849 VSSD.n1432 1.69188
R13468 VSSD.n2300 VSSD.n1431 1.69188
R13469 VSSD.n2300 VSSD.n2299 1.69188
R13470 VSSD.n2468 VSSD.n1314 1.69188
R13471 VSSD.n2470 VSSD.n1314 1.69188
R13472 VSSD.n2848 VSSD.n1313 1.69188
R13473 VSSD.n2848 VSSD.n2847 1.69188
R13474 VSSD.n3002 VSSD.n1015 1.69188
R13475 VSSD.n2990 VSSD.n1015 1.69188
R13476 VSSD.n3332 VSSD.n1014 1.69188
R13477 VSSD.n3332 VSSD.n3331 1.69188
R13478 VSSD.n1013 VSSD.n735 1.69188
R13479 VSSD.n1013 VSSD.n1012 1.69188
R13480 VSSD.n734 VSSD.n537 1.69188
R13481 VSSD.n734 VSSD.n733 1.69188
R13482 VSSD.n3469 VSSD.n3468 1.69188
R13483 VSSD.n3468 VSSD.n3467 1.69188
R13484 VSSD.n426 VSSD.n99 1.69188
R13485 VSSD.n428 VSSD.n99 1.69188
R13486 VSSD.n1892 VSSD.n1454 1.69188
R13487 VSSD.n1894 VSSD.n1454 1.69188
R13488 VSSD.n2043 VSSD.n2042 1.69188
R13489 VSSD.n2042 VSSD.n2041 1.69188
R13490 VSSD.n2526 VSSD.n1374 1.69188
R13491 VSSD.n2526 VSSD.n2525 1.69188
R13492 VSSD.n2627 VSSD.n2626 1.69188
R13493 VSSD.n2626 VSSD.n2625 1.69188
R13494 VSSD.n2947 VSSD.n2946 1.69188
R13495 VSSD.n2946 VSSD.n2945 1.69188
R13496 VSSD.n1225 VSSD.n533 1.69188
R13497 VSSD.n1210 VSSD.n533 1.69188
R13498 VSSD.n3337 VSSD.n532 1.69188
R13499 VSSD.n3338 VSSD.n3337 1.69188
R13500 VSSD.n609 VSSD.n531 1.69188
R13501 VSSD.n611 VSSD.n531 1.69188
R13502 VSSD.n3423 VSSD.n3422 1.69188
R13503 VSSD.n3422 VSSD.n3421 1.69188
R13504 VSSD.n1953 VSSD.n1570 1.69188
R13505 VSSD.n1953 VSSD.n1952 1.69188
R13506 VSSD.n1987 VSSD.n1986 1.69188
R13507 VSSD.n1986 VSSD.n1985 1.69188
R13508 VSSD.n1568 VSSD.n1474 1.69188
R13509 VSSD.n1568 VSSD.n1567 1.69188
R13510 VSSD.n2578 VSSD.n1311 1.69188
R13511 VSSD.n2555 VSSD.n1311 1.69188
R13512 VSSD.n2890 VSSD.n2889 1.69188
R13513 VSSD.n2889 VSSD.n2888 1.69188
R13514 VSSD.n1310 VSSD.n1132 1.69188
R13515 VSSD.n1310 VSSD.n1309 1.69188
R13516 VSSD.n3380 VSSD.n510 1.69188
R13517 VSSD.n510 VSSD.n509 1.69188
R13518 VSSD.n658 VSSD.n579 1.69188
R13519 VSSD.n579 VSSD.n578 1.69188
R13520 VSSD.n151 VSSD.n125 1.69188
R13521 VSSD.n2267 VSSD.n2114 1.66625
R13522 VSSD.n3177 VSSD.n3176 1.64728
R13523 VSSD.n3044 VSSD.n3023 1.64728
R13524 VSSD.n2520 VSSD.n1381 1.64728
R13525 VSSD.n2231 VSSD.n2132 1.60837
R13526 VSSD.n928 VSSD.n872 1.50638
R13527 VSSD.n3204 VSSD.n1048 1.50638
R13528 VSSD.n2659 VSSD.n2658 1.50638
R13529 VSSD.n2670 VSSD.n2668 1.50638
R13530 VSSD.n2678 VSSD.n2676 1.50638
R13531 VSSD.n2811 VSSD.n2810 1.50638
R13532 VSSD.n1492 VSSD.n1490 1.50638
R13533 VSSD.n1976 VSSD.n1975 1.50638
R13534 VSSD.n2098 VSSD.n2097 1.50638
R13535 VSSD.n2059 VSSD.n2056 1.50638
R13536 VSSD.n1888 VSSD.n1625 1.50638
R13537 VSSD.n3043 VSSD.n3025 1.49758
R13538 VSSD.n1282 VSSD.n1233 1.43682
R13539 VSSD.n3227 VSSD.n3226 1.42272
R13540 VSSD.n3179 VSSD.n3178 1.42272
R13541 VSSD.n2326 VSSD.n2325 1.3622
R13542 VSSD.n371 VSSD.n370 1.3622
R13543 VSSD.n3679 VSSD.n3678 1.3622
R13544 VSSD.n2024 VSSD.n2023 1.29412
R13545 VSSD.n1655 VSSD.n1654 1.29412
R13546 VSSD.n784 VSSD.n742 1.27173
R13547 VSSD.n3766 VSSD.n3765 1.26739
R13548 VSSD.n2388 VSSD.n2387 1.25365
R13549 VSSD.n3156 VSSD.n3154 1.25267
R13550 VSSD.n3230 VSSD.n3229 1.25267
R13551 VSSD.n1207 VSSD.n1206 1.25033
R13552 VSSD.n982 VSSD.n981 1.18311
R13553 VSSD.n802 VSSD.n801 1.18311
R13554 VSSD.n1298 VSSD.n1297 1.18311
R13555 VSSD.n3015 VSSD.n3014 1.18311
R13556 VSSD.n3401 VSSD.n3400 1.18311
R13557 VSSD.n3411 VSSD.n130 1.18311
R13558 VSSD.n3476 VSSD.n93 1.18311
R13559 VSSD.n3537 VSSD.n70 1.18311
R13560 VSSD.n3610 VSSD.n3609 1.18311
R13561 VSSD.n2875 VSSD.n2874 1.15795
R13562 VSSD.n787 VSSD.n779 1.14023
R13563 VSSD.n3309 VSSD.n1029 1.14023
R13564 VSSD.n1273 VSSD.n1235 1.14023
R13565 VSSD.n2902 VSSD.n2901 1.14023
R13566 VSSD.n2264 VSSD.n2115 1.14023
R13567 VSSD.n2219 VSSD.n2137 1.14023
R13568 VSSD.n1819 VSSD.n1662 1.14023
R13569 VSSD.n3230 VSSD.n1039 1.08588
R13570 VSSD.n3180 VSSD.n3154 1.08588
R13571 VSSD.n3040 VSSD.n3026 1.08588
R13572 VSSD.n439 VSSD.n438 1.08588
R13573 VSSD.n177 VSSD.n176 1.00931
R13574 VSSD.n3165 VSSD.n3164 0.972393
R13575 VSSD.n1414 VSSD.n1413 0.952566
R13576 VSSD.n2026 VSSD.n2025 0.952566
R13577 VSSD.n3009 VSSD.n3008 0.951336
R13578 VSSD.n902 VSSD.n883 0.931411
R13579 VSSD.n1649 VSSD.n1639 0.931411
R13580 VSSD.n1451 VSSD.n1450 0.899674
R13581 VSSD.n790 VSSD.n778 0.877212
R13582 VSSD.n419 VSSD.n180 0.877212
R13583 VSSD.n790 VSSD.n789 0.833377
R13584 VSSD.n1275 VSSD.n1234 0.833377
R13585 VSSD.n2899 VSSD.n2898 0.833377
R13586 VSSD.n2267 VSSD.n2266 0.833377
R13587 VSSD.n2220 VSSD.n2138 0.833377
R13588 VSSD.n1820 VSSD.n1663 0.833377
R13589 VSSD.n422 VSSD.n421 0.833377
R13590 VSSD.n649 VSSD.n584 0.830425
R13591 VSSD.n1274 VSSD.n1273 0.789541
R13592 VSSD.n850 VSSD.n849 0.753441
R13593 VSSD.n976 VSSD.n835 0.753441
R13594 VSSD.n3193 VSSD.n3192 0.753441
R13595 VSSD.n1268 VSSD.n1239 0.753441
R13596 VSSD.n2932 VSSD.n1114 0.753441
R13597 VSSD.n2940 VSSD.n2939 0.753441
R13598 VSSD.n2961 VSSD.n2960 0.753441
R13599 VSSD.n2813 VSSD.n1340 0.753441
R13600 VSSD.n2476 VSSD.n1400 0.753441
R13601 VSSD.n2491 VSSD.n1391 0.753441
R13602 VSSD.n1531 VSSD.n1530 0.753441
R13603 VSSD.n2016 VSSD.n2015 0.753441
R13604 VSSD.n2258 VSSD.n2121 0.753441
R13605 VSSD.n2207 VSSD.n2145 0.753441
R13606 VSSD.n1784 VSSD.n1783 0.753441
R13607 VSSD.n1812 VSSD.n1669 0.753441
R13608 VSSD.n3768 VSSD.n5 0.743162
R13609 VSSD.n1927 VSSD.n1926 0.716584
R13610 VSSD.n895 VSSD.n894 0.69032
R13611 VSSD.n2223 VSSD.n2136 0.614199
R13612 VSSD.n650 VSSD.n583 0.606984
R13613 VSSD.n579 VSSD.n575 0.581224
R13614 VSSD.n2547 VSSD.n2546 0.558563
R13615 VSSD.n1569 VSSD.n1430 0.551088
R13616 VSSD.n2852 VSSD.n2851 0.551088
R13617 VSSD.n3335 VSSD.n534 0.551088
R13618 VSSD.n700 VSSD.n699 0.537563
R13619 VSSD.n711 VSSD.n44 0.537563
R13620 VSSD.n679 VSSD.n678 0.537563
R13621 VSSD.n696 VSSD.n546 0.537563
R13622 VSSD.n956 VSSD.n955 0.537563
R13623 VSSD.n942 VSSD.n941 0.537563
R13624 VSSD.n940 VSSD.n864 0.537563
R13625 VSSD.n3374 VSSD.n514 0.537563
R13626 VSSD.n3356 VSSD.n520 0.537563
R13627 VSSD.n3279 VSSD.n3241 0.537563
R13628 VSSD.n3278 VSSD.n3242 0.537563
R13629 VSSD.n3265 VSSD.n3264 0.537563
R13630 VSSD.n2906 VSSD.n1123 0.537563
R13631 VSSD.n2927 VSSD.n1115 0.537563
R13632 VSSD.n2789 VSSD.n1364 0.537563
R13633 VSSD.n2776 VSSD.n2775 0.537563
R13634 VSSD.n2767 VSSD.n2695 0.537563
R13635 VSSD.n2744 VSSD.n2706 0.537563
R13636 VSSD.n2743 VSSD.n2707 0.537563
R13637 VSSD.n2730 VSSD.n2729 0.537563
R13638 VSSD.n2387 VSSD.n2385 0.537563
R13639 VSSD.n2431 VSSD.n2394 0.537563
R13640 VSSD.n2428 VSSD.n2395 0.537563
R13641 VSSD.n2419 VSSD.n2418 0.537563
R13642 VSSD.n2068 VSSD.n2066 0.537563
R13643 VSSD.n2282 VSSD.n2281 0.537563
R13644 VSSD.n1742 VSSD.n1706 0.537563
R13645 VSSD.n1729 VSSD.n1728 0.537563
R13646 VSSD.n1743 VSSD.n1705 0.537563
R13647 VSSD.n1947 VSSD.n1946 0.537563
R13648 VSSD.n1920 VSSD.n1584 0.537563
R13649 VSSD.n1919 VSSD.n1585 0.537563
R13650 VSSD.n1618 VSSD.n1592 0.537563
R13651 VSSD.n1624 VSSD.n1619 0.537563
R13652 VSSD.n3416 VSSD.n120 0.537563
R13653 VSSD.n3444 VSSD.n114 0.537563
R13654 VSSD.n3445 VSSD.n113 0.537563
R13655 VSSD.n3461 VSSD.n95 0.537563
R13656 VSSD.n3481 VSSD.n92 0.537563
R13657 VSSD.n3500 VSSD.n86 0.537563
R13658 VSSD.n3502 VSSD.n3501 0.537563
R13659 VSSD.n3529 VSSD.n72 0.537563
R13660 VSSD.n3542 VSSD.n69 0.537563
R13661 VSSD.n3570 VSSD.n54 0.537563
R13662 VSSD.n3571 VSSD.n53 0.537563
R13663 VSSD.n3587 VSSD.n47 0.537563
R13664 VSSD.n3594 VSSD.n3592 0.537563
R13665 VSSD.n3635 VSSD.n3599 0.537563
R13666 VSSD.n3634 VSSD.n3600 0.537563
R13667 VSSD.n3615 VSSD.n3606 0.537563
R13668 VSSD.n332 VSSD.n331 0.537563
R13669 VSSD.n324 VSSD.n323 0.537563
R13670 VSSD.n3738 VSSD.n3737 0.537563
R13671 VSSD.n780 VSSD.n777 0.526527
R13672 VSSD.n3314 VSSD.n3313 0.526527
R13673 VSSD.n1031 VSSD.n1028 0.526527
R13674 VSSD.n2116 VSSD.n2111 0.526527
R13675 VSSD.n2224 VSSD.n2223 0.526527
R13676 VSSD.n1824 VSSD.n1823 0.526527
R13677 VSSD.n863 VSSD.n861 0.448052
R13678 VSSD.n3268 VSSD.n3267 0.448052
R13679 VSSD.n2779 VSSD.n2778 0.448052
R13680 VSSD.n2733 VSSD.n2732 0.448052
R13681 VSSD.n2423 VSSD.n2397 0.448052
R13682 VSSD.n1732 VSSD.n1731 0.448052
R13683 VSSD.n244 VSSD.n242 0.448052
R13684 VSSD.n3760 VSSD.n3757 0.448052
R13685 VSSD.n830 VSSD.n828 0.417891
R13686 VSSD.n981 VSSD.n980 0.417891
R13687 VSSD.n806 VSSD.n805 0.417891
R13688 VSSD.n801 VSSD.n800 0.417891
R13689 VSSD.n1144 VSSD.n1139 0.417891
R13690 VSSD.n1299 VSSD.n1298 0.417891
R13691 VSSD.n3009 VSSD.n1080 0.417891
R13692 VSSD.n3404 VSSD.n3403 0.417891
R13693 VSSD.n3410 VSSD.n3409 0.417891
R13694 VSSD.n3415 VSSD.n130 0.417891
R13695 VSSD.n3475 VSSD.n3474 0.417891
R13696 VSSD.n3480 VSSD.n93 0.417891
R13697 VSSD.n3536 VSSD.n3535 0.417891
R13698 VSSD.n3541 VSSD.n70 0.417891
R13699 VSSD.n3614 VSSD.n3607 0.417891
R13700 VSSD.n3702 VSSD.n27 0.410635
R13701 VSSD.n734 VSSD.n536 0.410635
R13702 VSSD.n575 VSSD.n531 0.410635
R13703 VSSD.n902 VSSD.n901 0.409011
R13704 VSSD.n995 VSSD.n994 0.409011
R13705 VSSD.n989 VSSD.n748 0.409011
R13706 VSSD.n776 VSSD.n774 0.409011
R13707 VSSD.n496 VSSD.n491 0.409011
R13708 VSSD.n3165 VSSD.n3160 0.409011
R13709 VSSD.n1250 VSSD.n1022 0.409011
R13710 VSSD.n2870 VSSD.n2869 0.409011
R13711 VSSD.n3020 VSSD.n1077 0.409011
R13712 VSSD.n2831 VSSD.n1327 0.409011
R13713 VSSD.n2825 VSSD.n2824 0.409011
R13714 VSSD.n2563 VSSD.n2558 0.409011
R13715 VSSD.n1361 VSSD.n1347 0.409011
R13716 VSSD.n2791 VSSD.n2790 0.409011
R13717 VSSD.n2322 VSSD.n2317 0.409011
R13718 VSSD.n2330 VSSD.n2329 0.409011
R13719 VSSD.n2372 VSSD.n1419 0.409011
R13720 VSSD.n2380 VSSD.n2379 0.409011
R13721 VSSD.n2464 VSSD.n2463 0.409011
R13722 VSSD.n2022 VSSD.n2021 0.409011
R13723 VSSD.n2276 VSSD.n2109 0.409011
R13724 VSSD.n2231 VSSD.n2230 0.409011
R13725 VSSD.n2176 VSSD.n2161 0.409011
R13726 VSSD.n2173 VSSD.n2162 0.409011
R13727 VSSD.n2169 VSSD.n2164 0.409011
R13728 VSSD.n1777 VSSD.n1776 0.409011
R13729 VSSD.n1770 VSSD.n1692 0.409011
R13730 VSSD.n1766 VSSD.n1694 0.409011
R13731 VSSD.n1660 VSSD.n1658 0.409011
R13732 VSSD.n1650 VSSD.n1649 0.409011
R13733 VSSD.n1615 VSSD.n1599 0.409011
R13734 VSSD.n1612 VSSD.n1611 0.409011
R13735 VSSD.n374 VSSD.n212 0.409011
R13736 VSSD.n367 VSSD.n366 0.409011
R13737 VSSD.n3682 VSSD.n39 0.409011
R13738 VSSD.n1281 VSSD.n1278 0.395021
R13739 VSSD.n654 VSSD.n653 0.383542
R13740 VSSD.n2304 VSSD.n2303 0.3805
R13741 VSSD.n1312 VSSD.n1054 0.3805
R13742 VSSD.n2850 VSSD.n2849 0.3805
R13743 VSSD.n2302 VSSD.n2301 0.3805
R13744 VSSD.n3334 VSSD.n3333 0.3805
R13745 VSSD.n1052 VSSD.n535 0.3805
R13746 VSSD.n3336 VSSD.n3335 0.3805
R13747 VSSD.n2851 VSSD.n1104 0.3805
R13748 VSSD.n1430 VSSD.n1375 0.3805
R13749 VSSD.n2080 VSSD.n2062 0.376971
R13750 VSSD.n680 VSSD.n551 0.358542
R13751 VSSD.n935 VSSD.n934 0.358542
R13752 VSSD.n3370 VSSD.n3369 0.358542
R13753 VSSD.n3235 VSSD.n3233 0.358542
R13754 VSSD.n2700 VSSD.n2698 0.358542
R13755 VSSD.n1763 VSSD.n1762 0.358542
R13756 VSSD.n3016 VSSD.n3015 0.348326
R13757 VSSD.n2303 VSSD 0.340994
R13758 VSSD.n1312 VSSD 0.340994
R13759 VSSD.n535 VSSD 0.340994
R13760 VSSD.n27 VSSD 0.340994
R13761 VSSD.n2377 VSSD.n2376 0.340926
R13762 VSSD.n1775 VSSD.n1774 0.340926
R13763 VSSD.n3675 VSSD.n3674 0.340926
R13764 VSSD.n3310 VSSD.n1031 0.307349
R13765 VSSD.n645 VSSD.n586 0.305262
R13766 VSSD.n635 VSSD.n589 0.305262
R13767 VSSD.n634 VSSD.n590 0.305262
R13768 VSSD.n624 VSSD.n593 0.305262
R13769 VSSD.n623 VSSD.n594 0.305262
R13770 VSSD.n596 VSSD.n556 0.305262
R13771 VSSD.n310 VSSD.n253 0.305262
R13772 VSSD.n291 VSSD.n259 0.305262
R13773 VSSD.n290 VSSD.n260 0.305262
R13774 VSSD.n271 VSSD.n266 0.305262
R13775 VSSD.n1607 VSSD.n1575 0.27284
R13776 VSSD.n3306 VSSD.n1033 0.263514
R13777 VSSD.n1270 VSSD.n1237 0.263514
R13778 VSSD.n2896 VSSD.n2895 0.263514
R13779 VSSD.n2897 VSSD.n2896 0.263514
R13780 VSSD.n2905 VSSD.n1124 0.263514
R13781 VSSD.n2263 VSSD.n2262 0.263514
R13782 VSSD.n2216 VSSD.n2139 0.263514
R13783 VSSD.n1816 VSSD.n1664 0.263514
R13784 VSSD.n180 VSSD.n178 0.263514
R13785 VSSD.n418 VSSD.n417 0.263514
R13786 VSSD.n3767 VSSD.n3766 0.262616
R13787 VSSD.n3772 VSSD.n5 0.262616
R13788 VSSD.n664 VSSD.n569 0.259086
R13789 VSSD.n1290 VSSD.n1289 0.259086
R13790 VSSD.n1287 VSSD.n1286 0.259086
R13791 VSSD.n1207 VSSD.n1153 0.259086
R13792 VSSD.n1215 VSSD.n1147 0.259086
R13793 VSSD.n3261 VSSD.n3260 0.259086
R13794 VSSD.n3255 VSSD.n3250 0.259086
R13795 VSSD.n2726 VSSD.n2725 0.259086
R13796 VSSD.n2720 VSSD.n2715 0.259086
R13797 VSSD.n2417 VSSD.n2399 0.259086
R13798 VSSD.n2407 VSSD.n2402 0.259086
R13799 VSSD.n1725 VSSD.n1724 0.259086
R13800 VSSD.n1719 VSSD.n1714 0.259086
R13801 VSSD.n1908 VSSD.n1590 0.259086
R13802 VSSD.n1901 VSSD.n1900 0.259086
R13803 VSSD.n322 VSSD.n245 0.259086
R13804 VSSD.n3773 VSSD.n4 0.259086
R13805 VSSD.n3787 VSSD.n0 0.259086
R13806 VSSD.n2459 VSSD.n2458 0.239726
R13807 VSSD.n892 VSSD 0.238178
R13808 VSSD VSSD.n3114 0.237784
R13809 VSSD.n3218 VSSD.n3217 0.225061
R13810 VSSD.n3226 VSSD.n1039 0.225061
R13811 VSSD.n3170 VSSD.n3169 0.225061
R13812 VSSD.n3180 VSSD.n3179 0.225061
R13813 VSSD.n3050 VSSD.n3049 0.225061
R13814 VSSD.n3026 VSSD.n3025 0.225061
R13815 VSSD.n1523 VSSD.n1516 0.225061
R13816 VSSD.n2519 VSSD.n2518 0.225061
R13817 VSSD.n438 VSSD.n163 0.225061
R13818 VSSD.n176 VSSD.n172 0.225061
R13819 VSSD.n786 VSSD.n785 0.219678
R13820 VSSD.n269 VSSD 0.217246
R13821 VSSD.n995 VSSD.n746 0.207909
R13822 VSSD.n1527 VSSD.n1514 0.204755
R13823 VSSD.n1515 VSSD.n1514 0.204755
R13824 VSSD.n3114 VSSD 0.200023
R13825 VSSD.n892 VSSD 0.199635
R13826 VSSD.n646 VSSD.n585 0.192021
R13827 VSSD.n315 VSSD.n314 0.180304
R13828 VSSD.n3253 VSSD 0.17983
R13829 VSSD.n3079 VSSD 0.17983
R13830 VSSD.n2718 VSSD 0.17983
R13831 VSSD.n2167 VSSD 0.17983
R13832 VSSD.n500 VSSD 0.17983
R13833 VSSD VSSD.n1292 0.17983
R13834 VSSD.n1446 VSSD 0.17983
R13835 VSSD VSSD.n557 0.17983
R13836 VSSD.n715 VSSD.n710 0.179521
R13837 VSSD.n936 VSSD.n935 0.179521
R13838 VSSD.n3300 VSSD.n3233 0.179521
R13839 VSSD.n2765 VSSD.n2698 0.179521
R13840 VSSD.n2069 VSSD.n1440 0.179521
R13841 VSSD.n2283 VSSD.n1444 0.179521
R13842 VSSD.n1763 VSSD.n1695 0.179521
R13843 VSSD.n1589 VSSD.n1587 0.179521
R13844 VSSD VSSD.n891 0.179485
R13845 VSSD.n2405 VSSD 0.179485
R13846 VSSD.n1716 VSSD 0.179485
R13847 VSSD VSSD.n3791 0.179485
R13848 VSSD.n2902 VSSD.n1126 0.175842
R13849 VSSD.n1663 VSSD.n1661 0.175842
R13850 VSSD.n493 VSSD 0.172576
R13851 VSSD.n1141 VSSD 0.172576
R13852 VSSD VSSD.n2866 0.172576
R13853 VSSD.n2560 VSSD 0.172576
R13854 VSSD VSSD.n1486 0.172576
R13855 VSSD VSSD.n1967 0.172576
R13856 VSSD VSSD.n1603 0.172576
R13857 VSSD VSSD.n564 0.172576
R13858 VSSD VSSD.n137 0.172233
R13859 VSSD.n2302 VSSD.n1430 0.171088
R13860 VSSD.n2303 VSSD.n2302 0.171088
R13861 VSSD.n2851 VSSD.n2850 0.171088
R13862 VSSD.n2850 VSSD.n1312 0.171088
R13863 VSSD.n3335 VSSD.n3334 0.171088
R13864 VSSD.n3334 VSSD.n535 0.171088
R13865 VSSD.n575 VSSD.n536 0.171088
R13866 VSSD.n536 VSSD.n27 0.171088
R13867 VSSD.n3702 VSSD.n28 0.1509
R13868 VSSD.n3199 VSSD.n3150 0.1509
R13869 VSSD.n2350 VSSD.n1356 0.1509
R13870 VSSD.n1681 VSSD.n1429 0.1509
R13871 VSSD.n1681 VSSD.n58 0.1509
R13872 VSSD.n3565 VSSD.n58 0.1509
R13873 VSSD.n1013 VSSD.n734 0.1509
R13874 VSSD.n3332 VSSD.n1015 0.1509
R13875 VSSD.n2848 VSSD.n1314 0.1509
R13876 VSSD.n2300 VSSD.n1432 0.1509
R13877 VSSD.n1432 VSSD.n81 0.1509
R13878 VSSD.n3517 VSSD.n81 0.1509
R13879 VSSD.n3337 VSSD.n531 0.1509
R13880 VSSD.n2946 VSSD.n533 0.1509
R13881 VSSD.n2626 VSSD.n2526 0.1509
R13882 VSSD.n2042 VSSD.n1454 0.1509
R13883 VSSD.n1454 VSSD.n99 0.1509
R13884 VSSD.n3468 VSSD.n99 0.1509
R13885 VSSD.n579 VSSD.n510 0.1509
R13886 VSSD.n2889 VSSD.n1310 0.1509
R13887 VSSD.n1568 VSSD.n1311 0.1509
R13888 VSSD.n1986 VSSD.n1953 0.1509
R13889 VSSD.n1953 VSSD.n125 0.1509
R13890 VSSD.n3422 VSSD.n125 0.1509
R13891 VSSD.n891 VSSD 0.14207
R13892 VSSD.n2405 VSSD 0.14207
R13893 VSSD.n1716 VSSD 0.14207
R13894 VSSD.n269 VSSD 0.14207
R13895 VSSD.n3791 VSSD 0.14207
R13896 VSSD.n1292 VSSD 0.141725
R13897 VSSD.n3253 VSSD 0.141725
R13898 VSSD.n3079 VSSD 0.141725
R13899 VSSD.n2718 VSSD 0.141725
R13900 VSSD.n2458 VSSD 0.141725
R13901 VSSD VSSD.n1446 0.141725
R13902 VSSD.n2167 VSSD 0.141725
R13903 VSSD.n557 VSSD 0.141725
R13904 VSSD.n899 VSSD.n886 0.13667
R13905 VSSD.n1843 VSSD.n1842 0.13667
R13906 VSSD.n1608 VSSD.n1607 0.13667
R13907 VSSD.n1282 VSSD.n1281 0.132007
R13908 VSSD.n506 VSSD.n500 0.122194
R13909 VSSD.n2570 VSSD 0.120408
R13910 VSSD VSSD.n667 0.120408
R13911 VSSD VSSD.n553 0.120408
R13912 VSSD.n3373 VSSD.n3372 0.120292
R13913 VSSD.n3372 VSSD.n515 0.120292
R13914 VSSD.n3367 VSSD.n515 0.120292
R13915 VSSD.n3367 VSSD.n3366 0.120292
R13916 VSSD.n3366 VSSD.n3365 0.120292
R13917 VSSD.n3365 VSSD.n517 0.120292
R13918 VSSD.n3359 VSSD.n517 0.120292
R13919 VSSD.n3359 VSSD.n3358 0.120292
R13920 VSSD.n3358 VSSD.n3357 0.120292
R13921 VSSD.n3354 VSSD.n3353 0.120292
R13922 VSSD.n3353 VSSD.n522 0.120292
R13923 VSSD.n3349 VSSD.n522 0.120292
R13924 VSSD.n3349 VSSD.n3348 0.120292
R13925 VSSD.n3348 VSSD.n3347 0.120292
R13926 VSSD.n3347 VSSD.n526 0.120292
R13927 VSSD.n3341 VSSD.n526 0.120292
R13928 VSSD.n823 VSSD.n822 0.120292
R13929 VSSD.n822 VSSD.n768 0.120292
R13930 VSSD.n818 VSSD.n768 0.120292
R13931 VSSD.n818 VSSD.n817 0.120292
R13932 VSSD.n817 VSSD.n816 0.120292
R13933 VSSD.n816 VSSD.n770 0.120292
R13934 VSSD.n809 VSSD.n770 0.120292
R13935 VSSD.n809 VSSD.n808 0.120292
R13936 VSSD.n807 VSSD.n772 0.120292
R13937 VSSD.n799 VSSD.n772 0.120292
R13938 VSSD.n798 VSSD.n797 0.120292
R13939 VSSD.n797 VSSD.n775 0.120292
R13940 VSSD.n793 VSSD.n775 0.120292
R13941 VSSD.n793 VSSD.n792 0.120292
R13942 VSSD.n792 VSSD.n791 0.120292
R13943 VSSD.n998 VSSD.n997 0.120292
R13944 VSSD.n996 VSSD.n745 0.120292
R13945 VSSD.n991 VSSD.n745 0.120292
R13946 VSSD.n991 VSSD.n990 0.120292
R13947 VSSD.n985 VSSD.n984 0.120292
R13948 VSSD.n984 VSSD.n829 0.120292
R13949 VSSD.n977 VSSD.n833 0.120292
R13950 VSSD.n973 VSSD.n833 0.120292
R13951 VSSD.n973 VSSD.n972 0.120292
R13952 VSSD.n972 VSSD.n971 0.120292
R13953 VSSD.n971 VSSD.n837 0.120292
R13954 VSSD.n967 VSSD.n837 0.120292
R13955 VSSD.n967 VSSD.n966 0.120292
R13956 VSSD.n957 VSSD.n845 0.120292
R13957 VSSD.n952 VSSD.n845 0.120292
R13958 VSSD.n952 VSSD.n951 0.120292
R13959 VSSD.n951 VSSD.n860 0.120292
R13960 VSSD.n947 VSSD.n860 0.120292
R13961 VSSD.n947 VSSD.n946 0.120292
R13962 VSSD.n946 VSSD.n945 0.120292
R13963 VSSD.n945 VSSD.n862 0.120292
R13964 VSSD.n939 VSSD.n938 0.120292
R13965 VSSD.n938 VSSD.n865 0.120292
R13966 VSSD.n930 VSSD.n868 0.120292
R13967 VSSD.n930 VSSD.n929 0.120292
R13968 VSSD.n929 VSSD.n871 0.120292
R13969 VSSD.n925 VSSD.n871 0.120292
R13970 VSSD.n925 VSSD.n924 0.120292
R13971 VSSD.n924 VSSD.n923 0.120292
R13972 VSSD.n923 VSSD.n874 0.120292
R13973 VSSD.n918 VSSD.n874 0.120292
R13974 VSSD.n918 VSSD.n917 0.120292
R13975 VSSD.n917 VSSD.n916 0.120292
R13976 VSSD.n916 VSSD.n879 0.120292
R13977 VSSD.n911 VSSD.n879 0.120292
R13978 VSSD.n911 VSSD.n910 0.120292
R13979 VSSD.n910 VSSD.n909 0.120292
R13980 VSSD.n909 VSSD.n882 0.120292
R13981 VSSD.n904 VSSD.n882 0.120292
R13982 VSSD.n903 VSSD.n884 0.120292
R13983 VSSD.n898 VSSD.n884 0.120292
R13984 VSSD.n898 VSSD.n897 0.120292
R13985 VSSD.n1302 VSSD.n1301 0.120292
R13986 VSSD.n1175 VSSD.n1164 0.120292
R13987 VSSD.n1180 VSSD.n1164 0.120292
R13988 VSSD.n1181 VSSD.n1180 0.120292
R13989 VSSD.n1182 VSSD.n1181 0.120292
R13990 VSSD.n1182 VSSD.n1162 0.120292
R13991 VSSD.n1189 VSSD.n1162 0.120292
R13992 VSSD.n1190 VSSD.n1189 0.120292
R13993 VSSD.n1191 VSSD.n1190 0.120292
R13994 VSSD.n1191 VSSD.n1160 0.120292
R13995 VSSD.n1195 VSSD.n1160 0.120292
R13996 VSSD.n1196 VSSD.n1195 0.120292
R13997 VSSD.n1197 VSSD.n1196 0.120292
R13998 VSSD.n1197 VSSD.n1158 0.120292
R13999 VSSD.n1201 VSSD.n1158 0.120292
R14000 VSSD.n1202 VSSD.n1201 0.120292
R14001 VSSD.n1203 VSSD.n1202 0.120292
R14002 VSSD.n1291 VSSD.n1230 0.120292
R14003 VSSD.n1285 VSSD.n1230 0.120292
R14004 VSSD.n1283 VSSD.n1232 0.120292
R14005 VSSD.n1272 VSSD.n1232 0.120292
R14006 VSSD.n1272 VSSD.n1271 0.120292
R14007 VSSD.n1266 VSSD.n1240 0.120292
R14008 VSSD.n1260 VSSD.n1240 0.120292
R14009 VSSD.n1260 VSSD.n1259 0.120292
R14010 VSSD.n1259 VSSD.n1245 0.120292
R14011 VSSD.n1253 VSSD.n1245 0.120292
R14012 VSSD.n3317 VSSD.n3316 0.120292
R14013 VSSD.n3316 VSSD.n3315 0.120292
R14014 VSSD.n3315 VSSD.n1025 0.120292
R14015 VSSD.n3308 VSSD.n1025 0.120292
R14016 VSSD.n3308 VSSD.n3307 0.120292
R14017 VSSD.n3162 VSSD.n3161 0.120292
R14018 VSSD.n3172 VSSD.n3159 0.120292
R14019 VSSD.n3173 VSSD.n3172 0.120292
R14020 VSSD.n3174 VSSD.n3173 0.120292
R14021 VSSD.n3174 VSSD.n3155 0.120292
R14022 VSSD.n3181 VSSD.n3155 0.120292
R14023 VSSD.n3209 VSSD.n1045 0.120292
R14024 VSSD.n3210 VSSD.n3209 0.120292
R14025 VSSD.n3211 VSSD.n3210 0.120292
R14026 VSSD.n3216 VSSD.n1041 0.120292
R14027 VSSD.n3221 VSSD.n1041 0.120292
R14028 VSSD.n3222 VSSD.n3221 0.120292
R14029 VSSD.n3224 VSSD.n3222 0.120292
R14030 VSSD.n3224 VSSD.n3223 0.120292
R14031 VSSD.n3299 VSSD.n3298 0.120292
R14032 VSSD.n3298 VSSD.n3234 0.120292
R14033 VSSD.n3293 VSSD.n3234 0.120292
R14034 VSSD.n3293 VSSD.n3292 0.120292
R14035 VSSD.n3292 VSSD.n3291 0.120292
R14036 VSSD.n3291 VSSD.n3237 0.120292
R14037 VSSD.n3287 VSSD.n3237 0.120292
R14038 VSSD.n3287 VSSD.n3286 0.120292
R14039 VSSD.n3286 VSSD.n3239 0.120292
R14040 VSSD.n3281 VSSD.n3239 0.120292
R14041 VSSD.n3281 VSSD.n3280 0.120292
R14042 VSSD.n3277 VSSD.n3276 0.120292
R14043 VSSD.n3276 VSSD.n3243 0.120292
R14044 VSSD.n3271 VSSD.n3243 0.120292
R14045 VSSD.n3271 VSSD.n3270 0.120292
R14046 VSSD.n3270 VSSD.n3269 0.120292
R14047 VSSD.n3269 VSSD.n3246 0.120292
R14048 VSSD.n3263 VSSD.n3246 0.120292
R14049 VSSD.n3262 VSSD.n3248 0.120292
R14050 VSSD.n3257 VSSD.n3248 0.120292
R14051 VSSD.n3257 VSSD.n3256 0.120292
R14052 VSSD.n2876 VSSD.n2860 0.120292
R14053 VSSD.n2894 VSSD.n1125 0.120292
R14054 VSSD.n2903 VSSD.n1125 0.120292
R14055 VSSD.n2904 VSSD.n2903 0.120292
R14056 VSSD.n2908 VSSD.n2907 0.120292
R14057 VSSD.n2908 VSSD.n1121 0.120292
R14058 VSSD.n2913 VSSD.n1121 0.120292
R14059 VSSD.n2914 VSSD.n2913 0.120292
R14060 VSSD.n2915 VSSD.n2914 0.120292
R14061 VSSD.n2915 VSSD.n1118 0.120292
R14062 VSSD.n2920 VSSD.n1118 0.120292
R14063 VSSD.n2921 VSSD.n2920 0.120292
R14064 VSSD.n2921 VSSD.n1116 0.120292
R14065 VSSD.n2925 VSSD.n1116 0.120292
R14066 VSSD.n2926 VSSD.n2925 0.120292
R14067 VSSD.n2956 VSSD.n2955 0.120292
R14068 VSSD.n2963 VSSD.n1095 0.120292
R14069 VSSD.n2964 VSSD.n2963 0.120292
R14070 VSSD.n2965 VSSD.n1093 0.120292
R14071 VSSD.n2969 VSSD.n1093 0.120292
R14072 VSSD.n2970 VSSD.n2969 0.120292
R14073 VSSD.n2971 VSSD.n2970 0.120292
R14074 VSSD.n2971 VSSD.n1091 0.120292
R14075 VSSD.n2978 VSSD.n1091 0.120292
R14076 VSSD.n2979 VSSD.n2978 0.120292
R14077 VSSD.n2980 VSSD.n2979 0.120292
R14078 VSSD.n2980 VSSD.n1089 0.120292
R14079 VSSD.n2987 VSSD.n1089 0.120292
R14080 VSSD.n2988 VSSD.n2987 0.120292
R14081 VSSD.n3006 VSSD.n3005 0.120292
R14082 VSSD.n3012 VSSD.n3010 0.120292
R14083 VSSD.n3012 VSSD.n3011 0.120292
R14084 VSSD.n3051 VSSD.n3022 0.120292
R14085 VSSD.n3046 VSSD.n3022 0.120292
R14086 VSSD.n3046 VSSD.n3045 0.120292
R14087 VSSD.n3045 VSSD.n3024 0.120292
R14088 VSSD.n3032 VSSD.n3030 0.120292
R14089 VSSD.n3034 VSSD.n3032 0.120292
R14090 VSSD.n3034 VSSD.n3033 0.120292
R14091 VSSD.n3137 VSSD.n1065 0.120292
R14092 VSSD.n3131 VSSD.n1065 0.120292
R14093 VSSD.n3131 VSSD.n3130 0.120292
R14094 VSSD.n3130 VSSD.n3129 0.120292
R14095 VSSD.n3129 VSSD.n1069 0.120292
R14096 VSSD.n3124 VSSD.n1069 0.120292
R14097 VSSD.n3124 VSSD.n3123 0.120292
R14098 VSSD.n3123 VSSD.n1073 0.120292
R14099 VSSD.n1074 VSSD.n1073 0.120292
R14100 VSSD.n1075 VSSD.n1074 0.120292
R14101 VSSD.n1076 VSSD.n1075 0.120292
R14102 VSSD.n3109 VSSD.n3061 0.120292
R14103 VSSD.n3109 VSSD.n3108 0.120292
R14104 VSSD.n3108 VSSD.n3107 0.120292
R14105 VSSD.n3107 VSSD.n3064 0.120292
R14106 VSSD.n3103 VSSD.n3064 0.120292
R14107 VSSD.n3103 VSSD.n3102 0.120292
R14108 VSSD.n3102 VSSD.n3101 0.120292
R14109 VSSD.n3101 VSSD.n3066 0.120292
R14110 VSSD.n3096 VSSD.n3066 0.120292
R14111 VSSD.n3096 VSSD.n3095 0.120292
R14112 VSSD.n3095 VSSD.n3094 0.120292
R14113 VSSD.n3094 VSSD.n3070 0.120292
R14114 VSSD.n3090 VSSD.n3070 0.120292
R14115 VSSD.n3090 VSSD.n3089 0.120292
R14116 VSSD.n3089 VSSD.n3074 0.120292
R14117 VSSD.n3085 VSSD.n3074 0.120292
R14118 VSSD.n3085 VSSD.n3084 0.120292
R14119 VSSD.n3084 VSSD.n3083 0.120292
R14120 VSSD.n3083 VSSD.n3076 0.120292
R14121 VSSD.n2585 VSSD.n2584 0.120292
R14122 VSSD.n2586 VSSD.n2585 0.120292
R14123 VSSD.n2586 VSSD.n2544 0.120292
R14124 VSSD.n2590 VSSD.n2544 0.120292
R14125 VSSD.n2591 VSSD.n2590 0.120292
R14126 VSSD.n2591 VSSD.n2541 0.120292
R14127 VSSD.n2597 VSSD.n2541 0.120292
R14128 VSSD.n2598 VSSD.n2597 0.120292
R14129 VSSD.n2599 VSSD.n2598 0.120292
R14130 VSSD.n2599 VSSD.n2539 0.120292
R14131 VSSD.n2607 VSSD.n2539 0.120292
R14132 VSSD.n2608 VSSD.n2607 0.120292
R14133 VSSD.n2609 VSSD.n2608 0.120292
R14134 VSSD.n2609 VSSD.n2537 0.120292
R14135 VSSD.n2613 VSSD.n2537 0.120292
R14136 VSSD.n2614 VSSD.n2613 0.120292
R14137 VSSD.n2615 VSSD.n2614 0.120292
R14138 VSSD.n2688 VSSD.n2687 0.120292
R14139 VSSD.n2682 VSSD.n2681 0.120292
R14140 VSSD.n2681 VSSD.n2635 0.120292
R14141 VSSD.n2673 VSSD.n2635 0.120292
R14142 VSSD.n2673 VSSD.n2672 0.120292
R14143 VSSD.n2672 VSSD.n2638 0.120292
R14144 VSSD.n2665 VSSD.n2638 0.120292
R14145 VSSD.n2664 VSSD.n2641 0.120292
R14146 VSSD.n2657 VSSD.n2641 0.120292
R14147 VSSD.n2657 VSSD.n2656 0.120292
R14148 VSSD.n2656 VSSD.n2655 0.120292
R14149 VSSD.n2655 VSSD.n2645 0.120292
R14150 VSSD.n2650 VSSD.n2645 0.120292
R14151 VSSD.n2834 VSSD.n2833 0.120292
R14152 VSSD.n2830 VSSD.n2829 0.120292
R14153 VSSD.n2829 VSSD.n1328 0.120292
R14154 VSSD.n2823 VSSD.n1328 0.120292
R14155 VSSD.n1333 VSSD.n1330 0.120292
R14156 VSSD.n1334 VSSD.n1333 0.120292
R14157 VSSD.n2814 VSSD.n1338 0.120292
R14158 VSSD.n1342 VSSD.n1338 0.120292
R14159 VSSD.n1343 VSSD.n1342 0.120292
R14160 VSSD.n2807 VSSD.n1343 0.120292
R14161 VSSD.n2807 VSSD.n2806 0.120292
R14162 VSSD.n2806 VSSD.n2805 0.120292
R14163 VSSD.n2794 VSSD.n1359 0.120292
R14164 VSSD.n2788 VSSD.n2787 0.120292
R14165 VSSD.n2787 VSSD.n1365 0.120292
R14166 VSSD.n2782 VSSD.n1365 0.120292
R14167 VSSD.n2782 VSSD.n2781 0.120292
R14168 VSSD.n2781 VSSD.n2780 0.120292
R14169 VSSD.n2780 VSSD.n1368 0.120292
R14170 VSSD.n2774 VSSD.n1368 0.120292
R14171 VSSD.n2773 VSSD.n1370 0.120292
R14172 VSSD.n2764 VSSD.n2763 0.120292
R14173 VSSD.n2763 VSSD.n2699 0.120292
R14174 VSSD.n2758 VSSD.n2699 0.120292
R14175 VSSD.n2758 VSSD.n2757 0.120292
R14176 VSSD.n2757 VSSD.n2756 0.120292
R14177 VSSD.n2756 VSSD.n2702 0.120292
R14178 VSSD.n2752 VSSD.n2702 0.120292
R14179 VSSD.n2752 VSSD.n2751 0.120292
R14180 VSSD.n2751 VSSD.n2704 0.120292
R14181 VSSD.n2746 VSSD.n2704 0.120292
R14182 VSSD.n2746 VSSD.n2745 0.120292
R14183 VSSD.n2742 VSSD.n2741 0.120292
R14184 VSSD.n2741 VSSD.n2708 0.120292
R14185 VSSD.n2736 VSSD.n2708 0.120292
R14186 VSSD.n2736 VSSD.n2735 0.120292
R14187 VSSD.n2735 VSSD.n2734 0.120292
R14188 VSSD.n2734 VSSD.n2711 0.120292
R14189 VSSD.n2728 VSSD.n2711 0.120292
R14190 VSSD.n2727 VSSD.n2713 0.120292
R14191 VSSD.n2722 VSSD.n2713 0.120292
R14192 VSSD.n2722 VSSD.n2721 0.120292
R14193 VSSD.n1494 VSSD.n1493 0.120292
R14194 VSSD.n1495 VSSD.n1494 0.120292
R14195 VSSD.n1551 VSSD.n1550 0.120292
R14196 VSSD.n1550 VSSD.n1499 0.120292
R14197 VSSD.n1546 VSSD.n1499 0.120292
R14198 VSSD.n1546 VSSD.n1545 0.120292
R14199 VSSD.n1545 VSSD.n1504 0.120292
R14200 VSSD.n1540 VSSD.n1504 0.120292
R14201 VSSD.n1540 VSSD.n1539 0.120292
R14202 VSSD.n1539 VSSD.n1538 0.120292
R14203 VSSD.n1538 VSSD.n1507 0.120292
R14204 VSSD.n1508 VSSD.n1507 0.120292
R14205 VSSD.n1533 VSSD.n1508 0.120292
R14206 VSSD.n1533 VSSD.n1532 0.120292
R14207 VSSD.n1532 VSSD.n1510 0.120292
R14208 VSSD.n1526 VSSD.n1525 0.120292
R14209 VSSD.n1522 VSSD.n1521 0.120292
R14210 VSSD.n1521 VSSD.n1517 0.120292
R14211 VSSD.n2506 VSSD.n2505 0.120292
R14212 VSSD.n2505 VSSD.n2504 0.120292
R14213 VSSD.n2504 VSSD.n1386 0.120292
R14214 VSSD.n2498 VSSD.n1386 0.120292
R14215 VSSD.n2497 VSSD.n2496 0.120292
R14216 VSSD.n2492 VSSD.n1392 0.120292
R14217 VSSD.n2487 VSSD.n1392 0.120292
R14218 VSSD.n2487 VSSD.n2486 0.120292
R14219 VSSD.n2486 VSSD.n2485 0.120292
R14220 VSSD.n2485 VSSD.n1395 0.120292
R14221 VSSD.n2481 VSSD.n1395 0.120292
R14222 VSSD.n2481 VSSD.n2480 0.120292
R14223 VSSD.n2480 VSSD.n2479 0.120292
R14224 VSSD.n2465 VSSD.n1406 0.120292
R14225 VSSD.n2459 VSSD.n1406 0.120292
R14226 VSSD.n2324 VSSD.n2323 0.120292
R14227 VSSD.n2324 VSSD.n2316 0.120292
R14228 VSSD.n2331 VSSD.n2316 0.120292
R14229 VSSD.n2333 VSSD.n2313 0.120292
R14230 VSSD.n2340 VSSD.n2313 0.120292
R14231 VSSD.n2341 VSSD.n2340 0.120292
R14232 VSSD.n2342 VSSD.n2341 0.120292
R14233 VSSD.n2362 VSSD.n1424 0.120292
R14234 VSSD.n2363 VSSD.n2362 0.120292
R14235 VSSD.n2364 VSSD.n2363 0.120292
R14236 VSSD.n2364 VSSD.n1422 0.120292
R14237 VSSD.n2369 VSSD.n1422 0.120292
R14238 VSSD.n2374 VSSD.n2373 0.120292
R14239 VSSD.n2374 VSSD.n1418 0.120292
R14240 VSSD.n2381 VSSD.n1418 0.120292
R14241 VSSD.n2450 VSSD.n2449 0.120292
R14242 VSSD.n2449 VSSD.n2386 0.120292
R14243 VSSD.n2445 VSSD.n2386 0.120292
R14244 VSSD.n2445 VSSD.n2444 0.120292
R14245 VSSD.n2444 VSSD.n2443 0.120292
R14246 VSSD.n2443 VSSD.n2390 0.120292
R14247 VSSD.n2438 VSSD.n2390 0.120292
R14248 VSSD.n2438 VSSD.n2437 0.120292
R14249 VSSD.n2437 VSSD.n2393 0.120292
R14250 VSSD.n2433 VSSD.n2393 0.120292
R14251 VSSD.n2433 VSSD.n2432 0.120292
R14252 VSSD.n2427 VSSD.n2426 0.120292
R14253 VSSD.n2426 VSSD.n2396 0.120292
R14254 VSSD.n2422 VSSD.n2396 0.120292
R14255 VSSD.n2422 VSSD.n2421 0.120292
R14256 VSSD.n2421 VSSD.n2398 0.120292
R14257 VSSD.n2416 VSSD.n2415 0.120292
R14258 VSSD.n2415 VSSD.n2400 0.120292
R14259 VSSD.n2410 VSSD.n2400 0.120292
R14260 VSSD.n2410 VSSD.n2409 0.120292
R14261 VSSD.n2409 VSSD.n2408 0.120292
R14262 VSSD.n1978 VSSD.n1977 0.120292
R14263 VSSD.n1990 VSSD.n1467 0.120292
R14264 VSSD.n1995 VSSD.n1467 0.120292
R14265 VSSD.n1996 VSSD.n1995 0.120292
R14266 VSSD.n1997 VSSD.n1996 0.120292
R14267 VSSD.n1997 VSSD.n1464 0.120292
R14268 VSSD.n2004 VSSD.n1464 0.120292
R14269 VSSD.n2005 VSSD.n2004 0.120292
R14270 VSSD.n2006 VSSD.n2005 0.120292
R14271 VSSD.n2006 VSSD.n1462 0.120292
R14272 VSSD.n2010 VSSD.n1462 0.120292
R14273 VSSD.n2011 VSSD.n2010 0.120292
R14274 VSSD.n2012 VSSD.n2011 0.120292
R14275 VSSD.n2012 VSSD.n1459 0.120292
R14276 VSSD.n2018 VSSD.n1459 0.120292
R14277 VSSD.n2028 VSSD.n1456 0.120292
R14278 VSSD.n2102 VSSD.n2101 0.120292
R14279 VSSD.n2101 VSSD.n2049 0.120292
R14280 VSSD.n2095 VSSD.n2049 0.120292
R14281 VSSD.n2095 VSSD.n2094 0.120292
R14282 VSSD.n2094 VSSD.n2053 0.120292
R14283 VSSD.n2088 VSSD.n2053 0.120292
R14284 VSSD.n2088 VSSD.n2087 0.120292
R14285 VSSD.n2087 VSSD.n2086 0.120292
R14286 VSSD.n2086 VSSD.n2057 0.120292
R14287 VSSD.n2082 VSSD.n2057 0.120292
R14288 VSSD.n2082 VSSD.n2081 0.120292
R14289 VSSD.n2081 VSSD.n2063 0.120292
R14290 VSSD.n2065 VSSD.n2063 0.120292
R14291 VSSD.n2075 VSSD.n2074 0.120292
R14292 VSSD.n2074 VSSD.n2067 0.120292
R14293 VSSD.n2284 VSSD.n1447 0.120292
R14294 VSSD.n2275 VSSD.n2274 0.120292
R14295 VSSD.n2274 VSSD.n2110 0.120292
R14296 VSSD.n2270 VSSD.n2110 0.120292
R14297 VSSD.n2270 VSSD.n2269 0.120292
R14298 VSSD.n2269 VSSD.n2268 0.120292
R14299 VSSD.n2268 VSSD.n2112 0.120292
R14300 VSSD.n2261 VSSD.n2112 0.120292
R14301 VSSD.n2259 VSSD.n2119 0.120292
R14302 VSSD.n2238 VSSD.n2128 0.120292
R14303 VSSD.n2234 VSSD.n2233 0.120292
R14304 VSSD.n2232 VSSD.n2130 0.120292
R14305 VSSD.n2227 VSSD.n2130 0.120292
R14306 VSSD.n2227 VSSD.n2226 0.120292
R14307 VSSD.n2226 VSSD.n2225 0.120292
R14308 VSSD.n2225 VSSD.n2134 0.120292
R14309 VSSD.n2218 VSSD.n2134 0.120292
R14310 VSSD.n2218 VSSD.n2217 0.120292
R14311 VSSD.n2208 VSSD.n2146 0.120292
R14312 VSSD.n2147 VSSD.n2146 0.120292
R14313 VSSD.n2202 VSSD.n2147 0.120292
R14314 VSSD.n2202 VSSD.n2201 0.120292
R14315 VSSD.n2201 VSSD.n2200 0.120292
R14316 VSSD.n2200 VSSD.n2149 0.120292
R14317 VSSD.n2195 VSSD.n2149 0.120292
R14318 VSSD.n2195 VSSD.n2194 0.120292
R14319 VSSD.n2194 VSSD.n2193 0.120292
R14320 VSSD.n2193 VSSD.n2152 0.120292
R14321 VSSD.n2189 VSSD.n2152 0.120292
R14322 VSSD.n2189 VSSD.n2188 0.120292
R14323 VSSD.n2188 VSSD.n2157 0.120292
R14324 VSSD.n2183 VSSD.n2157 0.120292
R14325 VSSD.n2183 VSSD.n2182 0.120292
R14326 VSSD.n2182 VSSD.n2181 0.120292
R14327 VSSD.n2181 VSSD.n2160 0.120292
R14328 VSSD.n2175 VSSD.n2174 0.120292
R14329 VSSD.n2171 VSSD.n2170 0.120292
R14330 VSSD.n1613 VSSD.n1606 0.120292
R14331 VSSD.n1606 VSSD.n1605 0.120292
R14332 VSSD.n1936 VSSD.n1935 0.120292
R14333 VSSD.n1935 VSSD.n1577 0.120292
R14334 VSSD.n1931 VSSD.n1577 0.120292
R14335 VSSD.n1931 VSSD.n1930 0.120292
R14336 VSSD.n1930 VSSD.n1929 0.120292
R14337 VSSD.n1929 VSSD.n1581 0.120292
R14338 VSSD.n1923 VSSD.n1581 0.120292
R14339 VSSD.n1923 VSSD.n1922 0.120292
R14340 VSSD.n1922 VSSD.n1921 0.120292
R14341 VSSD.n1918 VSSD.n1917 0.120292
R14342 VSSD.n1917 VSSD.n1586 0.120292
R14343 VSSD.n1912 VSSD.n1586 0.120292
R14344 VSSD.n1912 VSSD.n1911 0.120292
R14345 VSSD.n1911 VSSD.n1910 0.120292
R14346 VSSD.n1907 VSSD.n1906 0.120292
R14347 VSSD.n1906 VSSD.n1591 0.120292
R14348 VSSD.n1886 VSSD.n1885 0.120292
R14349 VSSD.n1884 VSSD.n1627 0.120292
R14350 VSSD.n1878 VSSD.n1627 0.120292
R14351 VSSD.n1878 VSSD.n1877 0.120292
R14352 VSSD.n1877 VSSD.n1876 0.120292
R14353 VSSD.n1876 VSSD.n1629 0.120292
R14354 VSSD.n1870 VSSD.n1629 0.120292
R14355 VSSD.n1870 VSSD.n1869 0.120292
R14356 VSSD.n1869 VSSD.n1868 0.120292
R14357 VSSD.n1868 VSSD.n1633 0.120292
R14358 VSSD.n1864 VSSD.n1633 0.120292
R14359 VSSD.n1864 VSSD.n1863 0.120292
R14360 VSSD.n1863 VSSD.n1636 0.120292
R14361 VSSD.n1859 VSSD.n1636 0.120292
R14362 VSSD.n1859 VSSD.n1858 0.120292
R14363 VSSD.n1858 VSSD.n1857 0.120292
R14364 VSSD.n1844 VSSD.n1645 0.120292
R14365 VSSD.n1839 VSSD.n1838 0.120292
R14366 VSSD.n1838 VSSD.n1837 0.120292
R14367 VSSD.n1826 VSSD.n1825 0.120292
R14368 VSSD.n1825 VSSD.n1659 0.120292
R14369 VSSD.n1818 VSSD.n1659 0.120292
R14370 VSSD.n1818 VSSD.n1817 0.120292
R14371 VSSD.n1813 VSSD.n1667 0.120292
R14372 VSSD.n1809 VSSD.n1667 0.120292
R14373 VSSD.n1809 VSSD.n1808 0.120292
R14374 VSSD.n1808 VSSD.n1807 0.120292
R14375 VSSD.n1794 VSSD.n1684 0.120292
R14376 VSSD.n1788 VSSD.n1684 0.120292
R14377 VSSD.n1788 VSSD.n1787 0.120292
R14378 VSSD.n1787 VSSD.n1786 0.120292
R14379 VSSD.n1786 VSSD.n1687 0.120292
R14380 VSSD.n1780 VSSD.n1687 0.120292
R14381 VSSD.n1778 VSSD.n1691 0.120292
R14382 VSSD.n1772 VSSD.n1691 0.120292
R14383 VSSD.n1772 VSSD.n1771 0.120292
R14384 VSSD.n1760 VSSD.n1698 0.120292
R14385 VSSD.n1760 VSSD.n1759 0.120292
R14386 VSSD.n1759 VSSD.n1758 0.120292
R14387 VSSD.n1758 VSSD.n1699 0.120292
R14388 VSSD.n1754 VSSD.n1699 0.120292
R14389 VSSD.n1754 VSSD.n1753 0.120292
R14390 VSSD.n1753 VSSD.n1752 0.120292
R14391 VSSD.n1752 VSSD.n1702 0.120292
R14392 VSSD.n1746 VSSD.n1702 0.120292
R14393 VSSD.n1746 VSSD.n1745 0.120292
R14394 VSSD.n1745 VSSD.n1744 0.120292
R14395 VSSD.n1741 VSSD.n1740 0.120292
R14396 VSSD.n1740 VSSD.n1707 0.120292
R14397 VSSD.n1735 VSSD.n1707 0.120292
R14398 VSSD.n1735 VSSD.n1734 0.120292
R14399 VSSD.n1734 VSSD.n1733 0.120292
R14400 VSSD.n1733 VSSD.n1710 0.120292
R14401 VSSD.n1727 VSSD.n1710 0.120292
R14402 VSSD.n1726 VSSD.n1712 0.120292
R14403 VSSD.n1721 VSSD.n1712 0.120292
R14404 VSSD.n1721 VSSD.n1720 0.120292
R14405 VSSD.n3405 VSSD.n3399 0.120292
R14406 VSSD.n3413 VSSD.n131 0.120292
R14407 VSSD.n3414 VSSD.n3413 0.120292
R14408 VSSD.n3431 VSSD.n119 0.120292
R14409 VSSD.n3432 VSSD.n3431 0.120292
R14410 VSSD.n3433 VSSD.n3432 0.120292
R14411 VSSD.n3433 VSSD.n117 0.120292
R14412 VSSD.n3437 VSSD.n117 0.120292
R14413 VSSD.n3438 VSSD.n3437 0.120292
R14414 VSSD.n3438 VSSD.n115 0.120292
R14415 VSSD.n3442 VSSD.n115 0.120292
R14416 VSSD.n3443 VSSD.n3442 0.120292
R14417 VSSD.n3447 VSSD.n3446 0.120292
R14418 VSSD.n3447 VSSD.n112 0.120292
R14419 VSSD.n3451 VSSD.n112 0.120292
R14420 VSSD.n3452 VSSD.n3451 0.120292
R14421 VSSD.n3453 VSSD.n3452 0.120292
R14422 VSSD.n3453 VSSD.n110 0.120292
R14423 VSSD.n3457 VSSD.n110 0.120292
R14424 VSSD.n3458 VSSD.n3457 0.120292
R14425 VSSD.n3478 VSSD.n94 0.120292
R14426 VSSD.n3479 VSSD.n3478 0.120292
R14427 VSSD.n3483 VSSD.n3482 0.120292
R14428 VSSD.n3483 VSSD.n91 0.120292
R14429 VSSD.n3487 VSSD.n91 0.120292
R14430 VSSD.n3488 VSSD.n3487 0.120292
R14431 VSSD.n3489 VSSD.n3488 0.120292
R14432 VSSD.n3489 VSSD.n89 0.120292
R14433 VSSD.n3493 VSSD.n89 0.120292
R14434 VSSD.n3494 VSSD.n3493 0.120292
R14435 VSSD.n3494 VSSD.n87 0.120292
R14436 VSSD.n3498 VSSD.n87 0.120292
R14437 VSSD.n3499 VSSD.n3498 0.120292
R14438 VSSD.n3504 VSSD.n3503 0.120292
R14439 VSSD.n3505 VSSD.n3504 0.120292
R14440 VSSD.n3525 VSSD.n76 0.120292
R14441 VSSD.n3526 VSSD.n3525 0.120292
R14442 VSSD.n3526 VSSD.n74 0.120292
R14443 VSSD.n3531 VSSD.n74 0.120292
R14444 VSSD.n3532 VSSD.n3531 0.120292
R14445 VSSD.n3539 VSSD.n71 0.120292
R14446 VSSD.n3540 VSSD.n3539 0.120292
R14447 VSSD.n3544 VSSD.n3543 0.120292
R14448 VSSD.n3544 VSSD.n68 0.120292
R14449 VSSD.n3548 VSSD.n68 0.120292
R14450 VSSD.n3549 VSSD.n3548 0.120292
R14451 VSSD.n3550 VSSD.n3549 0.120292
R14452 VSSD.n3550 VSSD.n66 0.120292
R14453 VSSD.n3554 VSSD.n66 0.120292
R14454 VSSD.n3555 VSSD.n3554 0.120292
R14455 VSSD.n3573 VSSD.n3572 0.120292
R14456 VSSD.n3573 VSSD.n52 0.120292
R14457 VSSD.n3577 VSSD.n52 0.120292
R14458 VSSD.n3578 VSSD.n3577 0.120292
R14459 VSSD.n3579 VSSD.n3578 0.120292
R14460 VSSD.n3579 VSSD.n50 0.120292
R14461 VSSD.n3583 VSSD.n50 0.120292
R14462 VSSD.n3584 VSSD.n3583 0.120292
R14463 VSSD.n3584 VSSD.n48 0.120292
R14464 VSSD.n3589 VSSD.n48 0.120292
R14465 VSSD.n3590 VSSD.n3589 0.120292
R14466 VSSD.n3653 VSSD.n3652 0.120292
R14467 VSSD.n3652 VSSD.n3593 0.120292
R14468 VSSD.n3648 VSSD.n3593 0.120292
R14469 VSSD.n3648 VSSD.n3647 0.120292
R14470 VSSD.n3647 VSSD.n3646 0.120292
R14471 VSSD.n3646 VSSD.n3596 0.120292
R14472 VSSD.n3642 VSSD.n3596 0.120292
R14473 VSSD.n3642 VSSD.n3641 0.120292
R14474 VSSD.n3641 VSSD.n3598 0.120292
R14475 VSSD.n3637 VSSD.n3598 0.120292
R14476 VSSD.n3637 VSSD.n3636 0.120292
R14477 VSSD.n3633 VSSD.n3632 0.120292
R14478 VSSD.n3632 VSSD.n3601 0.120292
R14479 VSSD.n3628 VSSD.n3601 0.120292
R14480 VSSD.n3628 VSSD.n3627 0.120292
R14481 VSSD.n3627 VSSD.n3626 0.120292
R14482 VSSD.n3626 VSSD.n3603 0.120292
R14483 VSSD.n3622 VSSD.n3603 0.120292
R14484 VSSD.n3622 VSSD.n3621 0.120292
R14485 VSSD.n3621 VSSD.n3605 0.120292
R14486 VSSD.n3617 VSSD.n3605 0.120292
R14487 VSSD.n3617 VSSD.n3616 0.120292
R14488 VSSD.n3613 VSSD.n3612 0.120292
R14489 VSSD.n3612 VSSD.n3608 0.120292
R14490 VSSD.n486 VSSD.n485 0.120292
R14491 VSSD.n485 VSSD.n484 0.120292
R14492 VSSD.n473 VSSD.n153 0.120292
R14493 VSSD.n467 VSSD.n153 0.120292
R14494 VSSD.n467 VSSD.n466 0.120292
R14495 VSSD.n466 VSSD.n465 0.120292
R14496 VSSD.n465 VSSD.n157 0.120292
R14497 VSSD.n457 VSSD.n157 0.120292
R14498 VSSD.n457 VSSD.n456 0.120292
R14499 VSSD.n456 VSSD.n455 0.120292
R14500 VSSD.n455 VSSD.n159 0.120292
R14501 VSSD.n451 VSSD.n159 0.120292
R14502 VSSD.n451 VSSD.n450 0.120292
R14503 VSSD.n450 VSSD.n449 0.120292
R14504 VSSD.n449 VSSD.n161 0.120292
R14505 VSSD.n443 VSSD.n161 0.120292
R14506 VSSD.n437 VSSD.n436 0.120292
R14507 VSSD.n416 VSSD.n182 0.120292
R14508 VSSD.n414 VSSD.n183 0.120292
R14509 VSSD.n410 VSSD.n183 0.120292
R14510 VSSD.n410 VSSD.n409 0.120292
R14511 VSSD.n409 VSSD.n186 0.120292
R14512 VSSD.n405 VSSD.n186 0.120292
R14513 VSSD.n405 VSSD.n404 0.120292
R14514 VSSD.n404 VSSD.n403 0.120292
R14515 VSSD.n403 VSSD.n190 0.120292
R14516 VSSD.n397 VSSD.n190 0.120292
R14517 VSSD.n397 VSSD.n396 0.120292
R14518 VSSD.n396 VSSD.n395 0.120292
R14519 VSSD.n395 VSSD.n194 0.120292
R14520 VSSD.n391 VSSD.n194 0.120292
R14521 VSSD.n391 VSSD.n390 0.120292
R14522 VSSD.n373 VSSD.n372 0.120292
R14523 VSSD.n372 VSSD.n213 0.120292
R14524 VSSD.n365 VSSD.n213 0.120292
R14525 VSSD.n359 VSSD.n215 0.120292
R14526 VSSD.n359 VSSD.n358 0.120292
R14527 VSSD.n358 VSSD.n219 0.120292
R14528 VSSD.n353 VSSD.n219 0.120292
R14529 VSSD.n353 VSSD.n352 0.120292
R14530 VSSD.n352 VSSD.n351 0.120292
R14531 VSSD.n351 VSSD.n221 0.120292
R14532 VSSD.n346 VSSD.n221 0.120292
R14533 VSSD.n346 VSSD.n345 0.120292
R14534 VSSD.n345 VSSD.n225 0.120292
R14535 VSSD.n333 VSSD.n238 0.120292
R14536 VSSD.n328 VSSD.n238 0.120292
R14537 VSSD.n328 VSSD.n327 0.120292
R14538 VSSD.n327 VSSD.n326 0.120292
R14539 VSSD.n326 VSSD.n243 0.120292
R14540 VSSD.n321 VSSD.n320 0.120292
R14541 VSSD.n320 VSSD.n246 0.120292
R14542 VSSD.n315 VSSD.n246 0.120292
R14543 VSSD.n309 VSSD.n308 0.120292
R14544 VSSD.n308 VSSD.n254 0.120292
R14545 VSSD.n304 VSSD.n254 0.120292
R14546 VSSD.n304 VSSD.n303 0.120292
R14547 VSSD.n303 VSSD.n302 0.120292
R14548 VSSD.n302 VSSD.n256 0.120292
R14549 VSSD.n298 VSSD.n256 0.120292
R14550 VSSD.n298 VSSD.n297 0.120292
R14551 VSSD.n297 VSSD.n258 0.120292
R14552 VSSD.n293 VSSD.n258 0.120292
R14553 VSSD.n293 VSSD.n292 0.120292
R14554 VSSD.n289 VSSD.n288 0.120292
R14555 VSSD.n288 VSSD.n261 0.120292
R14556 VSSD.n284 VSSD.n261 0.120292
R14557 VSSD.n284 VSSD.n283 0.120292
R14558 VSSD.n283 VSSD.n282 0.120292
R14559 VSSD.n282 VSSD.n263 0.120292
R14560 VSSD.n278 VSSD.n263 0.120292
R14561 VSSD.n278 VSSD.n277 0.120292
R14562 VSSD.n277 VSSD.n265 0.120292
R14563 VSSD.n273 VSSD.n265 0.120292
R14564 VSSD.n273 VSSD.n272 0.120292
R14565 VSSD.n655 VSSD.n581 0.120292
R14566 VSSD.n648 VSSD.n581 0.120292
R14567 VSSD.n648 VSSD.n647 0.120292
R14568 VSSD.n644 VSSD.n643 0.120292
R14569 VSSD.n643 VSSD.n587 0.120292
R14570 VSSD.n638 VSSD.n587 0.120292
R14571 VSSD.n638 VSSD.n637 0.120292
R14572 VSSD.n637 VSSD.n636 0.120292
R14573 VSSD.n633 VSSD.n632 0.120292
R14574 VSSD.n632 VSSD.n591 0.120292
R14575 VSSD.n627 VSSD.n591 0.120292
R14576 VSSD.n627 VSSD.n626 0.120292
R14577 VSSD.n626 VSSD.n625 0.120292
R14578 VSSD.n622 VSSD.n621 0.120292
R14579 VSSD.n621 VSSD.n595 0.120292
R14580 VSSD.n682 VSSD.n552 0.120292
R14581 VSSD.n683 VSSD.n682 0.120292
R14582 VSSD.n684 VSSD.n683 0.120292
R14583 VSSD.n684 VSSD.n550 0.120292
R14584 VSSD.n689 VSSD.n550 0.120292
R14585 VSSD.n690 VSSD.n689 0.120292
R14586 VSSD.n690 VSSD.n547 0.120292
R14587 VSSD.n694 VSSD.n547 0.120292
R14588 VSSD.n695 VSSD.n694 0.120292
R14589 VSSD.n702 VSSD.n701 0.120292
R14590 VSSD.n703 VSSD.n702 0.120292
R14591 VSSD.n720 VSSD.n719 0.120292
R14592 VSSD.n719 VSSD.n708 0.120292
R14593 VSSD.n714 VSSD.n708 0.120292
R14594 VSSD.n714 VSSD 0.120292
R14595 VSSD.n3672 VSSD.n40 0.120292
R14596 VSSD.n3680 VSSD.n40 0.120292
R14597 VSSD.n3681 VSSD.n3680 0.120292
R14598 VSSD.n3685 VSSD.n38 0.120292
R14599 VSSD.n3686 VSSD.n3685 0.120292
R14600 VSSD.n3687 VSSD.n3686 0.120292
R14601 VSSD.n3687 VSSD.n36 0.120292
R14602 VSSD.n3693 VSSD.n36 0.120292
R14603 VSSD.n3694 VSSD.n3693 0.120292
R14604 VSSD.n3715 VSSD.n3714 0.120292
R14605 VSSD.n3716 VSSD.n3715 0.120292
R14606 VSSD.n3716 VSSD.n20 0.120292
R14607 VSSD.n3720 VSSD.n20 0.120292
R14608 VSSD.n3721 VSSD.n3720 0.120292
R14609 VSSD.n3722 VSSD.n18 0.120292
R14610 VSSD.n3726 VSSD.n18 0.120292
R14611 VSSD.n3727 VSSD.n3726 0.120292
R14612 VSSD.n3728 VSSD.n3727 0.120292
R14613 VSSD.n3740 VSSD.n3739 0.120292
R14614 VSSD.n3741 VSSD.n3740 0.120292
R14615 VSSD.n3741 VSSD.n12 0.120292
R14616 VSSD.n3746 VSSD.n12 0.120292
R14617 VSSD.n3747 VSSD.n3746 0.120292
R14618 VSSD.n3748 VSSD.n3747 0.120292
R14619 VSSD.n3748 VSSD.n10 0.120292
R14620 VSSD.n3753 VSSD.n10 0.120292
R14621 VSSD.n3754 VSSD.n3753 0.120292
R14622 VSSD.n3754 VSSD.n8 0.120292
R14623 VSSD.n3762 VSSD.n8 0.120292
R14624 VSSD.n3770 VSSD.n6 0.120292
R14625 VSSD.n3771 VSSD.n3770 0.120292
R14626 VSSD.n3775 VSSD.n3774 0.120292
R14627 VSSD.n3775 VSSD.n3 0.120292
R14628 VSSD.n3779 VSSD.n3 0.120292
R14629 VSSD.n3780 VSSD.n3779 0.120292
R14630 VSSD.n3780 VSSD.n1 0.120292
R14631 VSSD.n3785 VSSD.n1 0.120292
R14632 VSSD.n3786 VSSD.n3785 0.120292
R14633 VSSD.n3138 VSSD.n3137 0.117688
R14634 VSSD.n2795 VSSD.n2794 0.117688
R14635 VSSD.n2353 VSSD.n1424 0.117688
R14636 VSSD.n2239 VSSD.n2238 0.117688
R14637 VSSD.n1795 VSSD.n1794 0.117688
R14638 VSSD.n3714 VSSD.n22 0.117688
R14639 VSSD.n137 VSSD 0.105581
R14640 VSSD.n493 VSSD 0.105238
R14641 VSSD.n1141 VSSD 0.105238
R14642 VSSD.n2866 VSSD 0.105238
R14643 VSSD.n2560 VSSD 0.105238
R14644 VSSD.n1486 VSSD 0.105238
R14645 VSSD.n1967 VSSD 0.105238
R14646 VSSD.n1603 VSSD 0.105238
R14647 VSSD.n564 VSSD 0.105238
R14648 VSSD.n2304 VSSD.n1429 0.103624
R14649 VSSD.n2301 VSSD.n2300 0.103624
R14650 VSSD.n2042 VSSD.n1375 0.103624
R14651 VSSD.n1986 VSSD.n1569 0.103624
R14652 VSSD.n3354 VSSD 0.0981562
R14653 VSSD VSSD.n977 0.0981562
R14654 VSSD.n867 VSSD 0.0981562
R14655 VSSD VSSD.n1284 0.0981562
R14656 VSSD VSSD.n1266 0.0981562
R14657 VSSD.n3183 VSSD 0.0981562
R14658 VSSD.n3277 VSSD 0.0981562
R14659 VSSD.n2930 VSSD 0.0981562
R14660 VSSD VSSD.n1095 0.0981562
R14661 VSSD.n3030 VSSD 0.0981562
R14662 VSSD.n3061 VSSD 0.0981562
R14663 VSSD VSSD.n2688 0.0981562
R14664 VSSD VSSD.n2682 0.0981562
R14665 VSSD VSSD.n2814 0.0981562
R14666 VSSD.n2764 VSSD 0.0981562
R14667 VSSD.n2742 VSSD 0.0981562
R14668 VSSD VSSD.n2492 0.0981562
R14669 VSSD.n2333 VSSD 0.0981562
R14670 VSSD.n2427 VSSD 0.0981562
R14671 VSSD VSSD.n2284 0.0981562
R14672 VSSD.n2279 VSSD 0.0981562
R14673 VSSD VSSD.n2259 0.0981562
R14674 VSSD.n2143 VSSD 0.0981562
R14675 VSSD VSSD.n2208 0.0981562
R14676 VSSD.n1918 VSSD 0.0981562
R14677 VSSD VSSD.n1813 0.0981562
R14678 VSSD.n1741 VSSD 0.0981562
R14679 VSSD VSSD.n3399 0.0981562
R14680 VSSD.n3446 VSSD 0.0981562
R14681 VSSD.n3503 VSSD 0.0981562
R14682 VSSD.n3533 VSSD 0.0981562
R14683 VSSD.n3572 VSSD 0.0981562
R14684 VSSD.n3591 VSSD 0.0981562
R14685 VSSD.n3633 VSSD 0.0981562
R14686 VSSD.n3613 VSSD 0.0981562
R14687 VSSD VSSD.n414 0.0981562
R14688 VSSD.n211 VSSD 0.0981562
R14689 VSSD.n215 VSSD 0.0981562
R14690 VSSD VSSD.n312 0.0981562
R14691 VSSD.n289 VSSD 0.0981562
R14692 VSSD.n633 VSSD 0.0981562
R14693 VSSD.n622 VSSD 0.0981562
R14694 VSSD VSSD.n552 0.0981562
R14695 VSSD.n701 VSSD 0.0981562
R14696 VSSD.n3763 VSSD 0.0981562
R14697 VSSD VSSD.n1283 0.0968542
R14698 VSSD.n2931 VSSD 0.0968542
R14699 VSSD.n1330 VSSD 0.0968542
R14700 VSSD.n1052 VSSD.n28 0.0964353
R14701 VSSD.n3333 VSSD.n1013 0.0964353
R14702 VSSD.n3337 VSSD.n3336 0.0964353
R14703 VSSD.n534 VSSD.n510 0.0964353
R14704 VSSD.n577 VSSD.n576 0.0950946
R14705 VSSD.n657 VSSD.n573 0.0950946
R14706 VSSD.n614 VSSD.n600 0.0950946
R14707 VSSD.n608 VSSD.n603 0.0950946
R14708 VSSD.n431 VSSD.n167 0.0950946
R14709 VSSD.n425 VSSD.n170 0.0950946
R14710 VSSD.n732 VSSD.n731 0.0950946
R14711 VSSD.n725 VSSD.n543 0.0950946
R14712 VSSD.n385 VSSD.n202 0.0950946
R14713 VSSD.n379 VSSD.n205 0.0950946
R14714 VSSD.n3700 VSSD.n3699 0.0950946
R14715 VSSD.n3705 VSSD.n3704 0.0950946
R14716 VSSD.n1011 VSSD.n1010 0.0950946
R14717 VSSD.n1004 VSSD.n741 0.0950946
R14718 VSSD.n3339 VSSD.n529 0.0950946
R14719 VSSD.n766 VSSD.n765 0.0950946
R14720 VSSD.n508 VSSD.n507 0.0950946
R14721 VSSD.n3379 VSSD.n504 0.0950946
R14722 VSSD.n964 VSSD.n840 0.0950946
R14723 VSSD.n959 VSSD.n843 0.0950946
R14724 VSSD.n3330 VSSD.n3329 0.0950946
R14725 VSSD.n3323 VSSD.n1020 0.0950946
R14726 VSSD.n1211 VSSD.n1209 0.0950946
R14727 VSSD.n1226 VSSD.n1149 0.0950946
R14728 VSSD.n1308 VSSD.n1307 0.0950946
R14729 VSSD.n1173 VSSD.n1172 0.0950946
R14730 VSSD.n3197 VSSD.n3196 0.0950946
R14731 VSSD.n3201 VSSD.n1050 0.0950946
R14732 VSSD.n2991 VSSD.n2989 0.0950946
R14733 VSSD.n3003 VSSD.n1083 0.0950946
R14734 VSSD.n2944 VSSD.n2943 0.0950946
R14735 VSSD.n2948 VSSD.n1102 0.0950946
R14736 VSSD.n2887 VSSD.n2886 0.0950946
R14737 VSSD.n2891 VSSD.n1130 0.0950946
R14738 VSSD.n3148 VSSD.n3147 0.0950946
R14739 VSSD.n3140 VSSD.n3139 0.0950946
R14740 VSSD.n2846 VSSD.n2845 0.0950946
R14741 VSSD.n2839 VSSD.n1320 0.0950946
R14742 VSSD.n2624 VSSD.n2623 0.0950946
R14743 VSSD.n2628 VSSD.n1372 0.0950946
R14744 VSSD.n2556 VSSD.n2554 0.0950946
R14745 VSSD.n2579 VSSD.n2548 0.0950946
R14746 VSSD.n1354 VSSD.n1353 0.0950946
R14747 VSSD.n2796 VSSD.n1351 0.0950946
R14748 VSSD.n2473 VSSD.n1402 0.0950946
R14749 VSSD.n2467 VSSD.n1405 0.0950946
R14750 VSSD.n2524 VSSD.n2523 0.0950946
R14751 VSSD.n2515 VSSD.n2514 0.0950946
R14752 VSSD.n1566 VSSD.n1565 0.0950946
R14753 VSSD.n1557 VSSD.n1556 0.0950946
R14754 VSSD.n2348 VSSD.n2347 0.0950946
R14755 VSSD.n2352 VSSD.n1427 0.0950946
R14756 VSSD.n2298 VSSD.n2297 0.0950946
R14757 VSSD.n2291 VSSD.n1438 0.0950946
R14758 VSSD.n2040 VSSD.n2039 0.0950946
R14759 VSSD.n2044 VSSD.n1452 0.0950946
R14760 VSSD.n1984 VSSD.n1983 0.0950946
R14761 VSSD.n1988 VSSD.n1472 0.0950946
R14762 VSSD.n2245 VSSD.n2244 0.0950946
R14763 VSSD.n2251 VSSD.n2250 0.0950946
R14764 VSSD.n1852 VSSD.n1640 0.0950946
R14765 VSSD.n1846 VSSD.n1643 0.0950946
R14766 VSSD.n1897 VSSD.n1594 0.0950946
R14767 VSSD.n1891 VSSD.n1597 0.0950946
R14768 VSSD.n1951 VSSD.n1950 0.0950946
R14769 VSSD.n1942 VSSD.n1941 0.0950946
R14770 VSSD.n1679 VSSD.n1678 0.0950946
R14771 VSSD.n1796 VSSD.n1676 0.0950946
R14772 VSSD.n233 VSSD.n232 0.0950946
R14773 VSSD.n335 VSSD.n230 0.0950946
R14774 VSSD.n3515 VSSD.n3514 0.0950946
R14775 VSSD.n3519 VSSD.n79 0.0950946
R14776 VSSD.n3466 VSSD.n3465 0.0950946
R14777 VSSD.n3470 VSSD.n97 0.0950946
R14778 VSSD.n3420 VSSD.n3419 0.0950946
R14779 VSSD.n3425 VSSD.n3424 0.0950946
R14780 VSSD.n3563 VSSD.n3562 0.0950946
R14781 VSSD.n3567 VSSD.n56 0.0950946
R14782 VSSD.n148 VSSD.n147 0.0950946
R14783 VSSD.n475 VSSD.n146 0.0950946
R14784 VSSD.n3341 VSSD.n3340 0.0916458
R14785 VSSD.n1212 VSSD.n1208 0.0916458
R14786 VSSD.n2931 VSSD.n1106 0.0916458
R14787 VSSD.n2615 VSSD.n2528 0.0916458
R14788 VSSD.n1517 VSSD.n1377 0.0916458
R14789 VSSD.n2029 VSSD.n2028 0.0916458
R14790 VSSD.n1593 VSSD.n1591 0.0916458
R14791 VSSD.n3458 VSSD.n101 0.0916458
R14792 VSSD.n436 VSSD.n164 0.0916458
R14793 VSSD.n598 VSSD.n595 0.0916458
R14794 VSSD.n3761 VSSD.n3760 0.0900105
R14795 VSSD.n3317 VSSD.n1021 0.0864375
R14796 VSSD.n3005 VSSD.n3004 0.0864375
R14797 VSSD.n2834 VSSD.n1321 0.0864375
R14798 VSSD.n1845 VSSD.n1844 0.0864375
R14799 VSSD.n3520 VSSD.n76 0.0864375
R14800 VSSD.n720 VSSD.n544 0.0864375
R14801 VSSD.n506 VSSD.n502 0.0838333
R14802 VSSD.n3378 VSSD.n511 0.0838333
R14803 VSSD.n764 VSSD.n757 0.0838333
R14804 VSSD.n1009 VSSD.n1008 0.0838333
R14805 VSSD.n965 VSSD.n839 0.0838333
R14806 VSSD.n1306 VSSD.n1134 0.0838333
R14807 VSSD.n1174 VSSD.n1168 0.0838333
R14808 VSSD.n1221 VSSD.n1220 0.0838333
R14809 VSSD.n2892 VSSD.n1129 0.0838333
R14810 VSSD.n2936 VSSD.n1111 0.0838333
R14811 VSSD.n2998 VSSD.n1086 0.0838333
R14812 VSSD.n3146 VSSD.n1056 0.0838333
R14813 VSSD.n2557 VSSD.n2553 0.0838333
R14814 VSSD.n2844 VSSD.n2843 0.0838333
R14815 VSSD.n1564 VSSD.n1476 0.0838333
R14816 VSSD.n1558 VSSD.n1552 0.0838333
R14817 VSSD.n1383 VSSD.n1380 0.0838333
R14818 VSSD.n2474 VSSD.n1401 0.0838333
R14819 VSSD.n2346 VSSD.n2306 0.0838333
R14820 VSSD.n1982 VSSD.n1955 0.0838333
R14821 VSSD.n1989 VSSD.n1471 0.0838333
R14822 VSSD.n2036 VSSD.n2033 0.0838333
R14823 VSSD.n2296 VSSD.n2295 0.0838333
R14824 VSSD.n2243 VSSD.n2242 0.0838333
R14825 VSSD.n1943 VSSD.n1937 0.0838333
R14826 VSSD.n1622 VSSD.n1621 0.0838333
R14827 VSSD.n1673 VSSD.n1671 0.0838333
R14828 VSSD.n3426 VSSD.n122 0.0838333
R14829 VSSD.n108 VSSD.n105 0.0838333
R14830 VSSD.n3513 VSSD.n3512 0.0838333
R14831 VSSD.n3561 VSSD.n60 0.0838333
R14832 VSSD.n143 VSSD.n141 0.0838333
R14833 VSSD.n474 VSSD.n152 0.0838333
R14834 VSSD.n174 VSSD.n173 0.0838333
R14835 VSSD.n386 VSSD.n201 0.0838333
R14836 VSSD.n231 VSSD.n227 0.0838333
R14837 VSSD.n656 VSSD.n580 0.0838333
R14838 VSSD.n605 VSSD.n604 0.0838333
R14839 VSSD.n730 VSSD.n729 0.0838333
R14840 VSSD.n3698 VSSD.n30 0.0838333
R14841 VSSD.n314 VSSD 0.082648
R14842 VSSD.n553 VSSD 0.082648
R14843 VSSD.n3203 VSSD.n1049 0.0812292
R14844 VSSD.n3141 VSSD.n1061 0.0812292
R14845 VSSD.n1358 VSSD.n1357 0.0812292
R14846 VSSD.n2354 VSSD.n1426 0.0812292
R14847 VSSD.n2252 VSSD.n2126 0.0812292
R14848 VSSD.n1683 VSSD.n1682 0.0812292
R14849 VSSD.n3569 VSSD.n55 0.0812292
R14850 VSSD.n3707 VSSD.n3706 0.0812292
R14851 VSSD.n1356 VSSD.n1054 0.0792941
R14852 VSSD.n2849 VSSD.n2848 0.0792941
R14853 VSSD.n2626 VSSD.n1104 0.0792941
R14854 VSSD.n2852 VSSD.n1311 0.0792941
R14855 VSSD.n853 VSSD.n851 0.0760208
R14856 VSSD.n3145 VSSD.n1058 0.0760208
R14857 VSSD.n2345 VSSD.n2311 0.0760208
R14858 VSSD.n2125 VSSD.n2123 0.0760208
R14859 VSSD.n1802 VSSD.n1801 0.0760208
R14860 VSSD.n3560 VSSD.n64 0.0760208
R14861 VSSD.n341 VSSD.n340 0.0760208
R14862 VSSD.n3697 VSSD.n33 0.0760208
R14863 VSSD.n3150 VSSD.n1054 0.0721059
R14864 VSSD.n2849 VSSD.n1015 0.0721059
R14865 VSSD.n2946 VSSD.n1104 0.0721059
R14866 VSSD.n2889 VSSD.n2852 0.0721059
R14867 VSSD.n1167 VSSD.n1136 0.0708125
R14868 VSSD.n3322 VSSD.n1019 0.0708125
R14869 VSSD.n2881 VSSD.n2858 0.0708125
R14870 VSSD.n2997 VSSD.n1087 0.0708125
R14871 VSSD.n2574 VSSD.n2573 0.0708125
R14872 VSSD.n2838 VSSD.n1319 0.0708125
R14873 VSSD.n1559 VSSD.n1478 0.0708125
R14874 VSSD.n1960 VSSD.n1959 0.0708125
R14875 VSSD.n2290 VSSD.n1437 0.0708125
R14876 VSSD.n1944 VSSD.n1574 0.0708125
R14877 VSSD.n1648 VSSD.n1647 0.0708125
R14878 VSSD.n3427 VSSD.n121 0.0708125
R14879 VSSD.n3509 VSSD.n78 0.0708125
R14880 VSSD.n480 VSSD.n144 0.0708125
R14881 VSSD.n207 VSSD.n206 0.0708125
R14882 VSSD.n662 VSSD.n571 0.0708125
R14883 VSSD.n724 VSSD.n542 0.0708125
R14884 VSSD.n3016 VSSD.n1079 0.0700652
R14885 VSSD.n3674 VSSD.n3673 0.0685851
R14886 VSSD.n661 VSSD.n572 0.0680676
R14887 VSSD.n661 VSSD.n660 0.0680676
R14888 VSSD.n613 VSSD.n601 0.0680676
R14889 VSSD.n602 VSSD.n601 0.0680676
R14890 VSSD.n430 VSSD.n168 0.0680676
R14891 VSSD.n169 VSSD.n168 0.0680676
R14892 VSSD.n728 VSSD.n540 0.0680676
R14893 VSSD.n728 VSSD.n727 0.0680676
R14894 VSSD.n384 VSSD.n203 0.0680676
R14895 VSSD.n204 VSSD.n203 0.0680676
R14896 VSSD.n32 VSSD.n31 0.0680676
R14897 VSSD.n32 VSSD.n25 0.0680676
R14898 VSSD.n1007 VSSD.n738 0.0680676
R14899 VSSD.n1007 VSSD.n1006 0.0680676
R14900 VSSD.n756 VSSD.n755 0.0680676
R14901 VSSD.n756 VSSD.n754 0.0680676
R14902 VSSD.n3383 VSSD.n503 0.0680676
R14903 VSSD.n3383 VSSD.n3382 0.0680676
R14904 VSSD.n852 VSSD.n841 0.0680676
R14905 VSSD.n852 VSSD.n842 0.0680676
R14906 VSSD.n3326 VSSD.n1017 0.0680676
R14907 VSSD.n3326 VSSD.n3325 0.0680676
R14908 VSSD.n1222 VSSD.n1151 0.0680676
R14909 VSSD.n1223 VSSD.n1222 0.0680676
R14910 VSSD.n1169 VSSD.n1135 0.0680676
R14911 VSSD.n1171 VSSD.n1169 0.0680676
R14912 VSSD.n3187 VSSD.n3153 0.0680676
R14913 VSSD.n3187 VSSD.n3186 0.0680676
R14914 VSSD.n2999 VSSD.n1085 0.0680676
R14915 VSSD.n3000 VSSD.n2999 0.0680676
R14916 VSSD.n1110 VSSD.n1107 0.0680676
R14917 VSSD.n1110 VSSD.n1109 0.0680676
R14918 VSSD.n2857 VSSD.n2855 0.0680676
R14919 VSSD.n2857 VSSD.n2856 0.0680676
R14920 VSSD.n1062 VSSD.n1057 0.0680676
R14921 VSSD.n1064 VSSD.n1062 0.0680676
R14922 VSSD.n2842 VSSD.n1317 0.0680676
R14923 VSSD.n2842 VSSD.n2841 0.0680676
R14924 VSSD.n2534 VSSD.n2529 0.0680676
R14925 VSSD.n2534 VSSD.n2533 0.0680676
R14926 VSSD.n2575 VSSD.n2550 0.0680676
R14927 VSSD.n2576 VSSD.n2575 0.0680676
R14928 VSSD.n2800 VSSD.n1350 0.0680676
R14929 VSSD.n2800 VSSD.n2799 0.0680676
R14930 VSSD.n2472 VSSD.n1403 0.0680676
R14931 VSSD.n1404 VSSD.n1403 0.0680676
R14932 VSSD.n2511 VSSD.n1378 0.0680676
R14933 VSSD.n2513 VSSD.n2511 0.0680676
R14934 VSSD.n1553 VSSD.n1477 0.0680676
R14935 VSSD.n1555 VSSD.n1553 0.0680676
R14936 VSSD.n2310 VSSD.n2307 0.0680676
R14937 VSSD.n2310 VSSD.n2309 0.0680676
R14938 VSSD.n2294 VSSD.n1435 0.0680676
R14939 VSSD.n2294 VSSD.n2293 0.0680676
R14940 VSSD.n2035 VSSD.n2030 0.0680676
R14941 VSSD.n2035 VSSD.n2034 0.0680676
R14942 VSSD.n1958 VSSD.n1956 0.0680676
R14943 VSSD.n1958 VSSD.n1957 0.0680676
R14944 VSSD.n2241 VSSD.n2240 0.0680676
R14945 VSSD.n2240 VSSD.n2127 0.0680676
R14946 VSSD.n1851 VSSD.n1641 0.0680676
R14947 VSSD.n1642 VSSD.n1641 0.0680676
R14948 VSSD.n1896 VSSD.n1595 0.0680676
R14949 VSSD.n1596 VSSD.n1595 0.0680676
R14950 VSSD.n1938 VSSD.n1573 0.0680676
R14951 VSSD.n1940 VSSD.n1938 0.0680676
R14952 VSSD.n1800 VSSD.n1675 0.0680676
R14953 VSSD.n1800 VSSD.n1799 0.0680676
R14954 VSSD.n339 VSSD.n229 0.0680676
R14955 VSSD.n339 VSSD.n338 0.0680676
R14956 VSSD.n3511 VSSD.n84 0.0680676
R14957 VSSD.n3511 VSSD.n3510 0.0680676
R14958 VSSD.n107 VSSD.n102 0.0680676
R14959 VSSD.n107 VSSD.n106 0.0680676
R14960 VSSD.n129 VSSD.n128 0.0680676
R14961 VSSD.n128 VSSD.n123 0.0680676
R14962 VSSD.n63 VSSD.n61 0.0680676
R14963 VSSD.n63 VSSD.n62 0.0680676
R14964 VSSD.n479 VSSD.n145 0.0680676
R14965 VSSD.n479 VSSD.n478 0.0680676
R14966 VSSD.n760 VSSD.n759 0.0656042
R14967 VSSD.n1218 VSSD.n1152 0.0656042
R14968 VSSD.n2942 VSSD.n2941 0.0656042
R14969 VSSD.n2622 VSSD.n2621 0.0656042
R14970 VSSD.n2522 VSSD.n2521 0.0656042
R14971 VSSD.n2038 VSSD.n2037 0.0656042
R14972 VSSD.n3464 VSSD.n3463 0.0656042
R14973 VSSD.n432 VSSD.n166 0.0656042
R14974 VSSD.n615 VSSD.n599 0.0656042
R14975 VSSD.n2570 VSSD.n2557 0.0631167
R14976 VSSD.n667 VSSD.n566 0.0631167
R14977 VSSD.n497 VSSD 0.0603958
R14978 VSSD.n498 VSSD 0.0603958
R14979 VSSD.n513 VSSD 0.0603958
R14980 VSSD.n3373 VSSD 0.0603958
R14981 VSSD VSSD.n823 0.0603958
R14982 VSSD VSSD.n807 0.0603958
R14983 VSSD VSSD.n798 0.0603958
R14984 VSSD.n791 VSSD.n737 0.0603958
R14985 VSSD.n739 VSSD.n737 0.0603958
R14986 VSSD.n998 VSSD 0.0603958
R14987 VSSD.n997 VSSD 0.0603958
R14988 VSSD VSSD.n996 0.0603958
R14989 VSSD.n986 VSSD 0.0603958
R14990 VSSD VSSD.n985 0.0603958
R14991 VSSD.n978 VSSD 0.0603958
R14992 VSSD VSSD.n844 0.0603958
R14993 VSSD VSSD.n957 0.0603958
R14994 VSSD VSSD.n862 0.0603958
R14995 VSSD.n939 VSSD 0.0603958
R14996 VSSD.n868 VSSD 0.0603958
R14997 VSSD VSSD.n903 0.0603958
R14998 VSSD.n1145 VSSD 0.0603958
R14999 VSSD.n1146 VSSD 0.0603958
R15000 VSSD.n1300 VSSD 0.0603958
R15001 VSSD.n1301 VSSD 0.0603958
R15002 VSSD VSSD.n1154 0.0603958
R15003 VSSD.n1208 VSSD 0.0603958
R15004 VSSD VSSD.n1291 0.0603958
R15005 VSSD.n1267 VSSD 0.0603958
R15006 VSSD.n1253 VSSD 0.0603958
R15007 VSSD.n1018 VSSD 0.0603958
R15008 VSSD.n1036 VSSD 0.0603958
R15009 VSSD.n3161 VSSD 0.0603958
R15010 VSSD.n3166 VSSD 0.0603958
R15011 VSSD VSSD.n3166 0.0603958
R15012 VSSD.n3167 VSSD 0.0603958
R15013 VSSD VSSD.n3159 0.0603958
R15014 VSSD.n3182 VSSD 0.0603958
R15015 VSSD VSSD.n1045 0.0603958
R15016 VSSD.n3211 VSSD 0.0603958
R15017 VSSD.n3214 VSSD 0.0603958
R15018 VSSD.n3215 VSSD 0.0603958
R15019 VSSD.n3216 VSSD 0.0603958
R15020 VSSD VSSD.n1038 0.0603958
R15021 VSSD VSSD.n1037 0.0603958
R15022 VSSD.n3299 VSSD 0.0603958
R15023 VSSD.n3263 VSSD 0.0603958
R15024 VSSD VSSD.n3262 0.0603958
R15025 VSSD.n2867 VSSD 0.0603958
R15026 VSSD.n2868 VSSD 0.0603958
R15027 VSSD VSSD.n2860 0.0603958
R15028 VSSD.n2877 VSSD 0.0603958
R15029 VSSD.n2894 VSSD 0.0603958
R15030 VSSD.n2907 VSSD 0.0603958
R15031 VSSD.n2955 VSSD 0.0603958
R15032 VSSD.n2957 VSSD 0.0603958
R15033 VSSD VSSD.n2964 0.0603958
R15034 VSSD.n2965 VSSD 0.0603958
R15035 VSSD.n2992 VSSD.n2988 0.0603958
R15036 VSSD.n2993 VSSD.n2992 0.0603958
R15037 VSSD.n3006 VSSD 0.0603958
R15038 VSSD.n3010 VSSD 0.0603958
R15039 VSSD.n3021 VSSD 0.0603958
R15040 VSSD.n3053 VSSD 0.0603958
R15041 VSSD VSSD.n3052 0.0603958
R15042 VSSD VSSD.n3051 0.0603958
R15043 VSSD.n3027 VSSD 0.0603958
R15044 VSSD.n3029 VSSD 0.0603958
R15045 VSSD VSSD.n1076 0.0603958
R15046 VSSD.n3115 VSSD 0.0603958
R15047 VSSD VSSD.n3113 0.0603958
R15048 VSSD VSSD.n3076 0.0603958
R15049 VSSD.n2564 VSSD 0.0603958
R15050 VSSD.n2565 VSSD 0.0603958
R15051 VSSD.n2569 VSSD 0.0603958
R15052 VSSD.n2584 VSSD 0.0603958
R15053 VSSD.n2689 VSSD 0.0603958
R15054 VSSD.n2683 VSSD 0.0603958
R15055 VSSD.n2665 VSSD 0.0603958
R15056 VSSD VSSD.n2664 0.0603958
R15057 VSSD.n2650 VSSD.n1316 0.0603958
R15058 VSSD.n1318 VSSD.n1316 0.0603958
R15059 VSSD.n2833 VSSD 0.0603958
R15060 VSSD.n2830 VSSD 0.0603958
R15061 VSSD VSSD.n2822 0.0603958
R15062 VSSD VSSD.n2821 0.0603958
R15063 VSSD.n2815 VSSD 0.0603958
R15064 VSSD.n2788 VSSD 0.0603958
R15065 VSSD.n2774 VSSD 0.0603958
R15066 VSSD VSSD.n2773 0.0603958
R15067 VSSD.n2769 VSSD 0.0603958
R15068 VSSD VSSD.n2768 0.0603958
R15069 VSSD.n2728 VSSD 0.0603958
R15070 VSSD VSSD.n2727 0.0603958
R15071 VSSD.n1487 VSSD 0.0603958
R15072 VSSD.n1488 VSSD 0.0603958
R15073 VSSD.n1493 VSSD 0.0603958
R15074 VSSD.n1526 VSSD 0.0603958
R15075 VSSD.n1522 VSSD 0.0603958
R15076 VSSD VSSD.n2509 0.0603958
R15077 VSSD.n2506 VSSD 0.0603958
R15078 VSSD VSSD.n2497 0.0603958
R15079 VSSD.n2493 VSSD 0.0603958
R15080 VSSD.n2479 VSSD.n1397 0.0603958
R15081 VSSD.n2475 VSSD.n1397 0.0603958
R15082 VSSD VSSD.n2465 0.0603958
R15083 VSSD VSSD.n2457 0.0603958
R15084 VSSD.n2318 VSSD 0.0603958
R15085 VSSD.n2319 VSSD 0.0603958
R15086 VSSD.n2323 VSSD 0.0603958
R15087 VSSD.n2332 VSSD 0.0603958
R15088 VSSD VSSD.n2369 0.0603958
R15089 VSSD.n2370 VSSD 0.0603958
R15090 VSSD.n2373 VSSD 0.0603958
R15091 VSSD.n2382 VSSD 0.0603958
R15092 VSSD.n2383 VSSD 0.0603958
R15093 VSSD.n2451 VSSD 0.0603958
R15094 VSSD VSSD.n2450 0.0603958
R15095 VSSD VSSD.n2398 0.0603958
R15096 VSSD.n2416 VSSD 0.0603958
R15097 VSSD.n1968 VSSD 0.0603958
R15098 VSSD.n1972 VSSD 0.0603958
R15099 VSSD.n1973 VSSD 0.0603958
R15100 VSSD.n1977 VSSD 0.0603958
R15101 VSSD.n2019 VSSD 0.0603958
R15102 VSSD.n2020 VSSD 0.0603958
R15103 VSSD VSSD.n1456 0.0603958
R15104 VSSD.n2102 VSSD 0.0603958
R15105 VSSD.n2076 VSSD 0.0603958
R15106 VSSD VSSD.n2075 0.0603958
R15107 VSSD.n2067 VSSD.n1434 0.0603958
R15108 VSSD.n1436 VSSD.n1434 0.0603958
R15109 VSSD.n2285 VSSD 0.0603958
R15110 VSSD VSSD.n2278 0.0603958
R15111 VSSD.n2275 VSSD 0.0603958
R15112 VSSD VSSD.n2260 0.0603958
R15113 VSSD VSSD.n2128 0.0603958
R15114 VSSD.n2234 VSSD 0.0603958
R15115 VSSD VSSD.n2232 0.0603958
R15116 VSSD.n2214 VSSD 0.0603958
R15117 VSSD VSSD.n2213 0.0603958
R15118 VSSD VSSD.n2143 0.0603958
R15119 VSSD.n2209 VSSD 0.0603958
R15120 VSSD VSSD.n2160 0.0603958
R15121 VSSD.n2175 VSSD 0.0603958
R15122 VSSD.n2174 VSSD 0.0603958
R15123 VSSD.n2171 VSSD 0.0603958
R15124 VSSD.n1604 VSSD 0.0603958
R15125 VSSD.n1614 VSSD 0.0603958
R15126 VSSD VSSD.n1613 0.0603958
R15127 VSSD.n1907 VSSD 0.0603958
R15128 VSSD.n1620 VSSD 0.0603958
R15129 VSSD.n1886 VSSD 0.0603958
R15130 VSSD VSSD.n1884 0.0603958
R15131 VSSD.n1854 VSSD 0.0603958
R15132 VSSD.n1839 VSSD 0.0603958
R15133 VSSD.n1831 VSSD 0.0603958
R15134 VSSD VSSD.n1830 0.0603958
R15135 VSSD.n1827 VSSD 0.0603958
R15136 VSSD VSSD.n1826 0.0603958
R15137 VSSD.n1814 VSSD 0.0603958
R15138 VSSD VSSD.n1779 0.0603958
R15139 VSSD VSSD.n1778 0.0603958
R15140 VSSD.n1771 VSSD 0.0603958
R15141 VSSD.n1768 VSSD 0.0603958
R15142 VSSD VSSD.n1767 0.0603958
R15143 VSSD.n1698 VSSD 0.0603958
R15144 VSSD.n1727 VSSD 0.0603958
R15145 VSSD VSSD.n1726 0.0603958
R15146 VSSD VSSD.n3405 0.0603958
R15147 VSSD.n3406 VSSD 0.0603958
R15148 VSSD.n3407 VSSD 0.0603958
R15149 VSSD VSSD.n131 0.0603958
R15150 VSSD VSSD.n94 0.0603958
R15151 VSSD.n3482 VSSD 0.0603958
R15152 VSSD.n3505 VSSD.n83 0.0603958
R15153 VSSD.n3508 VSSD.n83 0.0603958
R15154 VSSD VSSD.n71 0.0603958
R15155 VSSD.n3543 VSSD 0.0603958
R15156 VSSD.n3654 VSSD 0.0603958
R15157 VSSD VSSD.n3653 0.0603958
R15158 VSSD.n138 VSSD 0.0603958
R15159 VSSD.n139 VSSD 0.0603958
R15160 VSSD.n486 VSSD 0.0603958
R15161 VSSD VSSD.n442 0.0603958
R15162 VSSD VSSD.n441 0.0603958
R15163 VSSD.n437 VSSD 0.0603958
R15164 VSSD.n182 VSSD 0.0603958
R15165 VSSD VSSD.n415 0.0603958
R15166 VSSD.n390 VSSD.n197 0.0603958
R15167 VSSD.n387 VSSD.n197 0.0603958
R15168 VSSD VSSD.n377 0.0603958
R15169 VSSD VSSD.n211 0.0603958
R15170 VSSD.n373 VSSD 0.0603958
R15171 VSSD VSSD.n364 0.0603958
R15172 VSSD VSSD.n363 0.0603958
R15173 VSSD.n237 VSSD 0.0603958
R15174 VSSD VSSD.n333 0.0603958
R15175 VSSD VSSD.n243 0.0603958
R15176 VSSD.n321 VSSD 0.0603958
R15177 VSSD.n250 VSSD 0.0603958
R15178 VSSD.n309 VSSD 0.0603958
R15179 VSSD.n565 VSSD 0.0603958
R15180 VSSD.n669 VSSD 0.0603958
R15181 VSSD VSSD.n668 0.0603958
R15182 VSSD.n644 VSSD 0.0603958
R15183 VSSD.n703 VSSD.n539 0.0603958
R15184 VSSD.n541 VSSD.n539 0.0603958
R15185 VSSD VSSD.n713 0.0603958
R15186 VSSD VSSD.n45 0.0603958
R15187 VSSD.n3671 VSSD 0.0603958
R15188 VSSD.n3672 VSSD 0.0603958
R15189 VSSD VSSD.n38 0.0603958
R15190 VSSD VSSD.n3721 0.0603958
R15191 VSSD.n3722 VSSD 0.0603958
R15192 VSSD.n3733 VSSD 0.0603958
R15193 VSSD.n3734 VSSD 0.0603958
R15194 VSSD.n3735 VSSD 0.0603958
R15195 VSSD.n3739 VSSD 0.0603958
R15196 VSSD VSSD.n6 0.0603958
R15197 VSSD.n3774 VSSD 0.0603958
R15198 VSSD.n3202 VSSD 0.0577917
R15199 VSSD.n659 VSSD.n574 0.0574697
R15200 VSSD.n612 VSSD.n610 0.0574697
R15201 VSSD.n429 VSSD.n427 0.0574697
R15202 VSSD.n726 VSSD.n538 0.0574697
R15203 VSSD.n383 VSSD.n381 0.0574697
R15204 VSSD.n29 VSSD.n26 0.0574697
R15205 VSSD.n1005 VSSD.n736 0.0574697
R15206 VSSD.n753 VSSD.n530 0.0574697
R15207 VSSD.n3381 VSSD.n505 0.0574697
R15208 VSSD.n962 VSSD.n961 0.0574697
R15209 VSSD.n3324 VSSD.n1016 0.0574697
R15210 VSSD.n1224 VSSD.n1150 0.0574697
R15211 VSSD.n1170 VSSD.n1133 0.0574697
R15212 VSSD.n3151 VSSD.n1051 0.0574697
R15213 VSSD.n3001 VSSD.n1084 0.0574697
R15214 VSSD.n1105 VSSD.n1103 0.0574697
R15215 VSSD.n2853 VSSD.n1131 0.0574697
R15216 VSSD.n1063 VSSD.n1055 0.0574697
R15217 VSSD.n2840 VSSD.n1315 0.0574697
R15218 VSSD.n2527 VSSD.n1373 0.0574697
R15219 VSSD.n2577 VSSD.n2549 0.0574697
R15220 VSSD.n2798 VSSD.n1352 0.0574697
R15221 VSSD.n2471 VSSD.n2469 0.0574697
R15222 VSSD.n2512 VSSD.n1376 0.0574697
R15223 VSSD.n1554 VSSD.n1475 0.0574697
R15224 VSSD.n2305 VSSD.n1428 0.0574697
R15225 VSSD.n2292 VSSD.n1433 0.0574697
R15226 VSSD.n1455 VSSD.n1453 0.0574697
R15227 VSSD.n1954 VSSD.n1473 0.0574697
R15228 VSSD.n2248 VSSD.n2247 0.0574697
R15229 VSSD.n1850 VSSD.n1848 0.0574697
R15230 VSSD.n1895 VSSD.n1893 0.0574697
R15231 VSSD.n1939 VSSD.n1571 0.0574697
R15232 VSSD.n1798 VSSD.n1677 0.0574697
R15233 VSSD.n337 VSSD.n235 0.0574697
R15234 VSSD.n82 VSSD.n80 0.0574697
R15235 VSSD.n100 VSSD.n98 0.0574697
R15236 VSSD.n126 VSSD.n124 0.0574697
R15237 VSSD.n59 VSSD.n57 0.0574697
R15238 VSSD.n150 VSSD.n149 0.0574697
R15239 VSSD.n477 VSSD.n476 0.0574697
R15240 VSSD.n759 VSSD.n528 0.0551875
R15241 VSSD.n824 VSSD.n767 0.0551875
R15242 VSSD.n1213 VSSD.n1152 0.0551875
R15243 VSSD.n1293 VSSD.n1227 0.0551875
R15244 VSSD.n2942 VSSD.n1108 0.0551875
R15245 VSSD.n2950 VSSD.n2949 0.0551875
R15246 VSSD.n2622 VSSD.n2530 0.0551875
R15247 VSSD.n2630 VSSD.n2629 0.0551875
R15248 VSSD.n2522 VSSD.n1379 0.0551875
R15249 VSSD.n2516 VSSD.n2510 0.0551875
R15250 VSSD.n2038 VSSD.n2031 0.0551875
R15251 VSSD.n2046 VSSD.n2045 0.0551875
R15252 VSSD.n1890 VSSD.n1889 0.0551875
R15253 VSSD.n3464 VSSD.n103 0.0551875
R15254 VSSD.n3472 VSSD.n3471 0.0551875
R15255 VSSD.n433 VSSD.n432 0.0551875
R15256 VSSD.n424 VSSD.n423 0.0551875
R15257 VSSD.n616 VSSD.n615 0.0551875
R15258 VSSD.n607 VSSD.n558 0.0551875
R15259 VSSD.n3199 VSSD.n1052 0.0549647
R15260 VSSD.n3333 VSSD.n3332 0.0549647
R15261 VSSD.n3336 VSSD.n533 0.0549647
R15262 VSSD.n1310 VSSD.n534 0.0549647
R15263 VSSD.n3188 VSSD 0.0538854
R15264 VSSD.n3195 VSSD 0.0525833
R15265 VSSD.n1348 VSSD 0.0525833
R15266 VSSD.n1003 VSSD.n1002 0.0499792
R15267 VSSD.n1305 VSSD.n1136 0.0499792
R15268 VSSD.n3322 VSSD.n3321 0.0499792
R15269 VSSD.n2884 VSSD.n2858 0.0499792
R15270 VSSD.n1087 VSSD.n1082 0.0499792
R15271 VSSD.n2574 VSSD.n2551 0.0499792
R15272 VSSD.n2838 VSSD.n2837 0.0499792
R15273 VSSD.n1563 VSSD.n1478 0.0499792
R15274 VSSD.n1410 VSSD.n1409 0.0499792
R15275 VSSD.n1981 VSSD.n1959 0.0499792
R15276 VSSD.n2290 VSSD.n2289 0.0499792
R15277 VSSD.n1948 VSSD.n1574 0.0499792
R15278 VSSD.n1647 VSSD.n1644 0.0499792
R15279 VSSD.n3417 VSSD.n121 0.0499792
R15280 VSSD.n3521 VSSD.n78 0.0499792
R15281 VSSD.n481 VSSD.n480 0.0499792
R15282 VSSD.n208 VSSD.n207 0.0499792
R15283 VSSD.n663 VSSD.n662 0.0499792
R15284 VSSD.n724 VSSD.n723 0.0499792
R15285 VSSD.n2350 VSSD.n2304 0.0477765
R15286 VSSD.n2301 VSSD.n1314 0.0477765
R15287 VSSD.n2526 VSSD.n1375 0.0477765
R15288 VSSD.n1569 VSSD.n1568 0.0477765
R15289 VSSD VSSD.n3327 0.047375
R15290 VSSD.n1646 VSSD 0.047375
R15291 VSSD.n855 VSSD.n853 0.0447708
R15292 VSSD.n3189 VSSD.n3188 0.0447708
R15293 VSSD.n3142 VSSD.n1058 0.0447708
R15294 VSSD.n2801 VSSD.n1349 0.0447708
R15295 VSSD.n2311 VSSD.n2308 0.0447708
R15296 VSSD.n2253 VSSD.n2125 0.0447708
R15297 VSSD.n1801 VSSD.n1674 0.0447708
R15298 VSSD.n3557 VSSD.n64 0.0447708
R15299 VSSD.n340 VSSD.n228 0.0447708
R15300 VSSD.n33 VSSD.n24 0.0447708
R15301 VSSD.n785 VSSD.n784 0.0443356
R15302 VSSD.n1890 VSSD 0.0434688
R15303 VSSD.n3471 VSSD 0.0434688
R15304 VSSD.n607 VSSD 0.0434688
R15305 VSSD VSSD.n2532 0.0421667
R15306 VSSD.n576 VSSD.n572 0.0410405
R15307 VSSD.n660 VSSD.n573 0.0410405
R15308 VSSD.n614 VSSD.n613 0.0410405
R15309 VSSD.n603 VSSD.n602 0.0410405
R15310 VSSD.n431 VSSD.n430 0.0410405
R15311 VSSD.n170 VSSD.n169 0.0410405
R15312 VSSD.n731 VSSD.n540 0.0410405
R15313 VSSD.n727 VSSD.n725 0.0410405
R15314 VSSD.n385 VSSD.n384 0.0410405
R15315 VSSD.n205 VSSD.n204 0.0410405
R15316 VSSD.n3699 VSSD.n31 0.0410405
R15317 VSSD.n3705 VSSD.n25 0.0410405
R15318 VSSD.n1010 VSSD.n738 0.0410405
R15319 VSSD.n1006 VSSD.n1004 0.0410405
R15320 VSSD.n755 VSSD.n529 0.0410405
R15321 VSSD.n765 VSSD.n754 0.0410405
R15322 VSSD.n507 VSSD.n503 0.0410405
R15323 VSSD.n3382 VSSD.n504 0.0410405
R15324 VSSD.n841 VSSD.n840 0.0410405
R15325 VSSD.n843 VSSD.n842 0.0410405
R15326 VSSD.n3329 VSSD.n1017 0.0410405
R15327 VSSD.n3325 VSSD.n3323 0.0410405
R15328 VSSD.n1209 VSSD.n1151 0.0410405
R15329 VSSD.n1223 VSSD.n1149 0.0410405
R15330 VSSD.n1307 VSSD.n1135 0.0410405
R15331 VSSD.n1172 VSSD.n1171 0.0410405
R15332 VSSD.n3196 VSSD.n3153 0.0410405
R15333 VSSD.n3186 VSSD.n1050 0.0410405
R15334 VSSD.n2989 VSSD.n1085 0.0410405
R15335 VSSD.n3000 VSSD.n1083 0.0410405
R15336 VSSD.n2943 VSSD.n1107 0.0410405
R15337 VSSD.n1109 VSSD.n1102 0.0410405
R15338 VSSD.n2886 VSSD.n2855 0.0410405
R15339 VSSD.n2856 VSSD.n1130 0.0410405
R15340 VSSD.n3147 VSSD.n1057 0.0410405
R15341 VSSD.n3140 VSSD.n1064 0.0410405
R15342 VSSD.n2845 VSSD.n1317 0.0410405
R15343 VSSD.n2841 VSSD.n2839 0.0410405
R15344 VSSD.n2623 VSSD.n2529 0.0410405
R15345 VSSD.n2533 VSSD.n1372 0.0410405
R15346 VSSD.n2554 VSSD.n2550 0.0410405
R15347 VSSD.n2576 VSSD.n2548 0.0410405
R15348 VSSD.n1353 VSSD.n1350 0.0410405
R15349 VSSD.n2799 VSSD.n1351 0.0410405
R15350 VSSD.n2473 VSSD.n2472 0.0410405
R15351 VSSD.n1405 VSSD.n1404 0.0410405
R15352 VSSD.n2523 VSSD.n1378 0.0410405
R15353 VSSD.n2514 VSSD.n2513 0.0410405
R15354 VSSD.n1565 VSSD.n1477 0.0410405
R15355 VSSD.n1557 VSSD.n1555 0.0410405
R15356 VSSD.n2347 VSSD.n2307 0.0410405
R15357 VSSD.n2309 VSSD.n1427 0.0410405
R15358 VSSD.n2297 VSSD.n1435 0.0410405
R15359 VSSD.n2293 VSSD.n2291 0.0410405
R15360 VSSD.n2039 VSSD.n2030 0.0410405
R15361 VSSD.n2034 VSSD.n1452 0.0410405
R15362 VSSD.n1983 VSSD.n1956 0.0410405
R15363 VSSD.n1957 VSSD.n1472 0.0410405
R15364 VSSD.n2244 VSSD.n2241 0.0410405
R15365 VSSD.n2251 VSSD.n2127 0.0410405
R15366 VSSD.n1852 VSSD.n1851 0.0410405
R15367 VSSD.n1643 VSSD.n1642 0.0410405
R15368 VSSD.n1897 VSSD.n1896 0.0410405
R15369 VSSD.n1597 VSSD.n1596 0.0410405
R15370 VSSD.n1950 VSSD.n1573 0.0410405
R15371 VSSD.n1942 VSSD.n1940 0.0410405
R15372 VSSD.n1678 VSSD.n1675 0.0410405
R15373 VSSD.n1799 VSSD.n1676 0.0410405
R15374 VSSD.n232 VSSD.n229 0.0410405
R15375 VSSD.n338 VSSD.n230 0.0410405
R15376 VSSD.n3514 VSSD.n84 0.0410405
R15377 VSSD.n3510 VSSD.n79 0.0410405
R15378 VSSD.n3465 VSSD.n102 0.0410405
R15379 VSSD.n106 VSSD.n97 0.0410405
R15380 VSSD.n3419 VSSD.n129 0.0410405
R15381 VSSD.n3425 VSSD.n123 0.0410405
R15382 VSSD.n3562 VSSD.n61 0.0410405
R15383 VSSD.n62 VSSD.n56 0.0410405
R15384 VSSD.n147 VSSD.n145 0.0410405
R15385 VSSD.n478 VSSD.n146 0.0410405
R15386 VSSD.n3189 VSSD.n1049 0.0395625
R15387 VSSD.n3142 VSSD.n3141 0.0395625
R15388 VSSD.n1357 VSSD.n1349 0.0395625
R15389 VSSD.n2308 VSSD.n1426 0.0395625
R15390 VSSD.n2253 VSSD.n2252 0.0395625
R15391 VSSD.n1682 VSSD.n1674 0.0395625
R15392 VSSD.n3557 VSSD.n55 0.0395625
R15393 VSSD.n236 VSSD.n228 0.0395625
R15394 VSSD.n3706 VSSD.n24 0.0395625
R15395 VSSD.n2580 VSSD 0.0369583
R15396 VSSD.n3385 VSSD.n502 0.0343542
R15397 VSSD.n1306 VSSD.n1305 0.0343542
R15398 VSSD.n3321 VSSD.n1021 0.0343542
R15399 VSSD.n3162 VSSD 0.0343542
R15400 VSSD VSSD.n2876 0.0343542
R15401 VSSD.n2885 VSSD.n2884 0.0343542
R15402 VSSD VSSD.n2956 0.0343542
R15403 VSSD.n3004 VSSD.n1082 0.0343542
R15404 VSSD.n2553 VSSD.n2551 0.0343542
R15405 VSSD.n2837 VSSD.n1321 0.0343542
R15406 VSSD VSSD.n1370 0.0343542
R15407 VSSD.n1564 VSSD.n1563 0.0343542
R15408 VSSD.n2496 VSSD 0.0343542
R15409 VSSD.n1982 VSSD.n1981 0.0343542
R15410 VSSD.n2233 VSSD 0.0343542
R15411 VSSD.n1949 VSSD.n1948 0.0343542
R15412 VSSD.n1885 VSSD 0.0343542
R15413 VSSD.n1845 VSSD.n1644 0.0343542
R15414 VSSD.n3418 VSSD.n3417 0.0343542
R15415 VSSD.n3521 VSSD.n3520 0.0343542
R15416 VSSD.n481 VSSD.n143 0.0343542
R15417 VSSD.n663 VSSD.n570 0.0343542
R15418 VSSD.n723 VSSD.n544 0.0343542
R15419 VSSD VSSD.n498 0.0330521
R15420 VSSD.n824 VSSD 0.0330521
R15421 VSSD.n986 VSSD 0.0330521
R15422 VSSD VSSD.n867 0.0330521
R15423 VSSD.n1146 VSSD 0.0330521
R15424 VSSD.n1293 VSSD 0.0330521
R15425 VSSD VSSD.n1036 0.0330521
R15426 VSSD.n1038 VSSD 0.0330521
R15427 VSSD.n2868 VSSD 0.0330521
R15428 VSSD.n2950 VSSD 0.0330521
R15429 VSSD.n3053 VSSD 0.0330521
R15430 VSSD.n3115 VSSD 0.0330521
R15431 VSSD.n2565 VSSD 0.0330521
R15432 VSSD VSSD.n2630 0.0330521
R15433 VSSD.n2822 VSSD 0.0330521
R15434 VSSD.n2769 VSSD 0.0330521
R15435 VSSD.n1488 VSSD 0.0330521
R15436 VSSD.n2510 VSSD 0.0330521
R15437 VSSD.n2457 VSSD 0.0330521
R15438 VSSD VSSD.n2383 0.0330521
R15439 VSSD VSSD.n1972 0.0330521
R15440 VSSD VSSD.n2046 0.0330521
R15441 VSSD.n2279 VSSD 0.0330521
R15442 VSSD.n2214 VSSD 0.0330521
R15443 VSSD.n1614 VSSD 0.0330521
R15444 VSSD VSSD.n1898 0.0330521
R15445 VSSD.n1889 VSSD 0.0330521
R15446 VSSD.n1830 VSSD 0.0330521
R15447 VSSD.n1768 VSSD 0.0330521
R15448 VSSD.n3407 VSSD 0.0330521
R15449 VSSD.n3472 VSSD 0.0330521
R15450 VSSD.n3533 VSSD 0.0330521
R15451 VSSD VSSD.n3591 0.0330521
R15452 VSSD VSSD.n139 0.0330521
R15453 VSSD.n423 VSSD 0.0330521
R15454 VSSD.n364 VSSD 0.0330521
R15455 VSSD.n312 VSSD 0.0330521
R15456 VSSD.n669 VSSD 0.0330521
R15457 VSSD.n558 VSSD 0.0330521
R15458 VSSD.n45 VSSD 0.0330521
R15459 VSSD VSSD.n3734 0.0330521
R15460 VSSD VSSD.n497 0.03175
R15461 VSSD VSSD.n1145 0.03175
R15462 VSSD.n1154 VSSD 0.03175
R15463 VSSD.n3167 VSSD 0.03175
R15464 VSSD VSSD.n3152 0.03175
R15465 VSSD VSSD.n3215 0.03175
R15466 VSSD VSSD.n2867 0.03175
R15467 VSSD.n3052 VSSD 0.03175
R15468 VSSD VSSD.n2564 0.03175
R15469 VSSD VSSD.n2569 0.03175
R15470 VSSD VSSD.n1346 0.03175
R15471 VSSD.n2802 VSSD 0.03175
R15472 VSSD VSSD.n1487 0.03175
R15473 VSSD.n2509 VSSD 0.03175
R15474 VSSD.n1410 VSSD 0.03175
R15475 VSSD.n2319 VSSD 0.03175
R15476 VSSD.n2370 VSSD 0.03175
R15477 VSSD.n2451 VSSD 0.03175
R15478 VSSD.n1968 VSSD 0.03175
R15479 VSSD.n1973 VSSD 0.03175
R15480 VSSD VSSD.n2019 0.03175
R15481 VSSD.n2076 VSSD 0.03175
R15482 VSSD.n2278 VSSD 0.03175
R15483 VSSD VSSD.n1604 0.03175
R15484 VSSD.n1827 VSSD 0.03175
R15485 VSSD.n1779 VSSD 0.03175
R15486 VSSD VSSD.n3406 0.03175
R15487 VSSD.n3654 VSSD 0.03175
R15488 VSSD VSSD.n138 0.03175
R15489 VSSD.n441 VSSD 0.03175
R15490 VSSD VSSD.n565 0.03175
R15491 VSSD.n668 VSSD 0.03175
R15492 VSSD VSSD.n3733 0.03175
R15493 VSSD.n3735 VSSD 0.03175
R15494 VSSD.n3564 VSSD.n59 0.0292489
R15495 VSSD.n3566 VSSD.n57 0.0292489
R15496 VSSD.n235 VSSD.n234 0.0292489
R15497 VSSD.n337 VSSD.n336 0.0292489
R15498 VSSD.n1680 VSSD.n1677 0.0292489
R15499 VSSD.n1798 VSSD.n1797 0.0292489
R15500 VSSD.n2247 VSSD.n2246 0.0292489
R15501 VSSD.n2249 VSSD.n2248 0.0292489
R15502 VSSD.n2349 VSSD.n2305 0.0292489
R15503 VSSD.n2351 VSSD.n1428 0.0292489
R15504 VSSD.n1355 VSSD.n1352 0.0292489
R15505 VSSD.n2798 VSSD.n2797 0.0292489
R15506 VSSD.n3149 VSSD.n1055 0.0292489
R15507 VSSD.n1063 VSSD.n1053 0.0292489
R15508 VSSD.n3198 VSSD.n3151 0.0292489
R15509 VSSD.n3200 VSSD.n1051 0.0292489
R15510 VSSD.n963 VSSD.n962 0.0292489
R15511 VSSD.n961 VSSD.n960 0.0292489
R15512 VSSD.n3701 VSSD.n29 0.0292489
R15513 VSSD.n3703 VSSD.n26 0.0292489
R15514 VSSD.n3516 VSSD.n82 0.0292489
R15515 VSSD.n3518 VSSD.n80 0.0292489
R15516 VSSD.n383 VSSD.n382 0.0292489
R15517 VSSD.n381 VSSD.n380 0.0292489
R15518 VSSD.n1850 VSSD.n1849 0.0292489
R15519 VSSD.n1848 VSSD.n1847 0.0292489
R15520 VSSD.n2299 VSSD.n1433 0.0292489
R15521 VSSD.n2292 VSSD.n1431 0.0292489
R15522 VSSD.n2471 VSSD.n2470 0.0292489
R15523 VSSD.n2469 VSSD.n2468 0.0292489
R15524 VSSD.n2847 VSSD.n1315 0.0292489
R15525 VSSD.n2840 VSSD.n1313 0.0292489
R15526 VSSD.n2990 VSSD.n1084 0.0292489
R15527 VSSD.n3002 VSSD.n3001 0.0292489
R15528 VSSD.n3331 VSSD.n1016 0.0292489
R15529 VSSD.n3324 VSSD.n1014 0.0292489
R15530 VSSD.n1012 VSSD.n736 0.0292489
R15531 VSSD.n1005 VSSD.n735 0.0292489
R15532 VSSD.n733 VSSD.n538 0.0292489
R15533 VSSD.n726 VSSD.n537 0.0292489
R15534 VSSD.n3467 VSSD.n100 0.0292489
R15535 VSSD.n3469 VSSD.n98 0.0292489
R15536 VSSD.n429 VSSD.n428 0.0292489
R15537 VSSD.n427 VSSD.n426 0.0292489
R15538 VSSD.n1895 VSSD.n1894 0.0292489
R15539 VSSD.n1893 VSSD.n1892 0.0292489
R15540 VSSD.n2041 VSSD.n1455 0.0292489
R15541 VSSD.n2043 VSSD.n1453 0.0292489
R15542 VSSD.n2525 VSSD.n1376 0.0292489
R15543 VSSD.n2512 VSSD.n1374 0.0292489
R15544 VSSD.n2625 VSSD.n2527 0.0292489
R15545 VSSD.n2627 VSSD.n1373 0.0292489
R15546 VSSD.n2945 VSSD.n1105 0.0292489
R15547 VSSD.n2947 VSSD.n1103 0.0292489
R15548 VSSD.n1210 VSSD.n1150 0.0292489
R15549 VSSD.n1225 VSSD.n1224 0.0292489
R15550 VSSD.n3338 VSSD.n530 0.0292489
R15551 VSSD.n753 VSSD.n532 0.0292489
R15552 VSSD.n612 VSSD.n611 0.0292489
R15553 VSSD.n610 VSSD.n609 0.0292489
R15554 VSSD.n3421 VSSD.n126 0.0292489
R15555 VSSD.n3423 VSSD.n124 0.0292489
R15556 VSSD.n1952 VSSD.n1571 0.0292489
R15557 VSSD.n1939 VSSD.n1570 0.0292489
R15558 VSSD.n1985 VSSD.n1954 0.0292489
R15559 VSSD.n1987 VSSD.n1473 0.0292489
R15560 VSSD.n1567 VSSD.n1475 0.0292489
R15561 VSSD.n1554 VSSD.n1474 0.0292489
R15562 VSSD.n2555 VSSD.n2549 0.0292489
R15563 VSSD.n2578 VSSD.n2577 0.0292489
R15564 VSSD.n2888 VSSD.n2853 0.0292489
R15565 VSSD.n2890 VSSD.n1131 0.0292489
R15566 VSSD.n1309 VSSD.n1133 0.0292489
R15567 VSSD.n1170 VSSD.n1132 0.0292489
R15568 VSSD.n509 VSSD.n505 0.0292489
R15569 VSSD.n3381 VSSD.n3380 0.0292489
R15570 VSSD.n578 VSSD.n574 0.0292489
R15571 VSSD.n659 VSSD.n658 0.0292489
R15572 VSSD.n477 VSSD.n151 0.0292489
R15573 VSSD.n151 VSSD.n150 0.0292489
R15574 VSSD.n3340 VSSD.n528 0.0291458
R15575 VSSD.n966 VSSD.n965 0.0291458
R15576 VSSD.n958 VSSD 0.0291458
R15577 VSSD.n1213 VSSD.n1212 0.0291458
R15578 VSSD.n1108 VSSD.n1106 0.0291458
R15579 VSSD.n3033 VSSD.n1056 0.0291458
R15580 VSSD.n2530 VSSD.n2528 0.0291458
R15581 VSSD.n2805 VSSD.n1346 0.0291458
R15582 VSSD.n1379 VSSD.n1377 0.0291458
R15583 VSSD.n2342 VSSD.n2306 0.0291458
R15584 VSSD.n2031 VSSD.n2029 0.0291458
R15585 VSSD.n2242 VSSD.n2119 0.0291458
R15586 VSSD.n1899 VSSD.n1593 0.0291458
R15587 VSSD.n1807 VSSD.n1671 0.0291458
R15588 VSSD.n103 VSSD.n101 0.0291458
R15589 VSSD.n3555 VSSD.n60 0.0291458
R15590 VSSD.n433 VSSD.n164 0.0291458
R15591 VSSD.n231 VSSD.n225 0.0291458
R15592 VSSD.n334 VSSD 0.0291458
R15593 VSSD.n616 VSSD.n598 0.0291458
R15594 VSSD.n3694 VSSD.n30 0.0291458
R15595 VSSD VSSD.n3384 0.0278438
R15596 VSSD VSSD.n744 0.0265417
R15597 VSSD.n2885 VSSD 0.0265417
R15598 VSSD.n2466 VSSD 0.0265417
R15599 VSSD VSSD.n1445 0.0265417
R15600 VSSD.n1949 VSSD 0.0265417
R15601 VSSD.n3418 VSSD 0.0265417
R15602 VSSD.n378 VSSD 0.0265417
R15603 VSSD.n570 VSSD 0.0265417
R15604 VSSD.n3378 VSSD.n3377 0.0239375
R15605 VSSD.n1009 VSSD.n739 0.0239375
R15606 VSSD.n1175 VSSD.n1174 0.0239375
R15607 VSSD.n1284 VSSD 0.0239375
R15608 VSSD.n3328 VSSD.n1018 0.0239375
R15609 VSSD.n2893 VSSD.n2892 0.0239375
R15610 VSSD VSSD.n2930 0.0239375
R15611 VSSD.n2993 VSSD.n1086 0.0239375
R15612 VSSD.n2581 VSSD.n2580 0.0239375
R15613 VSSD.n2844 VSSD.n1318 0.0239375
R15614 VSSD.n2821 VSSD 0.0239375
R15615 VSSD.n1552 VSSD.n1551 0.0239375
R15616 VSSD.n2475 VSSD.n2474 0.0239375
R15617 VSSD.n1990 VSSD.n1989 0.0239375
R15618 VSSD.n2296 VSSD.n1436 0.0239375
R15619 VSSD.n1937 VSSD.n1936 0.0239375
R15620 VSSD.n1854 VSSD.n1853 0.0239375
R15621 VSSD.n122 VSSD.n119 0.0239375
R15622 VSSD.n3513 VSSD.n3508 0.0239375
R15623 VSSD.n474 VSSD.n473 0.0239375
R15624 VSSD.n387 VSSD.n386 0.0239375
R15625 VSSD.n656 VSSD.n655 0.0239375
R15626 VSSD.n730 VSSD.n541 0.0239375
R15627 VSSD.n3385 VSSD 0.0226354
R15628 VSSD.n3377 VSSD 0.0226354
R15629 VSSD.n3357 VSSD 0.0226354
R15630 VSSD.n763 VSSD 0.0226354
R15631 VSSD.n808 VSSD 0.0226354
R15632 VSSD.n799 VSSD 0.0226354
R15633 VSSD VSSD.n740 0.0226354
R15634 VSSD.n1002 VSSD 0.0226354
R15635 VSSD.n990 VSSD 0.0226354
R15636 VSSD VSSD.n829 0.0226354
R15637 VSSD.n978 VSSD 0.0226354
R15638 VSSD.n855 VSSD 0.0226354
R15639 VSSD VSSD.n865 0.0226354
R15640 VSSD.n904 VSSD 0.0226354
R15641 VSSD.n897 VSSD 0.0226354
R15642 VSSD VSSD.n1300 0.0226354
R15643 VSSD.n1203 VSSD 0.0226354
R15644 VSSD.n1219 VSSD 0.0226354
R15645 VSSD.n1285 VSSD 0.0226354
R15646 VSSD.n1271 VSSD 0.0226354
R15647 VSSD.n1267 VSSD 0.0226354
R15648 VSSD.n3307 VSSD 0.0226354
R15649 VSSD VSSD.n3181 0.0226354
R15650 VSSD VSSD.n3182 0.0226354
R15651 VSSD.n3183 VSSD 0.0226354
R15652 VSSD.n3194 VSSD 0.0226354
R15653 VSSD VSSD.n3214 0.0226354
R15654 VSSD.n3223 VSSD 0.0226354
R15655 VSSD VSSD.n1037 0.0226354
R15656 VSSD.n3280 VSSD 0.0226354
R15657 VSSD.n3256 VSSD 0.0226354
R15658 VSSD VSSD.n2893 0.0226354
R15659 VSSD.n2904 VSSD 0.0226354
R15660 VSSD.n2926 VSSD 0.0226354
R15661 VSSD.n2937 VSSD 0.0226354
R15662 VSSD.n2957 VSSD 0.0226354
R15663 VSSD.n3011 VSSD 0.0226354
R15664 VSSD VSSD.n3021 0.0226354
R15665 VSSD VSSD.n3024 0.0226354
R15666 VSSD VSSD.n3027 0.0226354
R15667 VSSD VSSD.n3029 0.0226354
R15668 VSSD.n3113 VSSD 0.0226354
R15669 VSSD.n2581 VSSD 0.0226354
R15670 VSSD.n2531 VSSD 0.0226354
R15671 VSSD.n2689 VSSD 0.0226354
R15672 VSSD.n2687 VSSD 0.0226354
R15673 VSSD.n2683 VSSD 0.0226354
R15674 VSSD.n2823 VSSD 0.0226354
R15675 VSSD VSSD.n1334 0.0226354
R15676 VSSD.n2815 VSSD 0.0226354
R15677 VSSD VSSD.n1359 0.0226354
R15678 VSSD.n2768 VSSD 0.0226354
R15679 VSSD.n2745 VSSD 0.0226354
R15680 VSSD.n2721 VSSD 0.0226354
R15681 VSSD VSSD.n1510 0.0226354
R15682 VSSD.n1525 VSSD 0.0226354
R15683 VSSD.n2517 VSSD 0.0226354
R15684 VSSD.n2498 VSSD 0.0226354
R15685 VSSD.n2493 VSSD 0.0226354
R15686 VSSD VSSD.n1408 0.0226354
R15687 VSSD VSSD.n2318 0.0226354
R15688 VSSD VSSD.n2331 0.0226354
R15689 VSSD VSSD.n2332 0.0226354
R15690 VSSD VSSD.n2381 0.0226354
R15691 VSSD VSSD.n2382 0.0226354
R15692 VSSD.n2432 VSSD 0.0226354
R15693 VSSD.n2408 VSSD 0.0226354
R15694 VSSD VSSD.n2018 0.0226354
R15695 VSSD.n2020 VSSD 0.0226354
R15696 VSSD.n2032 VSSD 0.0226354
R15697 VSSD VSSD.n2065 0.0226354
R15698 VSSD.n2289 VSSD 0.0226354
R15699 VSSD.n2285 VSSD 0.0226354
R15700 VSSD VSSD.n1447 0.0226354
R15701 VSSD.n2261 VSSD 0.0226354
R15702 VSSD.n2260 VSSD 0.0226354
R15703 VSSD.n2217 VSSD 0.0226354
R15704 VSSD.n2213 VSSD 0.0226354
R15705 VSSD.n2209 VSSD 0.0226354
R15706 VSSD.n2170 VSSD 0.0226354
R15707 VSSD.n1921 VSSD 0.0226354
R15708 VSSD.n1910 VSSD 0.0226354
R15709 VSSD.n1899 VSSD 0.0226354
R15710 VSSD.n1623 VSSD 0.0226354
R15711 VSSD.n1857 VSSD 0.0226354
R15712 VSSD VSSD.n1645 0.0226354
R15713 VSSD.n1837 VSSD 0.0226354
R15714 VSSD.n1831 VSSD 0.0226354
R15715 VSSD.n1817 VSSD 0.0226354
R15716 VSSD.n1814 VSSD 0.0226354
R15717 VSSD.n1780 VSSD 0.0226354
R15718 VSSD.n1767 VSSD 0.0226354
R15719 VSSD.n1744 VSSD 0.0226354
R15720 VSSD.n1720 VSSD 0.0226354
R15721 VSSD.n3443 VSSD 0.0226354
R15722 VSSD.n104 VSSD 0.0226354
R15723 VSSD.n3479 VSSD 0.0226354
R15724 VSSD.n3499 VSSD 0.0226354
R15725 VSSD VSSD.n3532 0.0226354
R15726 VSSD.n3540 VSSD 0.0226354
R15727 VSSD VSSD.n3590 0.0226354
R15728 VSSD.n3636 VSSD 0.0226354
R15729 VSSD.n3616 VSSD 0.0226354
R15730 VSSD.n3608 VSSD 0.0226354
R15731 VSSD.n443 VSSD 0.0226354
R15732 VSSD.n442 VSSD 0.0226354
R15733 VSSD.n175 VSSD 0.0226354
R15734 VSSD.n416 VSSD 0.0226354
R15735 VSSD.n415 VSSD 0.0226354
R15736 VSSD.n208 VSSD 0.0226354
R15737 VSSD.n377 VSSD 0.0226354
R15738 VSSD.n365 VSSD 0.0226354
R15739 VSSD.n363 VSSD 0.0226354
R15740 VSSD VSSD.n250 0.0226354
R15741 VSSD.n292 VSSD 0.0226354
R15742 VSSD.n272 VSSD 0.0226354
R15743 VSSD.n647 VSSD 0.0226354
R15744 VSSD.n636 VSSD 0.0226354
R15745 VSSD.n625 VSSD 0.0226354
R15746 VSSD VSSD.n606 0.0226354
R15747 VSSD.n695 VSSD 0.0226354
R15748 VSSD.n713 VSSD 0.0226354
R15749 VSSD VSSD.n3671 0.0226354
R15750 VSSD.n3681 VSSD 0.0226354
R15751 VSSD.n3728 VSSD 0.0226354
R15752 VSSD VSSD.n3762 0.0226354
R15753 VSSD.n3763 VSSD 0.0226354
R15754 VSSD.n3771 VSSD 0.0226354
R15755 VSSD.n3786 VSSD 0.0226354
R15756 VSSD.n854 VSSD 0.0213333
R15757 VSSD VSSD.n236 0.0213333
R15758 VSSD VSSD.n2854 0.0200312
R15759 VSSD VSSD.n1572 0.0200312
R15760 VSSD VSSD.n127 0.0200312
R15761 VSSD.n3568 VSSD 0.0200312
R15762 VSSD VSSD.n566 0.0200312
R15763 VSSD.n760 VSSD.n757 0.0187292
R15764 VSSD.n764 VSSD.n763 0.0187292
R15765 VSSD.n1221 VSSD.n1218 0.0187292
R15766 VSSD.n1220 VSSD.n1219 0.0187292
R15767 VSSD.n2941 VSSD.n1111 0.0187292
R15768 VSSD.n2937 VSSD.n2936 0.0187292
R15769 VSSD.n2621 VSSD.n2535 0.0187292
R15770 VSSD.n2532 VSSD.n2531 0.0187292
R15771 VSSD.n2521 VSSD.n1380 0.0187292
R15772 VSSD.n2517 VSSD.n1383 0.0187292
R15773 VSSD.n2037 VSSD.n2036 0.0187292
R15774 VSSD.n2033 VSSD.n2032 0.0187292
R15775 VSSD.n1621 VSSD.n1620 0.0187292
R15776 VSSD.n1623 VSSD.n1622 0.0187292
R15777 VSSD.n3463 VSSD.n108 0.0187292
R15778 VSSD.n105 VSSD.n104 0.0187292
R15779 VSSD.n173 VSSD.n166 0.0187292
R15780 VSSD.n175 VSSD.n174 0.0187292
R15781 VSSD.n604 VSSD.n599 0.0187292
R15782 VSSD.n606 VSSD.n605 0.0187292
R15783 VSSD VSSD.n854 0.0174271
R15784 VSSD VSSD.n2801 0.016125
R15785 VSSD.n513 VSSD.n511 0.0135208
R15786 VSSD.n1008 VSSD.n740 0.0135208
R15787 VSSD.n1168 VSSD.n1167 0.0135208
R15788 VSSD.n3327 VSSD.n1019 0.0135208
R15789 VSSD.n2881 VSSD.n1129 0.0135208
R15790 VSSD.n2998 VSSD.n2997 0.0135208
R15791 VSSD.n2573 VSSD.n2552 0.0135208
R15792 VSSD.n2843 VSSD.n1319 0.0135208
R15793 VSSD.n1559 VSSD.n1558 0.0135208
R15794 VSSD.n1408 VSSD.n1401 0.0135208
R15795 VSSD.n1960 VSSD.n1471 0.0135208
R15796 VSSD.n2295 VSSD.n1437 0.0135208
R15797 VSSD.n1944 VSSD.n1943 0.0135208
R15798 VSSD.n1648 VSSD.n1646 0.0135208
R15799 VSSD.n3427 VSSD.n3426 0.0135208
R15800 VSSD.n3512 VSSD.n3509 0.0135208
R15801 VSSD.n152 VSSD.n144 0.0135208
R15802 VSSD.n206 VSSD.n201 0.0135208
R15803 VSSD.n580 VSSD.n571 0.0135208
R15804 VSSD.n729 VSSD.n542 0.0135208
R15805 VSSD.n744 VSSD 0.0122188
R15806 VSSD.n1445 VSSD 0.0122188
R15807 VSSD.n378 VSSD 0.0122188
R15808 VSSD.n3384 VSSD 0.0109167
R15809 VSSD.n1003 VSSD 0.0109167
R15810 VSSD.n1409 VSSD 0.0109167
R15811 VSSD.n2552 VSSD 0.00961458
R15812 VSSD.n851 VSSD.n839 0.0083125
R15813 VSSD.n3328 VSSD 0.0083125
R15814 VSSD.n3195 VSSD.n3194 0.0083125
R15815 VSSD.n3146 VSSD.n3145 0.0083125
R15816 VSSD.n2802 VSSD.n1348 0.0083125
R15817 VSSD.n2346 VSSD.n2345 0.0083125
R15818 VSSD.n2243 VSSD.n2123 0.0083125
R15819 VSSD.n1853 VSSD 0.0083125
R15820 VSSD.n1802 VSSD.n1673 0.0083125
R15821 VSSD.n3561 VSSD.n3560 0.0083125
R15822 VSSD.n341 VSSD.n227 0.0083125
R15823 VSSD.n3698 VSSD.n3697 0.0083125
R15824 VSSD.n3565 VSSD 0.00713529
R15825 VSSD.n3517 VSSD 0.00713529
R15826 VSSD.n3468 VSSD 0.00713529
R15827 VSSD.n3422 VSSD 0.00713529
R15828 VSSD VSSD.n3152 0.00701042
R15829 VSSD.n767 VSSD 0.00570833
R15830 VSSD.n1227 VSSD 0.00570833
R15831 VSSD.n2949 VSSD 0.00570833
R15832 VSSD.n2629 VSSD 0.00570833
R15833 VSSD VSSD.n2516 0.00570833
R15834 VSSD.n2045 VSSD 0.00570833
R15835 VSSD.n1898 VSSD 0.00570833
R15836 VSSD.n424 VSSD 0.00570833
R15837 VSSD.n2535 VSSD 0.00440625
R15838 VSSD.n958 VSSD.n844 0.00310417
R15839 VSSD.n1302 VSSD.n1134 0.00310417
R15840 VSSD.n3203 VSSD.n3202 0.00310417
R15841 VSSD.n2877 VSSD.n2854 0.00310417
R15842 VSSD.n3138 VSSD.n1061 0.00310417
R15843 VSSD.n2795 VSSD.n1358 0.00310417
R15844 VSSD.n1495 VSSD.n1476 0.00310417
R15845 VSSD.n2466 VSSD 0.00310417
R15846 VSSD.n2354 VSSD.n2353 0.00310417
R15847 VSSD.n1978 VSSD.n1955 0.00310417
R15848 VSSD.n2239 VSSD.n2126 0.00310417
R15849 VSSD.n1605 VSSD.n1572 0.00310417
R15850 VSSD.n1795 VSSD.n1683 0.00310417
R15851 VSSD.n3414 VSSD.n127 0.00310417
R15852 VSSD.n3569 VSSD.n3568 0.00310417
R15853 VSSD.n484 VSSD.n141 0.00310417
R15854 VSSD.n334 VSSD.n237 0.00310417
R15855 VSSD.n3707 VSSD.n22 0.00310417
R15856 a_6077_9813.n50 a_6077_9813.n49 330.05
R15857 a_6077_9813.n48 a_6077_9813.n3 327.253
R15858 a_6077_9813.n49 a_6077_9813.n2 217.256
R15859 a_6077_9813.n48 a_6077_9813.n4 217.256
R15860 a_6077_9813.n6 a_6077_9813.t34 212.081
R15861 a_6077_9813.n45 a_6077_9813.t21 212.081
R15862 a_6077_9813.n43 a_6077_9813.t39 212.081
R15863 a_6077_9813.n9 a_6077_9813.t37 212.081
R15864 a_6077_9813.n37 a_6077_9813.t22 212.081
R15865 a_6077_9813.n35 a_6077_9813.t12 212.081
R15866 a_6077_9813.n0 a_6077_9813.t25 212.081
R15867 a_6077_9813.n30 a_6077_9813.t14 212.081
R15868 a_6077_9813.n11 a_6077_9813.t26 212.081
R15869 a_6077_9813.n25 a_6077_9813.t35 212.081
R15870 a_6077_9813.n1 a_6077_9813.t33 212.081
R15871 a_6077_9813.n20 a_6077_9813.t20 212.081
R15872 a_6077_9813.n18 a_6077_9813.t38 212.081
R15873 a_6077_9813.n16 a_6077_9813.t28 212.081
R15874 a_6077_9813.n15 a_6077_9813.t8 212.081
R15875 a_6077_9813.n14 a_6077_9813.t30 212.081
R15876 a_6077_9813.n17 a_6077_9813.n13 169.409
R15877 a_6077_9813.n6 a_6077_9813.t36 162.274
R15878 a_6077_9813.n45 a_6077_9813.t13 162.274
R15879 a_6077_9813.n43 a_6077_9813.t9 162.274
R15880 a_6077_9813.n9 a_6077_9813.t31 162.274
R15881 a_6077_9813.n37 a_6077_9813.t32 162.274
R15882 a_6077_9813.n35 a_6077_9813.t24 162.274
R15883 a_6077_9813.n0 a_6077_9813.t29 162.274
R15884 a_6077_9813.n30 a_6077_9813.t27 162.274
R15885 a_6077_9813.n11 a_6077_9813.t17 162.274
R15886 a_6077_9813.n25 a_6077_9813.t23 162.274
R15887 a_6077_9813.n1 a_6077_9813.t10 162.274
R15888 a_6077_9813.n20 a_6077_9813.t18 162.274
R15889 a_6077_9813.n18 a_6077_9813.t15 162.274
R15890 a_6077_9813.n16 a_6077_9813.t11 162.274
R15891 a_6077_9813.n15 a_6077_9813.t19 162.274
R15892 a_6077_9813.n14 a_6077_9813.t16 162.274
R15893 a_6077_9813.n19 a_6077_9813.n13 152
R15894 a_6077_9813.n22 a_6077_9813.n21 152
R15895 a_6077_9813.n1 a_6077_9813.n23 152
R15896 a_6077_9813.n24 a_6077_9813.n12 152
R15897 a_6077_9813.n27 a_6077_9813.n26 152
R15898 a_6077_9813.n29 a_6077_9813.n28 152
R15899 a_6077_9813.n31 a_6077_9813.n10 152
R15900 a_6077_9813.n32 a_6077_9813.n0 152
R15901 a_6077_9813.n34 a_6077_9813.n33 152
R15902 a_6077_9813.n36 a_6077_9813.n8 152
R15903 a_6077_9813.n39 a_6077_9813.n38 152
R15904 a_6077_9813.n40 a_6077_9813.n7 152
R15905 a_6077_9813.n42 a_6077_9813.n41 152
R15906 a_6077_9813.n44 a_6077_9813.n5 152
R15907 a_6077_9813.n47 a_6077_9813.n46 152
R15908 a_6077_9813.n16 a_6077_9813.n15 55.2698
R15909 a_6077_9813.n15 a_6077_9813.n14 55.2698
R15910 a_6077_9813.n49 a_6077_9813.n48 44.0325
R15911 a_6077_9813.n21 a_6077_9813.n1 43.7018
R15912 a_6077_9813.n42 a_6077_9813.n7 43.7018
R15913 a_6077_9813.n0 a_6077_9813.n31 43.7018
R15914 a_6077_9813.n24 a_6077_9813.n1 43.7018
R15915 a_6077_9813.n34 a_6077_9813.n0 43.7018
R15916 a_6077_9813.n48 a_6077_9813.n47 43.5205
R15917 a_6077_9813.n2 a_6077_9813.t7 40.0005
R15918 a_6077_9813.n2 a_6077_9813.t6 40.0005
R15919 a_6077_9813.n4 a_6077_9813.t3 40.0005
R15920 a_6077_9813.n4 a_6077_9813.t4 40.0005
R15921 a_6077_9813.n44 a_6077_9813.n43 39.8458
R15922 a_6077_9813.n38 a_6077_9813.n9 35.9898
R15923 a_6077_9813.n17 a_6077_9813.n16 35.3472
R15924 a_6077_9813.n30 a_6077_9813.n29 33.4192
R15925 a_6077_9813.n26 a_6077_9813.n25 32.7765
R15926 a_6077_9813.n20 a_6077_9813.n19 31.4912
R15927 a_6077_9813.n36 a_6077_9813.n35 30.8485
R15928 a_6077_9813.n46 a_6077_9813.n45 28.2778
R15929 a_6077_9813.n3 a_6077_9813.t5 27.5805
R15930 a_6077_9813.n3 a_6077_9813.t1 27.5805
R15931 a_6077_9813.n50 a_6077_9813.t2 27.5805
R15932 a_6077_9813.t0 a_6077_9813.n50 27.5805
R15933 a_6077_9813.n46 a_6077_9813.n6 26.9925
R15934 a_6077_9813.n37 a_6077_9813.n36 24.4218
R15935 a_6077_9813.n19 a_6077_9813.n18 23.7792
R15936 a_6077_9813.n26 a_6077_9813.n11 22.4938
R15937 a_6077_9813.n29 a_6077_9813.n11 21.2085
R15938 a_6077_9813.n18 a_6077_9813.n17 19.9232
R15939 a_6077_9813.n38 a_6077_9813.n37 19.2805
R15940 a_6077_9813.n47 a_6077_9813.n5 17.4085
R15941 a_6077_9813.n41 a_6077_9813.n5 17.4085
R15942 a_6077_9813.n41 a_6077_9813.n40 17.4085
R15943 a_6077_9813.n40 a_6077_9813.n39 17.4085
R15944 a_6077_9813.n39 a_6077_9813.n8 17.4085
R15945 a_6077_9813.n33 a_6077_9813.n8 17.4085
R15946 a_6077_9813.n33 a_6077_9813.n32 17.4085
R15947 a_6077_9813.n32 a_6077_9813.n10 17.4085
R15948 a_6077_9813.n28 a_6077_9813.n10 17.4085
R15949 a_6077_9813.n28 a_6077_9813.n27 17.4085
R15950 a_6077_9813.n27 a_6077_9813.n12 17.4085
R15951 a_6077_9813.n23 a_6077_9813.n12 17.4085
R15952 a_6077_9813.n23 a_6077_9813.n22 17.4085
R15953 a_6077_9813.n22 a_6077_9813.n13 17.4085
R15954 a_6077_9813.n45 a_6077_9813.n44 15.4245
R15955 a_6077_9813.n35 a_6077_9813.n34 12.8538
R15956 a_6077_9813.n21 a_6077_9813.n20 12.2112
R15957 a_6077_9813.n25 a_6077_9813.n24 10.9258
R15958 a_6077_9813.n31 a_6077_9813.n30 10.2832
R15959 a_6077_9813.n9 a_6077_9813.n7 7.7125
R15960 a_6077_9813.n43 a_6077_9813.n42 3.8565
R15961 clknet_1_1__leaf_CLK.n2 clknet_1_1__leaf_CLK.n0 333.392
R15962 clknet_1_1__leaf_CLK.n2 clknet_1_1__leaf_CLK.n1 301.392
R15963 clknet_1_1__leaf_CLK.n4 clknet_1_1__leaf_CLK.n3 301.392
R15964 clknet_1_1__leaf_CLK.n6 clknet_1_1__leaf_CLK.n5 301.392
R15965 clknet_1_1__leaf_CLK.n8 clknet_1_1__leaf_CLK.n7 301.392
R15966 clknet_1_1__leaf_CLK.n49 clknet_1_1__leaf_CLK.n48 301.392
R15967 clknet_1_1__leaf_CLK.n51 clknet_1_1__leaf_CLK.n50 297.863
R15968 clknet_1_1__leaf_CLK.n42 clknet_1_1__leaf_CLK.t50 294.557
R15969 clknet_1_1__leaf_CLK.n37 clknet_1_1__leaf_CLK.t53 294.557
R15970 clknet_1_1__leaf_CLK.n27 clknet_1_1__leaf_CLK.t36 294.557
R15971 clknet_1_1__leaf_CLK.n24 clknet_1_1__leaf_CLK.t39 294.557
R15972 clknet_1_1__leaf_CLK.n32 clknet_1_1__leaf_CLK.t51 294.557
R15973 clknet_1_1__leaf_CLK.n30 clknet_1_1__leaf_CLK.t34 294.557
R15974 clknet_1_1__leaf_CLK.n22 clknet_1_1__leaf_CLK.t48 294.557
R15975 clknet_1_1__leaf_CLK.n19 clknet_1_1__leaf_CLK.t45 294.557
R15976 clknet_1_1__leaf_CLK.n16 clknet_1_1__leaf_CLK.t38 294.557
R15977 clknet_1_1__leaf_CLK.n14 clknet_1_1__leaf_CLK.t33 294.557
R15978 clknet_1_1__leaf_CLK.n9 clknet_1_1__leaf_CLK.t35 294.557
R15979 clknet_1_1__leaf_CLK.n11 clknet_1_1__leaf_CLK.t40 294.557
R15980 clknet_1_1__leaf_CLK.n46 clknet_1_1__leaf_CLK.n45 287.303
R15981 clknet_1_1__leaf_CLK.n54 clknet_1_1__leaf_CLK.n52 248.638
R15982 clknet_1_1__leaf_CLK.n42 clknet_1_1__leaf_CLK.t54 211.01
R15983 clknet_1_1__leaf_CLK.n37 clknet_1_1__leaf_CLK.t52 211.01
R15984 clknet_1_1__leaf_CLK.n27 clknet_1_1__leaf_CLK.t41 211.01
R15985 clknet_1_1__leaf_CLK.n24 clknet_1_1__leaf_CLK.t42 211.01
R15986 clknet_1_1__leaf_CLK.n32 clknet_1_1__leaf_CLK.t55 211.01
R15987 clknet_1_1__leaf_CLK.n30 clknet_1_1__leaf_CLK.t49 211.01
R15988 clknet_1_1__leaf_CLK.n22 clknet_1_1__leaf_CLK.t46 211.01
R15989 clknet_1_1__leaf_CLK.n19 clknet_1_1__leaf_CLK.t43 211.01
R15990 clknet_1_1__leaf_CLK.n16 clknet_1_1__leaf_CLK.t44 211.01
R15991 clknet_1_1__leaf_CLK.n14 clknet_1_1__leaf_CLK.t32 211.01
R15992 clknet_1_1__leaf_CLK.n9 clknet_1_1__leaf_CLK.t37 211.01
R15993 clknet_1_1__leaf_CLK.n11 clknet_1_1__leaf_CLK.t47 211.01
R15994 clknet_1_1__leaf_CLK.n54 clknet_1_1__leaf_CLK.n53 203.463
R15995 clknet_1_1__leaf_CLK.n56 clknet_1_1__leaf_CLK.n55 203.463
R15996 clknet_1_1__leaf_CLK.n60 clknet_1_1__leaf_CLK.n59 203.463
R15997 clknet_1_1__leaf_CLK.n62 clknet_1_1__leaf_CLK.n61 203.463
R15998 clknet_1_1__leaf_CLK.n64 clknet_1_1__leaf_CLK.n63 203.463
R15999 clknet_1_1__leaf_CLK.n58 clknet_1_1__leaf_CLK.n57 202.456
R16000 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n65 199.607
R16001 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n32 156.207
R16002 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n9 156.207
R16003 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n11 156.207
R16004 clknet_1_1__leaf_CLK.n43 clknet_1_1__leaf_CLK.n42 153.097
R16005 clknet_1_1__leaf_CLK.n28 clknet_1_1__leaf_CLK.n27 153.097
R16006 clknet_1_1__leaf_CLK.n17 clknet_1_1__leaf_CLK.n16 153.097
R16007 clknet_1_1__leaf_CLK.n38 clknet_1_1__leaf_CLK.n37 152
R16008 clknet_1_1__leaf_CLK.n25 clknet_1_1__leaf_CLK.n24 152
R16009 clknet_1_1__leaf_CLK.n31 clknet_1_1__leaf_CLK.n30 152
R16010 clknet_1_1__leaf_CLK.n23 clknet_1_1__leaf_CLK.n22 152
R16011 clknet_1_1__leaf_CLK.n20 clknet_1_1__leaf_CLK.n19 152
R16012 clknet_1_1__leaf_CLK.n15 clknet_1_1__leaf_CLK.n14 152
R16013 clknet_1_1__leaf_CLK.n56 clknet_1_1__leaf_CLK.n54 45.177
R16014 clknet_1_1__leaf_CLK.n62 clknet_1_1__leaf_CLK.n60 45.177
R16015 clknet_1_1__leaf_CLK.n64 clknet_1_1__leaf_CLK.n62 45.177
R16016 clknet_1_1__leaf_CLK.n58 clknet_1_1__leaf_CLK.n56 44.0476
R16017 clknet_1_1__leaf_CLK.n60 clknet_1_1__leaf_CLK.n58 44.0476
R16018 clknet_1_1__leaf_CLK.n52 clknet_1_1__leaf_CLK.t16 40.0005
R16019 clknet_1_1__leaf_CLK.n52 clknet_1_1__leaf_CLK.t28 40.0005
R16020 clknet_1_1__leaf_CLK.n53 clknet_1_1__leaf_CLK.t31 40.0005
R16021 clknet_1_1__leaf_CLK.n53 clknet_1_1__leaf_CLK.t18 40.0005
R16022 clknet_1_1__leaf_CLK.n55 clknet_1_1__leaf_CLK.t17 40.0005
R16023 clknet_1_1__leaf_CLK.n55 clknet_1_1__leaf_CLK.t21 40.0005
R16024 clknet_1_1__leaf_CLK.n57 clknet_1_1__leaf_CLK.t19 40.0005
R16025 clknet_1_1__leaf_CLK.n57 clknet_1_1__leaf_CLK.t20 40.0005
R16026 clknet_1_1__leaf_CLK.n59 clknet_1_1__leaf_CLK.t25 40.0005
R16027 clknet_1_1__leaf_CLK.n59 clknet_1_1__leaf_CLK.t22 40.0005
R16028 clknet_1_1__leaf_CLK.n61 clknet_1_1__leaf_CLK.t30 40.0005
R16029 clknet_1_1__leaf_CLK.n61 clknet_1_1__leaf_CLK.t24 40.0005
R16030 clknet_1_1__leaf_CLK.n63 clknet_1_1__leaf_CLK.t27 40.0005
R16031 clknet_1_1__leaf_CLK.n63 clknet_1_1__leaf_CLK.t29 40.0005
R16032 clknet_1_1__leaf_CLK.n65 clknet_1_1__leaf_CLK.t23 40.0005
R16033 clknet_1_1__leaf_CLK.n65 clknet_1_1__leaf_CLK.t26 40.0005
R16034 clknet_1_1__leaf_CLK.n4 clknet_1_1__leaf_CLK.n2 32.0005
R16035 clknet_1_1__leaf_CLK.n6 clknet_1_1__leaf_CLK.n4 32.0005
R16036 clknet_1_1__leaf_CLK.n47 clknet_1_1__leaf_CLK.n8 32.0005
R16037 clknet_1_1__leaf_CLK.n49 clknet_1_1__leaf_CLK.n47 32.0005
R16038 clknet_1_1__leaf_CLK.n8 clknet_1_1__leaf_CLK.n6 31.2005
R16039 clknet_1_1__leaf_CLK.n46 clknet_1_1__leaf_CLK.n44 30.612
R16040 clknet_1_1__leaf_CLK.n48 clknet_1_1__leaf_CLK.t1 27.5805
R16041 clknet_1_1__leaf_CLK.n48 clknet_1_1__leaf_CLK.t7 27.5805
R16042 clknet_1_1__leaf_CLK.n0 clknet_1_1__leaf_CLK.t4 27.5805
R16043 clknet_1_1__leaf_CLK.n0 clknet_1_1__leaf_CLK.t11 27.5805
R16044 clknet_1_1__leaf_CLK.n1 clknet_1_1__leaf_CLK.t0 27.5805
R16045 clknet_1_1__leaf_CLK.n1 clknet_1_1__leaf_CLK.t2 27.5805
R16046 clknet_1_1__leaf_CLK.n3 clknet_1_1__leaf_CLK.t10 27.5805
R16047 clknet_1_1__leaf_CLK.n3 clknet_1_1__leaf_CLK.t14 27.5805
R16048 clknet_1_1__leaf_CLK.n5 clknet_1_1__leaf_CLK.t9 27.5805
R16049 clknet_1_1__leaf_CLK.n5 clknet_1_1__leaf_CLK.t13 27.5805
R16050 clknet_1_1__leaf_CLK.n7 clknet_1_1__leaf_CLK.t8 27.5805
R16051 clknet_1_1__leaf_CLK.n7 clknet_1_1__leaf_CLK.t3 27.5805
R16052 clknet_1_1__leaf_CLK.n45 clknet_1_1__leaf_CLK.t5 27.5805
R16053 clknet_1_1__leaf_CLK.n45 clknet_1_1__leaf_CLK.t12 27.5805
R16054 clknet_1_1__leaf_CLK.n50 clknet_1_1__leaf_CLK.t15 27.5805
R16055 clknet_1_1__leaf_CLK.n50 clknet_1_1__leaf_CLK.t6 27.5805
R16056 clknet_1_1__leaf_CLK.n18 clknet_1_1__leaf_CLK.n17 21.2371
R16057 clknet_1_1__leaf_CLK.n34 clknet_1_1__leaf_CLK.n33 20.7375
R16058 clknet_1_1__leaf_CLK.n36 clknet_1_1__leaf_CLK 20.5068
R16059 clknet_1_1__leaf_CLK.n34 clknet_1_1__leaf_CLK 18.2951
R16060 clknet_1_1__leaf_CLK.n44 clknet_1_1__leaf_CLK.n43 16.5589
R16061 clknet_1_1__leaf_CLK.n29 clknet_1_1__leaf_CLK.n26 16.302
R16062 clknet_1_1__leaf_CLK.n18 clknet_1_1__leaf_CLK 15.5782
R16063 clknet_1_1__leaf_CLK.n47 clknet_1_1__leaf_CLK.n46 14.0898
R16064 clknet_1_1__leaf_CLK.n66 clknet_1_1__leaf_CLK.n64 13.177
R16065 clknet_1_1__leaf_CLK.n39 clknet_1_1__leaf_CLK 12.4091
R16066 clknet_1_1__leaf_CLK.n21 clknet_1_1__leaf_CLK 12.4091
R16067 clknet_1_1__leaf_CLK.n51 clknet_1_1__leaf_CLK.n49 10.4484
R16068 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n38 10.4234
R16069 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n31 10.4234
R16070 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n23 10.4234
R16071 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n20 10.4234
R16072 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n15 10.4234
R16073 clknet_1_1__leaf_CLK.n13 clknet_1_1__leaf_CLK.n12 10.416
R16074 clknet_1_1__leaf_CLK.n29 clknet_1_1__leaf_CLK 10.0149
R16075 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n28 9.55096
R16076 clknet_1_1__leaf_CLK.n26 clknet_1_1__leaf_CLK 9.32621
R16077 clknet_1_1__leaf_CLK.n33 clknet_1_1__leaf_CLK 9.32621
R16078 clknet_1_1__leaf_CLK.n10 clknet_1_1__leaf_CLK 9.32621
R16079 clknet_1_1__leaf_CLK.n12 clknet_1_1__leaf_CLK 9.32621
R16080 clknet_1_1__leaf_CLK.n13 clknet_1_1__leaf_CLK.n10 9.3005
R16081 clknet_1_1__leaf_CLK.n40 clknet_1_1__leaf_CLK.n39 6.86605
R16082 clknet_1_1__leaf_CLK.n41 clknet_1_1__leaf_CLK.n13 6.84249
R16083 clknet_1_1__leaf_CLK.n39 clknet_1_1__leaf_CLK.n36 6.04462
R16084 clknet_1_1__leaf_CLK.n21 clknet_1_1__leaf_CLK.n18 5.63391
R16085 clknet_1_1__leaf_CLK.n36 clknet_1_1__leaf_CLK.n35 4.5005
R16086 clknet_1_1__leaf_CLK.n41 clknet_1_1__leaf_CLK.n40 4.5005
R16087 clknet_1_1__leaf_CLK.n35 clknet_1_1__leaf_CLK.n34 3.20792
R16088 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n66 3.13183
R16089 clknet_1_1__leaf_CLK.n43 clknet_1_1__leaf_CLK 3.10907
R16090 clknet_1_1__leaf_CLK.n28 clknet_1_1__leaf_CLK 3.10907
R16091 clknet_1_1__leaf_CLK.n33 clknet_1_1__leaf_CLK 3.10907
R16092 clknet_1_1__leaf_CLK.n17 clknet_1_1__leaf_CLK 3.10907
R16093 clknet_1_1__leaf_CLK.n10 clknet_1_1__leaf_CLK 3.10907
R16094 clknet_1_1__leaf_CLK.n12 clknet_1_1__leaf_CLK 3.10907
R16095 clknet_1_1__leaf_CLK.n35 clknet_1_1__leaf_CLK.n29 2.90435
R16096 clknet_1_1__leaf_CLK.n44 clknet_1_1__leaf_CLK.n41 2.2972
R16097 clknet_1_1__leaf_CLK.n38 clknet_1_1__leaf_CLK 2.01193
R16098 clknet_1_1__leaf_CLK.n25 clknet_1_1__leaf_CLK 2.01193
R16099 clknet_1_1__leaf_CLK.n31 clknet_1_1__leaf_CLK 2.01193
R16100 clknet_1_1__leaf_CLK.n23 clknet_1_1__leaf_CLK 2.01193
R16101 clknet_1_1__leaf_CLK.n20 clknet_1_1__leaf_CLK 2.01193
R16102 clknet_1_1__leaf_CLK.n15 clknet_1_1__leaf_CLK 2.01193
R16103 clknet_1_1__leaf_CLK clknet_1_1__leaf_CLK.n51 1.75844
R16104 clknet_1_1__leaf_CLK.n40 clknet_1_1__leaf_CLK.n21 1.52676
R16105 clknet_1_1__leaf_CLK.n26 clknet_1_1__leaf_CLK.n25 1.09764
R16106 clknet_1_1__leaf_CLK.n66 clknet_1_1__leaf_CLK 0.604792
R16107 a_5515_4159.n4 a_5515_4159.n1 807.871
R16108 a_5515_4159.n0 a_5515_4159.t4 389.183
R16109 a_5515_4159.n5 a_5515_4159.n0 251.167
R16110 a_5515_4159.t0 a_5515_4159.n5 223.571
R16111 a_5515_4159.n2 a_5515_4159.t6 212.081
R16112 a_5515_4159.n3 a_5515_4159.t7 212.081
R16113 a_5515_4159.n4 a_5515_4159.n3 176.576
R16114 a_5515_4159.n0 a_5515_4159.t3 174.891
R16115 a_5515_4159.n2 a_5515_4159.t8 139.78
R16116 a_5515_4159.n3 a_5515_4159.t5 139.78
R16117 a_5515_4159.n1 a_5515_4159.t2 63.3219
R16118 a_5515_4159.n1 a_5515_4159.t1 63.3219
R16119 a_5515_4159.n3 a_5515_4159.n2 61.346
R16120 a_5515_4159.n5 a_5515_4159.n4 37.7195
R16121 a_5449_4233.n0 a_5449_4233.t0 68.3338
R16122 a_5449_4233.n0 a_5449_4233.t1 26.3935
R16123 a_5449_4233.n1 a_5449_4233.n0 14.4005
R16124 a_10329_5729.n3 a_10329_5729.n2 647.119
R16125 a_10329_5729.n1 a_10329_5729.t4 350.253
R16126 a_10329_5729.n2 a_10329_5729.n0 260.339
R16127 a_10329_5729.n2 a_10329_5729.n1 246.119
R16128 a_10329_5729.n1 a_10329_5729.t5 189.588
R16129 a_10329_5729.n3 a_10329_5729.t3 89.1195
R16130 a_10329_5729.n0 a_10329_5729.t1 63.3338
R16131 a_10329_5729.t2 a_10329_5729.n3 41.0422
R16132 a_10329_5729.n0 a_10329_5729.t0 31.9797
R16133 a_10207_5487.t0 a_10207_5487.t1 198.571
R16134 a_10373_5487.t0 a_10373_5487.t1 60.0005
R16135 CLKS.n365 CLKS.t57 408.63
R16136 CLKS.n42 CLKS.t50 408.63
R16137 CLKS.n34 CLKS.t66 408.63
R16138 CLKS.n351 CLKS.t87 408.63
R16139 CLKS.n118 CLKS.t56 408.63
R16140 CLKS.n104 CLKS.t119 408.63
R16141 CLKS.n98 CLKS.t130 408.63
R16142 CLKS.n78 CLKS.t74 408.63
R16143 CLKS.n51 CLKS.t34 408.63
R16144 CLKS.n320 CLKS.t109 408.63
R16145 CLKS.n254 CLKS.t107 408.63
R16146 CLKS.n238 CLKS.t31 408.63
R16147 CLKS.n227 CLKS.t112 408.63
R16148 CLKS.n221 CLKS.t91 408.63
R16149 CLKS.n199 CLKS.t76 408.63
R16150 CLKS.n177 CLKS.t52 408.63
R16151 CLKS.n185 CLKS.t30 408.63
R16152 CLKS.n171 CLKS.t93 408.63
R16153 CLKS.n308 CLKS.t140 408.63
R16154 CLKS.n284 CLKS.t85 408.63
R16155 CLKS.n278 CLKS.t55 408.63
R16156 CLKS.n266 CLKS.t105 408.63
R16157 CLKS.n302 CLKS.t46 408.63
R16158 CLKS.n153 CLKS.t24 408.63
R16159 CLKS.n335 CLKS.t90 408.63
R16160 CLKS.n148 CLKS.t23 408.63
R16161 CLKS.n136 CLKS.t70 408.63
R16162 CLKS.n20 CLKS.t123 408.63
R16163 CLKS.n10 CLKS.t60 408.63
R16164 CLKS.n8 CLKS.t94 408.63
R16165 CLKS.n361 CLKS.t127 347.577
R16166 CLKS.n45 CLKS.t49 347.577
R16167 CLKS.n39 CLKS.t137 347.577
R16168 CLKS.n347 CLKS.t38 347.577
R16169 CLKS.n122 CLKS.t89 347.577
R16170 CLKS.n110 CLKS.t117 347.577
R16171 CLKS.n94 CLKS.t82 347.577
R16172 CLKS.n84 CLKS.t19 347.577
R16173 CLKS.n57 CLKS.t106 347.577
R16174 CLKS.n325 CLKS.t78 347.577
R16175 CLKS.n249 CLKS.t36 347.577
R16176 CLKS.n243 CLKS.t32 347.577
R16177 CLKS.n232 CLKS.t115 347.577
R16178 CLKS.n216 CLKS.t18 347.577
R16179 CLKS.n204 CLKS.t111 347.577
R16180 CLKS.n182 CLKS.t20 347.577
R16181 CLKS.n190 CLKS.t58 347.577
R16182 CLKS.n166 CLKS.t120 347.577
R16183 CLKS.n312 CLKS.t68 347.577
R16184 CLKS.n289 CLKS.t86 347.577
R16185 CLKS.n274 CLKS.t98 347.577
R16186 CLKS.n261 CLKS.t33 347.577
R16187 CLKS.n297 CLKS.t48 347.577
R16188 CLKS.n158 CLKS.t81 347.577
R16189 CLKS.n331 CLKS.t16 347.577
R16190 CLKS.n145 CLKS.t21 347.577
R16191 CLKS.n132 CLKS.t101 347.577
R16192 CLKS.n26 CLKS.t135 347.577
R16193 CLKS.n14 CLKS.t103 347.577
R16194 CLKS.n4 CLKS.t104 347.577
R16195 CLKS.n209 CLKS.t121 261.887
R16196 CLKS.n196 CLKS.t100 261.887
R16197 CLKS.n161 CLKS.t51 230.576
R16198 CLKS.n74 CLKS.n63 205.28
R16199 CLKS.n73 CLKS.n64 205.28
R16200 CLKS.n62 CLKS.n61 205.28
R16201 CLKS.n361 CLKS.t35 193.337
R16202 CLKS.n45 CLKS.t75 193.337
R16203 CLKS.n39 CLKS.t114 193.337
R16204 CLKS.n347 CLKS.t132 193.337
R16205 CLKS.n122 CLKS.t139 193.337
R16206 CLKS.n110 CLKS.t122 193.337
R16207 CLKS.n94 CLKS.t47 193.337
R16208 CLKS.n84 CLKS.t26 193.337
R16209 CLKS.n57 CLKS.t84 193.337
R16210 CLKS.n325 CLKS.t54 193.337
R16211 CLKS.n249 CLKS.t62 193.337
R16212 CLKS.n243 CLKS.t129 193.337
R16213 CLKS.n232 CLKS.t92 193.337
R16214 CLKS.n216 CLKS.t71 193.337
R16215 CLKS.n204 CLKS.t118 193.337
R16216 CLKS.n182 CLKS.t72 193.337
R16217 CLKS.n190 CLKS.t40 193.337
R16218 CLKS.n166 CLKS.t102 193.337
R16219 CLKS.n312 CLKS.t128 193.337
R16220 CLKS.n289 CLKS.t69 193.337
R16221 CLKS.n274 CLKS.t42 193.337
R16222 CLKS.n261 CLKS.t96 193.337
R16223 CLKS.n297 CLKS.t28 193.337
R16224 CLKS.n158 CLKS.t17 193.337
R16225 CLKS.n331 CLKS.t83 193.337
R16226 CLKS.n145 CLKS.t126 193.337
R16227 CLKS.n132 CLKS.t44 193.337
R16228 CLKS.n26 CLKS.t113 193.337
R16229 CLKS.n14 CLKS.t27 193.337
R16230 CLKS.n4 CLKS.t79 193.337
R16231 CLKS.n77 CLKS.n76 190.911
R16232 CLKS CLKS.n34 165.201
R16233 CLKS CLKS.n104 165.201
R16234 CLKS CLKS.n51 165.201
R16235 CLKS CLKS.n148 165.201
R16236 CLKS CLKS.n20 165.201
R16237 CLKS CLKS.n10 165.201
R16238 CLKS CLKS.n8 165.201
R16239 CLKS.n119 CLKS.n118 165.117
R16240 CLKS.n79 CLKS.n78 165.117
R16241 CLKS.n49 CLKS.n42 165.072
R16242 CLKS.n321 CLKS.n320 165.072
R16243 CLKS.n255 CLKS.n254 165.072
R16244 CLKS.n239 CLKS.n238 165.072
R16245 CLKS.n228 CLKS.n227 165.072
R16246 CLKS.n222 CLKS.n221 165.072
R16247 CLKS.n208 CLKS.n199 165.072
R16248 CLKS.n178 CLKS.n177 165.072
R16249 CLKS.n194 CLKS.n185 165.072
R16250 CLKS.n172 CLKS.n171 165.072
R16251 CLKS.n309 CLKS.n308 165.072
R16252 CLKS.n285 CLKS.n284 165.072
R16253 CLKS.n267 CLKS.n266 165.072
R16254 CLKS.n303 CLKS.n302 165.072
R16255 CLKS.n154 CLKS.n153 165.072
R16256 CLKS.n336 CLKS.n335 165.072
R16257 CLKS.n161 CLKS.t108 158.275
R16258 CLKS.n366 CLKS.n365 158.144
R16259 CLKS.n352 CLKS.n351 158.144
R16260 CLKS.n99 CLKS.n98 158.144
R16261 CLKS.n279 CLKS.n278 158.144
R16262 CLKS.n137 CLKS.n136 158.144
R16263 CLKS.n162 CLKS.n161 156.268
R16264 CLKS.n209 CLKS.t73 155.847
R16265 CLKS.n196 CLKS.t37 155.847
R16266 CLKS.n210 CLKS.n209 153.13
R16267 CLKS.n197 CLKS.n196 152.512
R16268 CLKS.n362 CLKS.n361 152
R16269 CLKS.n46 CLKS.n45 152
R16270 CLKS.n40 CLKS.n39 152
R16271 CLKS.n348 CLKS.n347 152
R16272 CLKS.n123 CLKS.n122 152
R16273 CLKS.n111 CLKS.n110 152
R16274 CLKS.n95 CLKS.n94 152
R16275 CLKS.n85 CLKS.n84 152
R16276 CLKS.n58 CLKS.n57 152
R16277 CLKS.n326 CLKS.n325 152
R16278 CLKS.n250 CLKS.n249 152
R16279 CLKS.n244 CLKS.n243 152
R16280 CLKS.n233 CLKS.n232 152
R16281 CLKS.n217 CLKS.n216 152
R16282 CLKS.n205 CLKS.n204 152
R16283 CLKS.n183 CLKS.n182 152
R16284 CLKS.n191 CLKS.n190 152
R16285 CLKS.n167 CLKS.n166 152
R16286 CLKS.n313 CLKS.n312 152
R16287 CLKS.n290 CLKS.n289 152
R16288 CLKS.n275 CLKS.n274 152
R16289 CLKS.n262 CLKS.n261 152
R16290 CLKS.n298 CLKS.n297 152
R16291 CLKS.n159 CLKS.n158 152
R16292 CLKS.n332 CLKS.n331 152
R16293 CLKS.n146 CLKS.n145 152
R16294 CLKS.n133 CLKS.n132 152
R16295 CLKS.n27 CLKS.n26 152
R16296 CLKS.n15 CLKS.n14 152
R16297 CLKS.n5 CLKS.n4 152
R16298 CLKS.n365 CLKS.t141 132.282
R16299 CLKS.n42 CLKS.t125 132.282
R16300 CLKS.n34 CLKS.t99 132.282
R16301 CLKS.n351 CLKS.t116 132.282
R16302 CLKS.n118 CLKS.t43 132.282
R16303 CLKS.n104 CLKS.t59 132.282
R16304 CLKS.n98 CLKS.t25 132.282
R16305 CLKS.n78 CLKS.t131 132.282
R16306 CLKS.n51 CLKS.t64 132.282
R16307 CLKS.n320 CLKS.t29 132.282
R16308 CLKS.n254 CLKS.t80 132.282
R16309 CLKS.n238 CLKS.t77 132.282
R16310 CLKS.n227 CLKS.t39 132.282
R16311 CLKS.n221 CLKS.t88 132.282
R16312 CLKS.n199 CLKS.t133 132.282
R16313 CLKS.n177 CLKS.t138 132.282
R16314 CLKS.n185 CLKS.t61 132.282
R16315 CLKS.n171 CLKS.t136 132.282
R16316 CLKS.n308 CLKS.t22 132.282
R16317 CLKS.n284 CLKS.t134 132.282
R16318 CLKS.n278 CLKS.t53 132.282
R16319 CLKS.n266 CLKS.t110 132.282
R16320 CLKS.n302 CLKS.t97 132.282
R16321 CLKS.n153 CLKS.t41 132.282
R16322 CLKS.n335 CLKS.t67 132.282
R16323 CLKS.n148 CLKS.t63 132.282
R16324 CLKS.n136 CLKS.t65 132.282
R16325 CLKS.n20 CLKS.t124 132.282
R16326 CLKS.n10 CLKS.t45 132.282
R16327 CLKS.n8 CLKS.t95 132.282
R16328 CLKS.n69 CLKS.n68 99.1759
R16329 CLKS.n72 CLKS.n65 99.1749
R16330 CLKS.n71 CLKS.n66 99.1749
R16331 CLKS.n70 CLKS.n67 99.1749
R16332 CLKS.n74 CLKS.n73 38.4005
R16333 CLKS.n75 CLKS.n62 38.4005
R16334 CLKS.n75 CLKS.n74 38.4005
R16335 CLKS.n72 CLKS.n71 34.3584
R16336 CLKS.n71 CLKS.n70 34.3584
R16337 CLKS.n70 CLKS.n69 34.3584
R16338 CLKS CLKS.n72 34.0948
R16339 CLKS.n69 CLKS 32.411
R16340 CLKS.n73 CLKS 30.14
R16341 CLKS.n366 CLKS.n358 27.7325
R16342 CLKS.n352 CLKS.n342 27.7325
R16343 CLKS.n99 CLKS.n91 27.7325
R16344 CLKS.n279 CLKS.n271 27.7325
R16345 CLKS.n137 CLKS.n129 27.7325
R16346 CLKS CLKS.n62 27.6358
R16347 CLKS.n76 CLKS.t9 26.5955
R16348 CLKS.n76 CLKS.t14 26.5955
R16349 CLKS.n63 CLKS.t0 26.5955
R16350 CLKS.n63 CLKS.t12 26.5955
R16351 CLKS.n64 CLKS.t3 26.5955
R16352 CLKS.n64 CLKS.t7 26.5955
R16353 CLKS.n61 CLKS.t1 26.5955
R16354 CLKS.n61 CLKS.t4 26.5955
R16355 CLKS.n90 CLKS.n77 25.4745
R16356 CLKS.n65 CLKS.t5 24.9236
R16357 CLKS.n65 CLKS.t11 24.9236
R16358 CLKS.n66 CLKS.t13 24.9236
R16359 CLKS.n66 CLKS.t8 24.9236
R16360 CLKS.n67 CLKS.t2 24.9236
R16361 CLKS.n67 CLKS.t10 24.9236
R16362 CLKS.n68 CLKS.t15 24.9236
R16363 CLKS.n68 CLKS.t6 24.9236
R16364 CLKS.n211 CLKS.n208 19.5495
R16365 CLKS.n163 CLKS.n162 17.2898
R16366 CLKS.n357 CLKS.n356 15.2364
R16367 CLKS.n247 CLKS.n246 14.9196
R16368 CLKS.n294 CLKS.n293 14.881
R16369 CLKS.n77 CLKS.n75 14.3703
R16370 CLKS.n327 CLKS 14.0185
R16371 CLKS.n245 CLKS 14.0185
R16372 CLKS CLKS.n231 14.0185
R16373 CLKS CLKS.n165 14.0185
R16374 CLKS.n291 CLKS 14.0185
R16375 CLKS CLKS.n296 14.0185
R16376 CLKS CLKS.n360 13.8338
R16377 CLKS CLKS.n44 13.8338
R16378 CLKS CLKS.n121 13.8338
R16379 CLKS CLKS.n93 13.8338
R16380 CLKS.n184 CLKS 13.8338
R16381 CLKS CLKS.n273 13.8338
R16382 CLKS.n160 CLKS 13.8338
R16383 CLKS CLKS.n131 13.8338
R16384 CLKS CLKS.n13 13.8338
R16385 CLKS.n293 CLKS.n282 13.0706
R16386 CLKS.n318 CLKS.n317 13.0596
R16387 CLKS.n213 CLKS.n212 12.5829
R16388 CLKS.n330 CLKS.n329 12.1444
R16389 CLKS.n363 CLKS.n362 12.0681
R16390 CLKS.n47 CLKS.n46 12.0681
R16391 CLKS.n41 CLKS.n40 12.0681
R16392 CLKS.n349 CLKS.n348 12.0681
R16393 CLKS.n124 CLKS.n123 12.0681
R16394 CLKS.n112 CLKS.n111 12.0681
R16395 CLKS.n96 CLKS.n95 12.0681
R16396 CLKS.n86 CLKS.n85 12.0681
R16397 CLKS.n59 CLKS.n58 12.0681
R16398 CLKS.n206 CLKS.n205 12.0681
R16399 CLKS.n192 CLKS.n191 12.0681
R16400 CLKS.n276 CLKS.n275 12.0681
R16401 CLKS.n147 CLKS.n146 12.0681
R16402 CLKS.n134 CLKS.n133 12.0681
R16403 CLKS.n28 CLKS.n27 12.0681
R16404 CLKS.n16 CLKS.n15 12.0681
R16405 CLKS.n6 CLKS.n5 12.0681
R16406 CLKS.n212 CLKS.n211 11.5913
R16407 CLKS.n195 CLKS.n184 10.7699
R16408 CLKS.n329 CLKS.n328 10.4663
R16409 CLKS.n38 CLKS.n37 9.86717
R16410 CLKS.n346 CLKS.n345 9.86717
R16411 CLKS.n109 CLKS.n108 9.86717
R16412 CLKS.n83 CLKS.n82 9.86717
R16413 CLKS.n56 CLKS.n55 9.86717
R16414 CLKS.n203 CLKS.n202 9.86717
R16415 CLKS.n189 CLKS.n188 9.86717
R16416 CLKS.n144 CLKS.n143 9.86717
R16417 CLKS.n25 CLKS.n24 9.86717
R16418 CLKS.n3 CLKS.n2 9.86717
R16419 CLKS.n198 CLKS.n197 9.66056
R16420 CLKS.n231 CLKS 9.37931
R16421 CLKS.n165 CLKS 9.37931
R16422 CLKS.n296 CLKS 9.37931
R16423 CLKS.n367 CLKS.n366 9.3005
R16424 CLKS.n37 CLKS.n36 9.3005
R16425 CLKS.n345 CLKS.n344 9.3005
R16426 CLKS.n353 CLKS.n352 9.3005
R16427 CLKS.n108 CLKS.n107 9.3005
R16428 CLKS.n100 CLKS.n99 9.3005
R16429 CLKS.n82 CLKS.n81 9.3005
R16430 CLKS.n55 CLKS.n54 9.3005
R16431 CLKS.n324 CLKS.n323 9.3005
R16432 CLKS.n328 CLKS.n327 9.3005
R16433 CLKS.n252 CLKS.n251 9.3005
R16434 CLKS.n242 CLKS.n241 9.3005
R16435 CLKS.n246 CLKS.n245 9.3005
R16436 CLKS.n235 CLKS.n234 9.3005
R16437 CLKS.n219 CLKS.n218 9.3005
R16438 CLKS.n202 CLKS.n201 9.3005
R16439 CLKS.n211 CLKS.n210 9.3005
R16440 CLKS.n181 CLKS.n180 9.3005
R16441 CLKS.n188 CLKS.n187 9.3005
R16442 CLKS.n169 CLKS.n168 9.3005
R16443 CLKS.n315 CLKS.n314 9.3005
R16444 CLKS.n288 CLKS.n287 9.3005
R16445 CLKS.n292 CLKS.n291 9.3005
R16446 CLKS.n280 CLKS.n279 9.3005
R16447 CLKS.n264 CLKS.n263 9.3005
R16448 CLKS.n300 CLKS.n299 9.3005
R16449 CLKS.n157 CLKS.n156 9.3005
R16450 CLKS.n334 CLKS.n333 9.3005
R16451 CLKS.n143 CLKS.n142 9.3005
R16452 CLKS.n138 CLKS.n137 9.3005
R16453 CLKS.n24 CLKS.n23 9.3005
R16454 CLKS.n2 CLKS.n1 9.3005
R16455 CLKS.n128 CLKS.n117 8.82605
R16456 CLKS.n362 CLKS 8.82212
R16457 CLKS.n46 CLKS 8.82212
R16458 CLKS.n40 CLKS.n38 8.82212
R16459 CLKS.n348 CLKS.n346 8.82212
R16460 CLKS.n123 CLKS 8.82212
R16461 CLKS.n111 CLKS.n109 8.82212
R16462 CLKS.n95 CLKS 8.82212
R16463 CLKS.n85 CLKS.n83 8.82212
R16464 CLKS.n58 CLKS.n56 8.82212
R16465 CLKS.n205 CLKS.n203 8.82212
R16466 CLKS.n191 CLKS.n189 8.82212
R16467 CLKS.n275 CLKS 8.82212
R16468 CLKS.n146 CLKS.n144 8.82212
R16469 CLKS.n133 CLKS 8.82212
R16470 CLKS.n27 CLKS.n25 8.82212
R16471 CLKS.n15 CLKS 8.82212
R16472 CLKS.n5 CLKS.n3 8.82212
R16473 CLKS.n117 CLKS.n116 8.61863
R16474 CLKS.n32 CLKS.n19 8.41671
R16475 CLKS.n340 CLKS.n128 8.36314
R16476 CLKS.n50 CLKS 7.58395
R16477 CLKS.n341 CLKS.n340 6.75425
R16478 CLKS.n356 CLKS.n355 6.49363
R16479 CLKS.n151 CLKS.n140 6.19006
R16480 CLKS.n371 CLKS 6.10421
R16481 CLKS.n214 CLKS.n163 5.92684
R16482 CLKS.n195 CLKS.n194 5.7623
R16483 CLKS.n294 CLKS.n270 5.58292
R16484 CLKS.n339 CLKS.n338 5.43457
R16485 CLKS.n50 CLKS.n49 5.33372
R16486 CLKS.n213 CLKS.n175 4.99885
R16487 CLKS.n307 CLKS.n306 4.83577
R16488 CLKS.n236 CLKS 4.76939
R16489 CLKS.n316 CLKS 4.76939
R16490 CLKS CLKS.n326 4.67077
R16491 CLKS.n250 CLKS 4.67077
R16492 CLKS CLKS.n244 4.67077
R16493 CLKS.n233 CLKS 4.67077
R16494 CLKS.n217 CLKS 4.67077
R16495 CLKS CLKS.n183 4.67077
R16496 CLKS.n167 CLKS 4.67077
R16497 CLKS.n313 CLKS 4.67077
R16498 CLKS CLKS.n290 4.67077
R16499 CLKS.n262 CLKS 4.67077
R16500 CLKS.n298 CLKS 4.67077
R16501 CLKS CLKS.n159 4.67077
R16502 CLKS.n332 CLKS 4.67077
R16503 CLKS.n37 CLKS 4.53383
R16504 CLKS.n345 CLKS 4.53383
R16505 CLKS.n108 CLKS 4.53383
R16506 CLKS.n82 CLKS 4.53383
R16507 CLKS.n55 CLKS 4.53383
R16508 CLKS.n327 CLKS 4.53383
R16509 CLKS.n245 CLKS 4.53383
R16510 CLKS.n231 CLKS 4.53383
R16511 CLKS.n202 CLKS 4.53383
R16512 CLKS.n188 CLKS 4.53383
R16513 CLKS.n165 CLKS 4.53383
R16514 CLKS.n291 CLKS 4.53383
R16515 CLKS.n296 CLKS 4.53383
R16516 CLKS.n143 CLKS 4.53383
R16517 CLKS.n24 CLKS 4.53383
R16518 CLKS.n2 CLKS 4.53383
R16519 CLKS.n151 CLKS.n150 4.50133
R16520 CLKS.n90 CLKS.n89 4.5005
R16521 CLKS.n103 CLKS.n102 4.5005
R16522 CLKS.n116 CLKS.n115 4.5005
R16523 CLKS.n128 CLKS.n127 4.5005
R16524 CLKS.n226 CLKS.n225 4.5005
R16525 CLKS.n259 CLKS.n258 4.5005
R16526 CLKS.n32 CLKS.n31 4.5005
R16527 CLKS.n370 CLKS.n369 4.5005
R16528 CLKS.n163 CLKS 4.49111
R16529 CLKS.n317 CLKS.n259 4.4222
R16530 CLKS.n197 CLKS 4.3525
R16531 CLKS.n236 CLKS.n226 3.2255
R16532 CLKS.n116 CLKS.n103 3.20792
R16533 CLKS.n339 CLKS.n151 3.20792
R16534 CLKS.n210 CLKS 3.2005
R16535 CLKS.n324 CLKS 2.94104
R16536 CLKS.n251 CLKS 2.94104
R16537 CLKS.n242 CLKS 2.94104
R16538 CLKS.n234 CLKS 2.94104
R16539 CLKS.n218 CLKS 2.94104
R16540 CLKS.n181 CLKS 2.94104
R16541 CLKS.n168 CLKS 2.94104
R16542 CLKS.n314 CLKS 2.94104
R16543 CLKS.n288 CLKS 2.94104
R16544 CLKS.n263 CLKS 2.94104
R16545 CLKS.n299 CLKS 2.94104
R16546 CLKS.n157 CLKS 2.94104
R16547 CLKS.n333 CLKS 2.94104
R16548 CLKS.n316 CLKS.n307 2.77907
R16549 CLKS.n326 CLKS.n324 2.76807
R16550 CLKS.n251 CLKS.n250 2.76807
R16551 CLKS.n244 CLKS.n242 2.76807
R16552 CLKS.n234 CLKS.n233 2.76807
R16553 CLKS.n218 CLKS.n217 2.76807
R16554 CLKS.n183 CLKS.n181 2.76807
R16555 CLKS.n168 CLKS.n167 2.76807
R16556 CLKS.n314 CLKS.n313 2.76807
R16557 CLKS.n290 CLKS.n288 2.76807
R16558 CLKS.n263 CLKS.n262 2.76807
R16559 CLKS.n299 CLKS.n298 2.76807
R16560 CLKS.n159 CLKS.n157 2.76807
R16561 CLKS.n333 CLKS.n332 2.76807
R16562 CLKS.n253 CLKS 2.75496
R16563 CLKS.n220 CLKS 2.75496
R16564 CLKS.n265 CLKS 2.75496
R16565 CLKS.n301 CLKS 2.75496
R16566 CLKS.n21 CLKS 2.64782
R16567 CLKS.n117 CLKS.n60 2.55957
R16568 CLKS.n162 CLKS 2.4005
R16569 CLKS CLKS.n364 2.36657
R16570 CLKS CLKS.n48 2.36657
R16571 CLKS.n35 CLKS 2.36657
R16572 CLKS CLKS.n350 2.36657
R16573 CLKS CLKS.n97 2.36657
R16574 CLKS.n52 CLKS 2.36657
R16575 CLKS CLKS.n322 2.36657
R16576 CLKS CLKS.n240 2.36657
R16577 CLKS CLKS.n229 2.36657
R16578 CLKS CLKS.n207 2.36657
R16579 CLKS CLKS.n179 2.36657
R16580 CLKS CLKS.n193 2.36657
R16581 CLKS CLKS.n310 2.36657
R16582 CLKS CLKS.n286 2.36657
R16583 CLKS CLKS.n277 2.36657
R16584 CLKS CLKS.n155 2.36657
R16585 CLKS CLKS.n337 2.36657
R16586 CLKS.n149 CLKS 2.36657
R16587 CLKS CLKS.n135 2.36657
R16588 CLKS.n126 CLKS.n125 2.24604
R16589 CLKS.n88 CLKS.n87 2.24604
R16590 CLKS.n105 CLKS 2.23711
R16591 CLKS.n9 CLKS 2.23711
R16592 CLKS.n226 CLKS.n214 2.14885
R16593 CLKS.n329 CLKS.n318 1.98814
R16594 CLKS CLKS.n370 1.90229
R16595 CLKS.n257 CLKS.n256 1.88889
R16596 CLKS.n224 CLKS.n223 1.88889
R16597 CLKS.n269 CLKS.n268 1.88889
R16598 CLKS.n305 CLKS.n304 1.88889
R16599 CLKS.n11 CLKS 1.88889
R16600 CLKS.n30 CLKS.n29 1.83532
R16601 CLKS.n38 CLKS 1.73023
R16602 CLKS.n346 CLKS 1.73023
R16603 CLKS.n109 CLKS 1.73023
R16604 CLKS.n83 CLKS 1.73023
R16605 CLKS.n56 CLKS 1.73023
R16606 CLKS.n203 CLKS 1.73023
R16607 CLKS.n189 CLKS 1.73023
R16608 CLKS.n144 CLKS 1.73023
R16609 CLKS.n25 CLKS 1.73023
R16610 CLKS.n3 CLKS 1.73023
R16611 CLKS.n170 CLKS 1.52282
R16612 CLKS.n126 CLKS 1.49329
R16613 CLKS.n88 CLKS 1.49329
R16614 CLKS.n114 CLKS.n113 1.42461
R16615 CLKS.n170 CLKS 1.42461
R16616 CLKS.n372 CLKS.n7 1.42461
R16617 CLKS.n103 CLKS.n90 1.38649
R16618 CLKS.n370 CLKS.n32 1.38649
R16619 CLKS.n356 CLKS.n50 1.38099
R16620 CLKS.n212 CLKS.n198 1.34528
R16621 CLKS.n257 CLKS 1.32983
R16622 CLKS.n224 CLKS 1.32983
R16623 CLKS.n269 CLKS 1.32983
R16624 CLKS.n305 CLKS 1.32983
R16625 CLKS.n30 CLKS 1.27213
R16626 CLKS.n247 CLKS.n236 1.13903
R16627 CLKS.n259 CLKS.n247 1.08292
R16628 CLKS.n340 CLKS.n339 1.08292
R16629 CLKS.n114 CLKS 1.05098
R16630 CLKS CLKS.n372 1.05098
R16631 CLKS.n11 CLKS 1.00496
R16632 CLKS.n317 CLKS.n316 0.728316
R16633 CLKS.n174 CLKS 0.666365
R16634 CLKS.n105 CLKS 0.65675
R16635 CLKS.n174 CLKS.n173 0.65675
R16636 CLKS.n9 CLKS 0.65675
R16637 CLKS.n318 CLKS.n160 0.628411
R16638 CLKS.n322 CLKS 0.580857
R16639 CLKS.n256 CLKS 0.580857
R16640 CLKS.n240 CLKS 0.580857
R16641 CLKS.n229 CLKS 0.580857
R16642 CLKS.n223 CLKS 0.580857
R16643 CLKS.n179 CLKS 0.580857
R16644 CLKS.n173 CLKS 0.580857
R16645 CLKS.n310 CLKS 0.580857
R16646 CLKS.n286 CLKS 0.580857
R16647 CLKS.n268 CLKS 0.580857
R16648 CLKS.n304 CLKS 0.580857
R16649 CLKS.n155 CLKS 0.580857
R16650 CLKS.n337 CLKS 0.580857
R16651 CLKS.n364 CLKS 0.527286
R16652 CLKS.n48 CLKS 0.527286
R16653 CLKS.n35 CLKS 0.527286
R16654 CLKS.n350 CLKS 0.527286
R16655 CLKS.n125 CLKS 0.527286
R16656 CLKS.n113 CLKS 0.527286
R16657 CLKS.n97 CLKS 0.527286
R16658 CLKS.n87 CLKS 0.527286
R16659 CLKS.n52 CLKS 0.527286
R16660 CLKS.n207 CLKS 0.527286
R16661 CLKS.n193 CLKS 0.527286
R16662 CLKS.n277 CLKS 0.527286
R16663 CLKS.n149 CLKS 0.527286
R16664 CLKS.n135 CLKS 0.527286
R16665 CLKS.n29 CLKS 0.527286
R16666 CLKS.n17 CLKS 0.527286
R16667 CLKS.n7 CLKS 0.527286
R16668 CLKS.n293 CLKS.n292 0.44984
R16669 CLKS.n91 CLKS 0.418351
R16670 CLKS.n271 CLKS 0.418351
R16671 CLKS.n129 CLKS 0.418351
R16672 CLKS.n214 CLKS.n213 0.401393
R16673 CLKS.n18 CLKS 0.387519
R16674 CLKS.n341 CLKS 0.351043
R16675 CLKS.n357 CLKS 0.351043
R16676 CLKS.n307 CLKS.n294 0.327423
R16677 CLKS.n21 CLKS 0.246036
R16678 CLKS.n321 CLKS 0.225552
R16679 CLKS.n255 CLKS 0.225552
R16680 CLKS.n239 CLKS 0.225552
R16681 CLKS.n228 CLKS 0.225552
R16682 CLKS.n222 CLKS 0.225552
R16683 CLKS.n178 CLKS 0.225552
R16684 CLKS.n172 CLKS 0.225552
R16685 CLKS.n309 CLKS 0.225552
R16686 CLKS.n285 CLKS 0.225552
R16687 CLKS.n267 CLKS 0.225552
R16688 CLKS.n303 CLKS 0.225552
R16689 CLKS.n154 CLKS 0.225552
R16690 CLKS.n336 CLKS 0.225552
R16691 CLKS.n359 CLKS 0.196446
R16692 CLKS.n43 CLKS 0.196446
R16693 CLKS.n33 CLKS 0.196446
R16694 CLKS.n343 CLKS 0.196446
R16695 CLKS.n120 CLKS 0.196446
R16696 CLKS.n106 CLKS 0.196446
R16697 CLKS.n92 CLKS 0.196446
R16698 CLKS.n80 CLKS 0.196446
R16699 CLKS.n53 CLKS 0.196446
R16700 CLKS.n319 CLKS 0.196446
R16701 CLKS.n248 CLKS 0.196446
R16702 CLKS.n237 CLKS 0.196446
R16703 CLKS.n230 CLKS 0.196446
R16704 CLKS.n215 CLKS 0.196446
R16705 CLKS.n200 CLKS 0.196446
R16706 CLKS.n176 CLKS 0.196446
R16707 CLKS.n186 CLKS 0.196446
R16708 CLKS.n164 CLKS 0.196446
R16709 CLKS.n311 CLKS 0.196446
R16710 CLKS.n283 CLKS 0.196446
R16711 CLKS.n272 CLKS 0.196446
R16712 CLKS.n260 CLKS 0.196446
R16713 CLKS.n295 CLKS 0.196446
R16714 CLKS.n152 CLKS 0.196446
R16715 CLKS.n330 CLKS 0.196446
R16716 CLKS.n141 CLKS 0.196446
R16717 CLKS.n130 CLKS 0.196446
R16718 CLKS.n22 CLKS 0.196446
R16719 CLKS.n12 CLKS 0.196446
R16720 CLKS.n0 CLKS 0.196446
R16721 CLKS.n253 CLKS 0.192464
R16722 CLKS.n220 CLKS 0.192464
R16723 CLKS.n265 CLKS 0.192464
R16724 CLKS.n301 CLKS 0.192464
R16725 CLKS.n18 CLKS.n17 0.192464
R16726 CLKS.n101 CLKS 0.15675
R16727 CLKS.n281 CLKS 0.15675
R16728 CLKS.n139 CLKS 0.15675
R16729 CLKS.n354 CLKS 0.15675
R16730 CLKS.n368 CLKS 0.15675
R16731 CLKS.n49 CLKS 0.128681
R16732 CLKS.n322 CLKS.n321 0.128681
R16733 CLKS.n256 CLKS.n255 0.128681
R16734 CLKS.n240 CLKS.n239 0.128681
R16735 CLKS.n229 CLKS.n228 0.128681
R16736 CLKS.n223 CLKS.n222 0.128681
R16737 CLKS.n208 CLKS 0.128681
R16738 CLKS.n179 CLKS.n178 0.128681
R16739 CLKS.n194 CLKS 0.128681
R16740 CLKS.n173 CLKS.n172 0.128681
R16741 CLKS.n310 CLKS.n309 0.128681
R16742 CLKS.n286 CLKS.n285 0.128681
R16743 CLKS.n268 CLKS.n267 0.128681
R16744 CLKS.n304 CLKS.n303 0.128681
R16745 CLKS.n155 CLKS.n154 0.128681
R16746 CLKS.n337 CLKS.n336 0.128681
R16747 CLKS.n198 CLKS.n195 0.1255
R16748 CLKS.n119 CLKS 0.11596
R16749 CLKS.n79 CLKS 0.11596
R16750 CLKS.n368 CLKS.n367 0.0983261
R16751 CLKS.n354 CLKS.n353 0.0983261
R16752 CLKS.n101 CLKS.n100 0.0983261
R16753 CLKS.n281 CLKS.n280 0.0983261
R16754 CLKS.n139 CLKS.n138 0.0983261
R16755 CLKS.n360 CLKS.n359 0.0793043
R16756 CLKS.n360 CLKS 0.0793043
R16757 CLKS.n367 CLKS 0.0793043
R16758 CLKS.n44 CLKS.n43 0.0793043
R16759 CLKS.n44 CLKS 0.0793043
R16760 CLKS.n36 CLKS.n33 0.0793043
R16761 CLKS.n36 CLKS 0.0793043
R16762 CLKS.n344 CLKS.n343 0.0793043
R16763 CLKS.n344 CLKS 0.0793043
R16764 CLKS.n353 CLKS 0.0793043
R16765 CLKS.n121 CLKS.n120 0.0793043
R16766 CLKS.n121 CLKS 0.0793043
R16767 CLKS.n107 CLKS.n106 0.0793043
R16768 CLKS.n107 CLKS 0.0793043
R16769 CLKS.n93 CLKS.n92 0.0793043
R16770 CLKS.n93 CLKS 0.0793043
R16771 CLKS.n100 CLKS 0.0793043
R16772 CLKS.n81 CLKS.n80 0.0793043
R16773 CLKS.n81 CLKS 0.0793043
R16774 CLKS.n54 CLKS.n53 0.0793043
R16775 CLKS.n54 CLKS 0.0793043
R16776 CLKS.n328 CLKS 0.0793043
R16777 CLKS.n246 CLKS 0.0793043
R16778 CLKS.n201 CLKS.n200 0.0793043
R16779 CLKS.n201 CLKS 0.0793043
R16780 CLKS.n184 CLKS 0.0793043
R16781 CLKS.n187 CLKS.n186 0.0793043
R16782 CLKS.n187 CLKS 0.0793043
R16783 CLKS.n292 CLKS 0.0793043
R16784 CLKS.n273 CLKS.n272 0.0793043
R16785 CLKS.n273 CLKS 0.0793043
R16786 CLKS.n280 CLKS 0.0793043
R16787 CLKS.n160 CLKS 0.0793043
R16788 CLKS.n142 CLKS.n141 0.0793043
R16789 CLKS.n142 CLKS 0.0793043
R16790 CLKS.n131 CLKS.n130 0.0793043
R16791 CLKS.n131 CLKS 0.0793043
R16792 CLKS.n138 CLKS 0.0793043
R16793 CLKS.n23 CLKS.n22 0.0793043
R16794 CLKS.n23 CLKS 0.0793043
R16795 CLKS.n13 CLKS.n12 0.0793043
R16796 CLKS.n13 CLKS 0.0793043
R16797 CLKS.n1 CLKS.n0 0.0793043
R16798 CLKS.n1 CLKS 0.0793043
R16799 CLKS.n115 CLKS.n105 0.0774231
R16800 CLKS.n115 CLKS.n114 0.0774231
R16801 CLKS.n102 CLKS.n101 0.0774231
R16802 CLKS.n258 CLKS.n253 0.0774231
R16803 CLKS.n258 CLKS.n257 0.0774231
R16804 CLKS.n225 CLKS.n220 0.0774231
R16805 CLKS.n225 CLKS.n224 0.0774231
R16806 CLKS.n175 CLKS.n170 0.0774231
R16807 CLKS.n175 CLKS.n174 0.0774231
R16808 CLKS.n282 CLKS.n281 0.0774231
R16809 CLKS.n270 CLKS.n265 0.0774231
R16810 CLKS.n270 CLKS.n269 0.0774231
R16811 CLKS.n306 CLKS.n301 0.0774231
R16812 CLKS.n306 CLKS.n305 0.0774231
R16813 CLKS.n140 CLKS.n139 0.0774231
R16814 CLKS.n355 CLKS.n354 0.0774231
R16815 CLKS.n369 CLKS.n368 0.0774231
R16816 CLKS.n31 CLKS.n21 0.0774231
R16817 CLKS.n31 CLKS.n30 0.0774231
R16818 CLKS.n19 CLKS.n11 0.0774231
R16819 CLKS.n19 CLKS.n18 0.0774231
R16820 CLKS.n371 CLKS.n9 0.0774231
R16821 CLKS.n372 CLKS.n371 0.0774231
R16822 CLKS.n342 CLKS.n341 0.0678077
R16823 CLKS.n358 CLKS.n357 0.0678077
R16824 CLKS CLKS.n126 0.0654038
R16825 CLKS CLKS.n88 0.0654038
R16826 CLKS.n127 CLKS.n119 0.0634968
R16827 CLKS.n89 CLKS.n79 0.0634968
R16828 CLKS.n364 CLKS.n363 0.03675
R16829 CLKS.n363 CLKS 0.03675
R16830 CLKS.n48 CLKS.n47 0.03675
R16831 CLKS.n47 CLKS 0.03675
R16832 CLKS.n41 CLKS.n35 0.03675
R16833 CLKS CLKS.n41 0.03675
R16834 CLKS.n350 CLKS.n349 0.03675
R16835 CLKS.n349 CLKS 0.03675
R16836 CLKS.n125 CLKS.n124 0.03675
R16837 CLKS.n124 CLKS 0.03675
R16838 CLKS.n113 CLKS.n112 0.03675
R16839 CLKS.n112 CLKS 0.03675
R16840 CLKS.n97 CLKS.n96 0.03675
R16841 CLKS.n96 CLKS 0.03675
R16842 CLKS.n87 CLKS.n86 0.03675
R16843 CLKS.n86 CLKS 0.03675
R16844 CLKS.n59 CLKS 0.03675
R16845 CLKS.n323 CLKS.n319 0.03675
R16846 CLKS.n323 CLKS 0.03675
R16847 CLKS.n252 CLKS.n248 0.03675
R16848 CLKS CLKS.n252 0.03675
R16849 CLKS.n241 CLKS.n237 0.03675
R16850 CLKS.n241 CLKS 0.03675
R16851 CLKS.n235 CLKS.n230 0.03675
R16852 CLKS CLKS.n235 0.03675
R16853 CLKS.n219 CLKS.n215 0.03675
R16854 CLKS CLKS.n219 0.03675
R16855 CLKS.n207 CLKS.n206 0.03675
R16856 CLKS.n206 CLKS 0.03675
R16857 CLKS.n180 CLKS.n176 0.03675
R16858 CLKS.n180 CLKS 0.03675
R16859 CLKS.n193 CLKS.n192 0.03675
R16860 CLKS.n192 CLKS 0.03675
R16861 CLKS.n169 CLKS.n164 0.03675
R16862 CLKS CLKS.n169 0.03675
R16863 CLKS.n315 CLKS.n311 0.03675
R16864 CLKS CLKS.n315 0.03675
R16865 CLKS.n287 CLKS.n283 0.03675
R16866 CLKS.n287 CLKS 0.03675
R16867 CLKS.n277 CLKS.n276 0.03675
R16868 CLKS.n276 CLKS 0.03675
R16869 CLKS.n264 CLKS.n260 0.03675
R16870 CLKS CLKS.n264 0.03675
R16871 CLKS.n300 CLKS.n295 0.03675
R16872 CLKS CLKS.n300 0.03675
R16873 CLKS.n156 CLKS.n152 0.03675
R16874 CLKS.n156 CLKS 0.03675
R16875 CLKS.n334 CLKS.n330 0.03675
R16876 CLKS.n147 CLKS 0.03675
R16877 CLKS.n135 CLKS.n134 0.03675
R16878 CLKS.n134 CLKS 0.03675
R16879 CLKS.n29 CLKS.n28 0.03675
R16880 CLKS.n28 CLKS 0.03675
R16881 CLKS.n17 CLKS.n16 0.03675
R16882 CLKS.n16 CLKS 0.03675
R16883 CLKS.n7 CLKS.n6 0.03675
R16884 CLKS.n6 CLKS 0.03675
R16885 CLKS.n60 CLKS.n52 0.02175
R16886 CLKS.n338 CLKS 0.02175
R16887 CLKS.n150 CLKS.n149 0.02121
R16888 CLKS.n150 CLKS.n147 0.0155106
R16889 CLKS.n60 CLKS.n59 0.0155
R16890 CLKS.n338 CLKS.n334 0.0155
R16891 CLKS.n127 CLKS 0.0125192
R16892 CLKS.n89 CLKS 0.0125192
R16893 CLKS.n102 CLKS.n91 0.0101154
R16894 CLKS.n282 CLKS.n271 0.0101154
R16895 CLKS.n140 CLKS.n129 0.0101154
R16896 CLKS.n355 CLKS.n342 0.0101154
R16897 CLKS.n369 CLKS.n358 0.0101154
R16898 CLKS.n359 CLKS 0.00725676
R16899 CLKS.n43 CLKS 0.00725676
R16900 CLKS CLKS.n33 0.00725676
R16901 CLKS.n343 CLKS 0.00725676
R16902 CLKS.n120 CLKS 0.00725676
R16903 CLKS.n106 CLKS 0.00725676
R16904 CLKS.n92 CLKS 0.00725676
R16905 CLKS.n80 CLKS 0.00725676
R16906 CLKS.n53 CLKS 0.00725676
R16907 CLKS.n319 CLKS 0.00725676
R16908 CLKS CLKS.n248 0.00725676
R16909 CLKS.n237 CLKS 0.00725676
R16910 CLKS CLKS.n230 0.00725676
R16911 CLKS CLKS.n215 0.00725676
R16912 CLKS.n200 CLKS 0.00725676
R16913 CLKS.n176 CLKS 0.00725676
R16914 CLKS.n186 CLKS 0.00725676
R16915 CLKS CLKS.n164 0.00725676
R16916 CLKS CLKS.n311 0.00725676
R16917 CLKS.n283 CLKS 0.00725676
R16918 CLKS.n272 CLKS 0.00725676
R16919 CLKS CLKS.n260 0.00725676
R16920 CLKS CLKS.n295 0.00725676
R16921 CLKS.n152 CLKS 0.00725676
R16922 CLKS CLKS.n330 0.00725676
R16923 CLKS.n141 CLKS 0.00725676
R16924 CLKS.n130 CLKS 0.00725676
R16925 CLKS.n22 CLKS 0.00725676
R16926 CLKS.n12 CLKS 0.00725676
R16927 CLKS.n0 CLKS 0.00725676
R16928 CF[0].n2 CF[0].t10 294.557
R16929 CF[0].n0 CF[0].t8 294.557
R16930 CF[0].n16 CF[0].n15 289.096
R16931 CF[0].n11 CF[0].t9 235.763
R16932 CF[0].n5 CF[0].t6 221.72
R16933 CF[0].n6 CF[0].t7 221.72
R16934 CF[0].n2 CF[0].t4 211.01
R16935 CF[0].n0 CF[0].t11 211.01
R16936 CF[0].n18 CF[0].n17 185
R16937 CF[0].n11 CF[0].t5 163.464
R16938 CF[0].n1 CF[0].n0 153.097
R16939 CF[0].n8 CF[0].n7 152
R16940 CF[0].n10 CF[0].n9 152
R16941 CF[0].n12 CF[0].n11 152
R16942 CF[0].n3 CF[0].n2 152
R16943 CF[0].n5 CF[0].t12 149.421
R16944 CF[0].n6 CF[0].t13 149.421
R16945 CF[0].n7 CF[0].n6 58.019
R16946 CF[0].n18 CF[0] 49.0339
R16947 CF[0].n10 CF[0].n5 43.7375
R16948 CF[0].n20 CF[0].n14 29.8563
R16949 CF[0].n15 CF[0].t3 26.5955
R16950 CF[0].n15 CF[0].t1 26.5955
R16951 CF[0] CF[0].n20 25.9746
R16952 CF[0].n17 CF[0].t0 24.9236
R16953 CF[0].n17 CF[0].t2 24.9236
R16954 CF[0].n13 CF[0].n4 24.6413
R16955 CF[0].n9 CF[0] 20.8005
R16956 CF[0].n13 CF[0].n12 20.1268
R16957 CF[0].n11 CF[0].n10 17.8524
R16958 CF[0].n7 CF[0].n5 16.9598
R16959 CF[0].n8 CF[0] 16.3205
R16960 CF[0] CF[0].n8 13.1205
R16961 CF[0].n14 CF[0].n13 10.6063
R16962 CF[0].n14 CF[0].n1 9.79203
R16963 CF[0] CF[0].n16 9.48653
R16964 CF[0].n4 CF[0] 9.32621
R16965 CF[0].n20 CF[0].n19 9.3005
R16966 CF[0].n9 CF[0] 8.6405
R16967 CF[0].n16 CF[0] 7.7181
R16968 CF[0].n19 CF[0].n18 6.1445
R16969 CF[0].n19 CF[0] 4.3525
R16970 CF[0].n1 CF[0] 3.10907
R16971 CF[0].n3 CF[0] 2.01193
R16972 CF[0].n4 CF[0].n3 1.09764
R16973 CF[0].n12 CF[0] 0.9605
R16974 a_4463_8893.n1 a_4463_8893.t6 530.01
R16975 a_4463_8893.t0 a_4463_8893.n5 421.021
R16976 a_4463_8893.n0 a_4463_8893.t4 337.171
R16977 a_4463_8893.n3 a_4463_8893.t1 280.223
R16978 a_4463_8893.n4 a_4463_8893.t2 263.173
R16979 a_4463_8893.n4 a_4463_8893.t5 227.826
R16980 a_4463_8893.n0 a_4463_8893.t3 199.762
R16981 a_4463_8893.n2 a_4463_8893.n1 170.81
R16982 a_4463_8893.n2 a_4463_8893.n0 167.321
R16983 a_4463_8893.n5 a_4463_8893.n4 152
R16984 a_4463_8893.n1 a_4463_8893.t7 141.923
R16985 a_4463_8893.n3 a_4463_8893.n2 10.8376
R16986 a_4463_8893.n5 a_4463_8893.n3 2.50485
R16987 a_10667_9813.n5 a_10667_9813.n4 807.871
R16988 a_10667_9813.n2 a_10667_9813.t3 389.183
R16989 a_10667_9813.n3 a_10667_9813.n2 251.167
R16990 a_10667_9813.n3 a_10667_9813.t1 223.571
R16991 a_10667_9813.n0 a_10667_9813.t6 212.081
R16992 a_10667_9813.n1 a_10667_9813.t8 212.081
R16993 a_10667_9813.n4 a_10667_9813.n1 176.576
R16994 a_10667_9813.n2 a_10667_9813.t5 174.891
R16995 a_10667_9813.n0 a_10667_9813.t4 139.78
R16996 a_10667_9813.n1 a_10667_9813.t7 139.78
R16997 a_10667_9813.t0 a_10667_9813.n5 63.3219
R16998 a_10667_9813.n5 a_10667_9813.t2 63.3219
R16999 a_10667_9813.n1 a_10667_9813.n0 61.346
R17000 a_10667_9813.n4 a_10667_9813.n3 37.7195
R17001 a_10654_10205.t0 a_10654_10205.t1 126.644
R17002 a_4259_3861.n1 a_4259_3861.t4 530.01
R17003 a_4259_3861.t0 a_4259_3861.n5 421.021
R17004 a_4259_3861.n0 a_4259_3861.t6 337.142
R17005 a_4259_3861.n3 a_4259_3861.t1 280.223
R17006 a_4259_3861.n4 a_4259_3861.t2 263.173
R17007 a_4259_3861.n4 a_4259_3861.t5 227.826
R17008 a_4259_3861.n0 a_4259_3861.t7 199.762
R17009 a_4259_3861.n2 a_4259_3861.n1 170.81
R17010 a_4259_3861.n2 a_4259_3861.n0 167.321
R17011 a_4259_3861.n5 a_4259_3861.n4 152
R17012 a_4259_3861.n1 a_4259_3861.t3 141.923
R17013 a_4259_3861.n3 a_4259_3861.n2 10.8376
R17014 a_4259_3861.n5 a_4259_3861.n3 2.50485
R17015 a_4425_3861.t0 a_4425_3861.n3 370.026
R17016 a_4425_3861.n0 a_4425_3861.t3 351.356
R17017 a_4425_3861.n1 a_4425_3861.t5 334.717
R17018 a_4425_3861.n3 a_4425_3861.t1 325.971
R17019 a_4425_3861.n1 a_4425_3861.t2 309.935
R17020 a_4425_3861.n0 a_4425_3861.t4 305.683
R17021 a_4425_3861.n2 a_4425_3861.n0 16.879
R17022 a_4425_3861.n3 a_4425_3861.n2 10.8867
R17023 a_4425_3861.n2 a_4425_3861.n1 9.3005
R17024 EN.n217 EN.t54 408.63
R17025 EN.n202 EN.t10 408.63
R17026 EN.n170 EN.t20 408.63
R17027 EN.n156 EN.t76 408.63
R17028 EN.n121 EN.t79 408.63
R17029 EN.n134 EN.t35 408.63
R17030 EN.n148 EN.t7 408.63
R17031 EN.n185 EN.t13 408.63
R17032 EN.n112 EN.t53 408.63
R17033 EN.n100 EN.t87 408.63
R17034 EN.n85 EN.t24 408.63
R17035 EN.n82 EN.t88 408.63
R17036 EN.n67 EN.t36 408.63
R17037 EN.n58 EN.t3 408.63
R17038 EN.n233 EN.t33 408.63
R17039 EN.n243 EN.t12 408.63
R17040 EN.n44 EN.t14 408.63
R17041 EN.n38 EN.t75 408.63
R17042 EN.n26 EN.t73 408.63
R17043 EN.n11 EN.t60 408.63
R17044 EN.n256 EN.t77 408.63
R17045 EN.n8 EN.t48 408.63
R17046 EN.n220 EN.t69 347.577
R17047 EN.n205 EN.t72 347.577
R17048 EN.n173 EN.t18 347.577
R17049 EN.n158 EN.t16 347.577
R17050 EN.n116 EN.t34 347.577
R17051 EN.n129 EN.t1 347.577
R17052 EN.n143 EN.t61 347.577
R17053 EN.n188 EN.t19 347.577
R17054 EN.n107 EN.t44 347.577
R17055 EN.n95 EN.t81 347.577
R17056 EN.n90 EN.t26 347.577
R17057 EN.n77 EN.t59 347.577
R17058 EN.n70 EN.t4 347.577
R17059 EN.n61 EN.t46 347.577
R17060 EN.n229 EN.t31 347.577
R17061 EN.n238 EN.t40 347.577
R17062 EN.n50 EN.t21 347.577
R17063 EN.n34 EN.t5 347.577
R17064 EN.n22 EN.t2 347.577
R17065 EN.n14 EN.t32 347.577
R17066 EN.n251 EN.t63 347.577
R17067 EN.n4 EN.t11 347.577
R17068 EN.n126 EN.t74 333.651
R17069 EN.n126 EN.t38 297.233
R17070 EN.n127 EN.n126 196.493
R17071 EN.n220 EN.t86 193.337
R17072 EN.n205 EN.t25 193.337
R17073 EN.n173 EN.t66 193.337
R17074 EN.n158 EN.t64 193.337
R17075 EN.n116 EN.t42 193.337
R17076 EN.n129 EN.t62 193.337
R17077 EN.n143 EN.t68 193.337
R17078 EN.n188 EN.t70 193.337
R17079 EN.n107 EN.t57 193.337
R17080 EN.n95 EN.t49 193.337
R17081 EN.n90 EN.t29 193.337
R17082 EN.n77 EN.t80 193.337
R17083 EN.n70 EN.t51 193.337
R17084 EN.n61 EN.t8 193.337
R17085 EN.n229 EN.t47 193.337
R17086 EN.n238 EN.t0 193.337
R17087 EN.n50 EN.t27 193.337
R17088 EN.n34 EN.t71 193.337
R17089 EN.n22 EN.t6 193.337
R17090 EN.n14 EN.t50 193.337
R17091 EN.n251 EN.t83 193.337
R17092 EN.n4 EN.t52 193.337
R17093 EN EN.n217 165.201
R17094 EN EN.n44 165.201
R17095 EN EN.n11 165.201
R17096 EN EN.n8 165.201
R17097 EN.n122 EN.n121 165.072
R17098 EN.n135 EN.n134 165.072
R17099 EN.n149 EN.n148 165.072
R17100 EN.n113 EN.n112 165.072
R17101 EN.n101 EN.n100 165.072
R17102 EN.n86 EN.n85 165.072
R17103 EN.n83 EN.n82 165.072
R17104 EN.n75 EN.n67 165.072
R17105 EN.n66 EN.n58 165.072
R17106 EN.n234 EN.n233 165.072
R17107 EN.n244 EN.n243 165.072
R17108 EN.n257 EN.n256 165.072
R17109 EN.n211 EN.n202 158.144
R17110 EN.n179 EN.n170 158.144
R17111 EN.n164 EN.n156 158.144
R17112 EN.n194 EN.n185 158.144
R17113 EN.n39 EN.n38 158.144
R17114 EN.n27 EN.n26 158.144
R17115 EN.n221 EN.n220 152
R17116 EN.n206 EN.n205 152
R17117 EN.n174 EN.n173 152
R17118 EN.n159 EN.n158 152
R17119 EN.n117 EN.n116 152
R17120 EN.n130 EN.n129 152
R17121 EN.n144 EN.n143 152
R17122 EN.n189 EN.n188 152
R17123 EN.n108 EN.n107 152
R17124 EN.n96 EN.n95 152
R17125 EN.n91 EN.n90 152
R17126 EN.n78 EN.n77 152
R17127 EN.n71 EN.n70 152
R17128 EN.n62 EN.n61 152
R17129 EN.n230 EN.n229 152
R17130 EN.n239 EN.n238 152
R17131 EN.n51 EN.n50 152
R17132 EN.n35 EN.n34 152
R17133 EN.n23 EN.n22 152
R17134 EN.n15 EN.n14 152
R17135 EN.n252 EN.n251 152
R17136 EN.n5 EN.n4 152
R17137 EN.n217 EN.t22 132.282
R17138 EN.n202 EN.t15 132.282
R17139 EN.n170 EN.t82 132.282
R17140 EN.n156 EN.t78 132.282
R17141 EN.n121 EN.t41 132.282
R17142 EN.n134 EN.t58 132.282
R17143 EN.n148 EN.t67 132.282
R17144 EN.n185 EN.t17 132.282
R17145 EN.n112 EN.t28 132.282
R17146 EN.n100 EN.t39 132.282
R17147 EN.n85 EN.t85 132.282
R17148 EN.n82 EN.t56 132.282
R17149 EN.n67 EN.t43 132.282
R17150 EN.n58 EN.t9 132.282
R17151 EN.n233 EN.t30 132.282
R17152 EN.n243 EN.t84 132.282
R17153 EN.n44 EN.t37 132.282
R17154 EN.n38 EN.t89 132.282
R17155 EN.n26 EN.t23 132.282
R17156 EN.n11 EN.t55 132.282
R17157 EN.n256 EN.t45 132.282
R17158 EN.n8 EN.t65 132.282
R17159 EN.n139 EN.n127 37.6104
R17160 EN.n57 EN.n56 30.0335
R17161 EN.n212 EN.n211 27.7325
R17162 EN.n180 EN.n179 27.7325
R17163 EN.n165 EN.n164 27.7325
R17164 EN.n195 EN.n194 27.7325
R17165 EN.n39 EN.n31 27.7325
R17166 EN.n27 EN.n17 27.7325
R17167 EN.n224 EN 14.8875
R17168 EN EN.n204 14.0185
R17169 EN EN.n172 14.0185
R17170 EN EN.n115 14.0185
R17171 EN EN.n142 14.0185
R17172 EN EN.n187 14.0185
R17173 EN.n92 EN 14.0185
R17174 EN EN.n69 14.0185
R17175 EN EN.n60 14.0185
R17176 EN EN.n237 14.0185
R17177 EN.n222 EN 13.8338
R17178 EN EN.n33 13.8338
R17179 EN EN.n13 13.8338
R17180 EN.n221 EN.n219 12.0681
R17181 EN.n52 EN.n51 12.0681
R17182 EN.n36 EN.n35 12.0681
R17183 EN.n24 EN.n23 12.0681
R17184 EN.n16 EN.n15 12.0681
R17185 EN.n6 EN.n5 12.0681
R17186 EN.n215 EN.n214 11.2313
R17187 EN.n223 EN.n215 10.4469
R17188 EN.n226 EN.n225 10.1186
R17189 EN.n197 EN.n196 10.0829
R17190 EN.n199 EN.n105 9.88649
R17191 EN.n49 EN.n48 9.86717
R17192 EN.n21 EN.n20 9.86717
R17193 EN.n3 EN.n2 9.86717
R17194 EN.n197 EN.n182 9.82056
R17195 EN.n204 EN 9.37931
R17196 EN.n172 EN 9.37931
R17197 EN.n115 EN 9.37931
R17198 EN.n142 EN 9.37931
R17199 EN.n187 EN 9.37931
R17200 EN.n69 EN 9.37931
R17201 EN.n60 EN 9.37931
R17202 EN.n237 EN 9.37931
R17203 EN.n208 EN.n207 9.3005
R17204 EN.n211 EN.n210 9.3005
R17205 EN.n176 EN.n175 9.3005
R17206 EN.n179 EN.n178 9.3005
R17207 EN.n161 EN.n160 9.3005
R17208 EN.n164 EN.n163 9.3005
R17209 EN.n119 EN.n118 9.3005
R17210 EN.n132 EN.n131 9.3005
R17211 EN.n146 EN.n145 9.3005
R17212 EN.n191 EN.n190 9.3005
R17213 EN.n194 EN.n193 9.3005
R17214 EN.n110 EN.n109 9.3005
R17215 EN.n98 EN.n97 9.3005
R17216 EN.n89 EN.n88 9.3005
R17217 EN.n93 EN.n92 9.3005
R17218 EN.n80 EN.n79 9.3005
R17219 EN.n73 EN.n72 9.3005
R17220 EN.n64 EN.n63 9.3005
R17221 EN.n228 EN.n227 9.3005
R17222 EN.n241 EN.n240 9.3005
R17223 EN.n48 EN.n47 9.3005
R17224 EN.n40 EN.n39 9.3005
R17225 EN.n20 EN.n19 9.3005
R17226 EN.n28 EN.n27 9.3005
R17227 EN.n254 EN.n253 9.3005
R17228 EN.n2 EN.n1 9.3005
R17229 EN.n199 EN.n198 8.95242
R17230 EN.n105 EN.n93 8.91275
R17231 EN EN.n221 8.82212
R17232 EN.n51 EN.n49 8.82212
R17233 EN.n35 EN 8.82212
R17234 EN.n23 EN.n21 8.82212
R17235 EN.n15 EN 8.82212
R17236 EN.n5 EN.n3 8.82212
R17237 EN.n226 EN 8.19287
R17238 EN.n259 EN.n258 7.70792
R17239 EN.n249 EN.n57 6.94555
R17240 EN.n224 EN.n223 6.89885
R17241 EN.n57 EN 6.09082
R17242 EN.n235 EN 5.9301
R17243 EN.n43 EN.n30 5.88649
R17244 EN.n225 EN.n224 5.58292
R17245 EN.n258 EN 5.10867
R17246 EN.n140 EN.n125 4.84592
R17247 EN.n153 EN.n152 4.84592
R17248 EN.n153 EN.n140 4.73264
R17249 EN.n206 EN 4.67077
R17250 EN.n174 EN 4.67077
R17251 EN.n159 EN 4.67077
R17252 EN.n117 EN 4.67077
R17253 EN.n130 EN 4.67077
R17254 EN.n144 EN 4.67077
R17255 EN.n189 EN 4.67077
R17256 EN.n108 EN 4.67077
R17257 EN.n96 EN 4.67077
R17258 EN EN.n91 4.67077
R17259 EN.n78 EN 4.67077
R17260 EN.n71 EN 4.67077
R17261 EN.n62 EN 4.67077
R17262 EN EN.n230 4.67077
R17263 EN.n239 EN 4.67077
R17264 EN.n252 EN 4.67077
R17265 EN.n204 EN 4.53383
R17266 EN.n172 EN 4.53383
R17267 EN.n115 EN 4.53383
R17268 EN.n142 EN 4.53383
R17269 EN.n187 EN 4.53383
R17270 EN.n92 EN 4.53383
R17271 EN.n69 EN 4.53383
R17272 EN.n60 EN 4.53383
R17273 EN.n237 EN 4.53383
R17274 EN.n48 EN 4.53383
R17275 EN.n20 EN 4.53383
R17276 EN.n2 EN 4.53383
R17277 EN.n139 EN.n138 4.5005
R17278 EN.n167 EN.n166 4.5005
R17279 EN.n182 EN.n181 4.5005
R17280 EN.n105 EN.n104 4.5005
R17281 EN.n214 EN.n213 4.5005
R17282 EN.n43 EN.n42 4.5005
R17283 EN.n56 EN.n55 4.5005
R17284 EN.n248 EN.n247 4.5005
R17285 EN.n198 EN.n197 4.45242
R17286 EN.n56 EN.n43 3.90435
R17287 EN.n167 EN.n153 3.21135
R17288 EN.n248 EN.n235 3.20792
R17289 EN.n207 EN 2.94104
R17290 EN.n175 EN 2.94104
R17291 EN.n160 EN 2.94104
R17292 EN.n118 EN 2.94104
R17293 EN.n131 EN 2.94104
R17294 EN.n145 EN 2.94104
R17295 EN.n190 EN 2.94104
R17296 EN.n109 EN 2.94104
R17297 EN.n97 EN 2.94104
R17298 EN.n89 EN 2.94104
R17299 EN.n79 EN 2.94104
R17300 EN.n72 EN 2.94104
R17301 EN.n63 EN 2.94104
R17302 EN.n228 EN 2.94104
R17303 EN.n240 EN 2.94104
R17304 EN.n253 EN 2.94104
R17305 EN.n207 EN.n206 2.76807
R17306 EN.n175 EN.n174 2.76807
R17307 EN.n160 EN.n159 2.76807
R17308 EN.n118 EN.n117 2.76807
R17309 EN.n131 EN.n130 2.76807
R17310 EN.n145 EN.n144 2.76807
R17311 EN.n190 EN.n189 2.76807
R17312 EN.n109 EN.n108 2.76807
R17313 EN.n97 EN.n96 2.76807
R17314 EN.n91 EN.n89 2.76807
R17315 EN.n79 EN.n78 2.76807
R17316 EN.n72 EN.n71 2.76807
R17317 EN.n63 EN.n62 2.76807
R17318 EN.n230 EN.n228 2.76807
R17319 EN.n240 EN.n239 2.76807
R17320 EN.n253 EN.n252 2.76807
R17321 EN.n120 EN 2.75496
R17322 EN.n147 EN 2.75496
R17323 EN.n99 EN 2.75496
R17324 EN.n45 EN 2.64782
R17325 EN.n9 EN 2.64782
R17326 EN.n225 EN 2.4301
R17327 EN.n218 EN 2.36657
R17328 EN.n209 EN 2.36657
R17329 EN.n177 EN 2.36657
R17330 EN.n162 EN 2.36657
R17331 EN.n192 EN 2.36657
R17332 EN.n111 EN 2.36657
R17333 EN EN.n87 2.36657
R17334 EN.n81 EN 2.36657
R17335 EN.n74 EN 2.36657
R17336 EN.n65 EN 2.36657
R17337 EN.n232 EN 2.36657
R17338 EN EN.n37 2.36657
R17339 EN EN.n25 2.36657
R17340 EN.n12 EN 2.36657
R17341 EN.n255 EN 2.36657
R17342 EN.n124 EN.n123 1.88889
R17343 EN.n151 EN.n150 1.88889
R17344 EN.n103 EN.n102 1.88889
R17345 EN.n54 EN.n53 1.83532
R17346 EN.n260 EN.n7 1.83532
R17347 EN.n140 EN.n139 1.80064
R17348 EN.n201 EN 1.7505
R17349 EN.n201 EN 1.7505
R17350 EN.n169 EN 1.7505
R17351 EN.n169 EN 1.7505
R17352 EN.n155 EN 1.7505
R17353 EN.n155 EN 1.7505
R17354 EN.n184 EN 1.7505
R17355 EN.n184 EN 1.7505
R17356 EN.n49 EN 1.73023
R17357 EN.n21 EN 1.73023
R17358 EN.n3 EN 1.73023
R17359 EN.n133 EN 1.52282
R17360 EN.n242 EN 1.52282
R17361 EN.n133 EN 1.42461
R17362 EN.n242 EN 1.42461
R17363 EN.n182 EN.n167 1.38649
R17364 EN.n124 EN 1.32983
R17365 EN.n151 EN 1.32983
R17366 EN.n103 EN 1.32983
R17367 EN.n54 EN 1.27213
R17368 EN EN.n260 1.27213
R17369 EN.n215 EN 1.26389
R17370 EN.n214 EN.n199 1.08292
R17371 EN.n235 EN.n226 1.08292
R17372 EN.n249 EN.n248 0.934566
R17373 EN.n258 EN.n249 0.738137
R17374 EN.n137 EN 0.666365
R17375 EN.n246 EN 0.666365
R17376 EN.n137 EN.n136 0.65675
R17377 EN.n246 EN.n245 0.65675
R17378 EN.n209 EN 0.580857
R17379 EN.n177 EN 0.580857
R17380 EN.n162 EN 0.580857
R17381 EN.n123 EN 0.580857
R17382 EN.n136 EN 0.580857
R17383 EN.n150 EN 0.580857
R17384 EN.n192 EN 0.580857
R17385 EN.n111 EN 0.580857
R17386 EN.n102 EN 0.580857
R17387 EN.n87 EN 0.580857
R17388 EN.n81 EN 0.580857
R17389 EN.n74 EN 0.580857
R17390 EN.n65 EN 0.580857
R17391 EN.n232 EN 0.580857
R17392 EN.n245 EN 0.580857
R17393 EN.n255 EN 0.580857
R17394 EN.n218 EN 0.527286
R17395 EN.n53 EN 0.527286
R17396 EN.n37 EN 0.527286
R17397 EN.n25 EN 0.527286
R17398 EN.n12 EN 0.527286
R17399 EN.n7 EN 0.527286
R17400 EN.n198 EN 0.442464
R17401 EN.n31 EN 0.418351
R17402 EN.n17 EN 0.418351
R17403 EN.n223 EN 0.371036
R17404 EN.n45 EN 0.246036
R17405 EN.n9 EN 0.246036
R17406 EN.n127 EN 0.24431
R17407 EN.n122 EN 0.225552
R17408 EN.n135 EN 0.225552
R17409 EN.n149 EN 0.225552
R17410 EN EN.n113 0.225552
R17411 EN.n101 EN 0.225552
R17412 EN.n86 EN 0.225552
R17413 EN EN.n83 0.225552
R17414 EN EN.n75 0.225552
R17415 EN EN.n66 0.225552
R17416 EN EN.n234 0.225552
R17417 EN.n244 EN 0.225552
R17418 EN EN.n257 0.225552
R17419 EN.n216 EN 0.196446
R17420 EN.n203 EN 0.196446
R17421 EN.n171 EN 0.196446
R17422 EN.n157 EN 0.196446
R17423 EN.n114 EN 0.196446
R17424 EN.n128 EN 0.196446
R17425 EN.n141 EN 0.196446
R17426 EN.n186 EN 0.196446
R17427 EN.n106 EN 0.196446
R17428 EN.n94 EN 0.196446
R17429 EN.n84 EN 0.196446
R17430 EN.n76 EN 0.196446
R17431 EN.n68 EN 0.196446
R17432 EN.n59 EN 0.196446
R17433 EN.n236 EN 0.196446
R17434 EN.n46 EN 0.196446
R17435 EN.n32 EN 0.196446
R17436 EN.n18 EN 0.196446
R17437 EN.n10 EN 0.196446
R17438 EN.n250 EN 0.196446
R17439 EN.n0 EN 0.196446
R17440 EN.n120 EN 0.192464
R17441 EN.n147 EN 0.192464
R17442 EN.n99 EN 0.192464
R17443 EN.n200 EN 0.17713
R17444 EN.n168 EN 0.17713
R17445 EN.n154 EN 0.17713
R17446 EN.n183 EN 0.17713
R17447 EN.n41 EN 0.15675
R17448 EN.n29 EN 0.15675
R17449 EN.n123 EN.n122 0.128681
R17450 EN.n136 EN.n135 0.128681
R17451 EN.n150 EN.n149 0.128681
R17452 EN.n113 EN.n111 0.128681
R17453 EN.n102 EN.n101 0.128681
R17454 EN.n87 EN.n86 0.128681
R17455 EN.n83 EN.n81 0.128681
R17456 EN.n75 EN.n74 0.128681
R17457 EN.n66 EN.n65 0.128681
R17458 EN.n234 EN.n232 0.128681
R17459 EN.n245 EN.n244 0.128681
R17460 EN.n257 EN.n255 0.128681
R17461 EN.n231 EN 0.10523
R17462 EN EN.n231 0.098473
R17463 EN.n210 EN.n200 0.0983261
R17464 EN.n178 EN.n168 0.0983261
R17465 EN.n163 EN.n154 0.0983261
R17466 EN.n193 EN.n183 0.0983261
R17467 EN.n41 EN.n40 0.0983261
R17468 EN.n29 EN.n28 0.0983261
R17469 EN.n231 EN.n227 0.0867069
R17470 EN.n222 EN.n216 0.0793043
R17471 EN EN.n222 0.0793043
R17472 EN.n210 EN.n209 0.0793043
R17473 EN.n178 EN.n177 0.0793043
R17474 EN.n163 EN.n162 0.0793043
R17475 EN.n193 EN.n192 0.0793043
R17476 EN.n93 EN 0.0793043
R17477 EN.n47 EN.n46 0.0793043
R17478 EN.n47 EN 0.0793043
R17479 EN.n33 EN.n32 0.0793043
R17480 EN.n33 EN 0.0793043
R17481 EN.n40 EN 0.0793043
R17482 EN.n19 EN.n18 0.0793043
R17483 EN.n19 EN 0.0793043
R17484 EN.n28 EN 0.0793043
R17485 EN.n13 EN.n10 0.0793043
R17486 EN.n13 EN 0.0793043
R17487 EN.n1 EN.n0 0.0793043
R17488 EN.n1 EN 0.0793043
R17489 EN.n213 EN.n200 0.0774231
R17490 EN.n181 EN.n168 0.0774231
R17491 EN.n166 EN.n154 0.0774231
R17492 EN.n125 EN.n120 0.0774231
R17493 EN.n125 EN.n124 0.0774231
R17494 EN.n138 EN.n133 0.0774231
R17495 EN.n138 EN.n137 0.0774231
R17496 EN.n152 EN.n147 0.0774231
R17497 EN.n152 EN.n151 0.0774231
R17498 EN.n196 EN.n183 0.0774231
R17499 EN.n104 EN.n99 0.0774231
R17500 EN.n104 EN.n103 0.0774231
R17501 EN.n247 EN.n242 0.0774231
R17502 EN.n247 EN.n246 0.0774231
R17503 EN.n55 EN.n45 0.0774231
R17504 EN.n55 EN.n54 0.0774231
R17505 EN.n42 EN.n41 0.0774231
R17506 EN.n30 EN.n29 0.0774231
R17507 EN.n259 EN.n9 0.0774231
R17508 EN.n260 EN.n259 0.0774231
R17509 EN.n212 EN.n201 0.0678077
R17510 EN.n180 EN.n169 0.0678077
R17511 EN.n165 EN.n155 0.0678077
R17512 EN.n195 EN.n184 0.0678077
R17513 EN.n227 EN 0.050069
R17514 EN.n219 EN.n218 0.03675
R17515 EN.n219 EN 0.03675
R17516 EN.n208 EN.n203 0.03675
R17517 EN EN.n208 0.03675
R17518 EN.n176 EN.n171 0.03675
R17519 EN EN.n176 0.03675
R17520 EN.n161 EN.n157 0.03675
R17521 EN EN.n161 0.03675
R17522 EN.n119 EN.n114 0.03675
R17523 EN EN.n119 0.03675
R17524 EN.n132 EN.n128 0.03675
R17525 EN EN.n132 0.03675
R17526 EN.n146 EN.n141 0.03675
R17527 EN EN.n146 0.03675
R17528 EN.n191 EN.n186 0.03675
R17529 EN EN.n191 0.03675
R17530 EN.n110 EN.n106 0.03675
R17531 EN EN.n110 0.03675
R17532 EN.n98 EN.n94 0.03675
R17533 EN EN.n98 0.03675
R17534 EN.n88 EN.n84 0.03675
R17535 EN.n88 EN 0.03675
R17536 EN.n80 EN.n76 0.03675
R17537 EN EN.n80 0.03675
R17538 EN.n73 EN.n68 0.03675
R17539 EN EN.n73 0.03675
R17540 EN.n64 EN.n59 0.03675
R17541 EN EN.n64 0.03675
R17542 EN.n241 EN.n236 0.03675
R17543 EN EN.n241 0.03675
R17544 EN.n53 EN.n52 0.03675
R17545 EN.n52 EN 0.03675
R17546 EN.n37 EN.n36 0.03675
R17547 EN.n36 EN 0.03675
R17548 EN.n25 EN.n24 0.03675
R17549 EN.n24 EN 0.03675
R17550 EN.n16 EN.n12 0.03675
R17551 EN EN.n16 0.03675
R17552 EN.n254 EN.n250 0.03675
R17553 EN EN.n254 0.03675
R17554 EN.n7 EN.n6 0.03675
R17555 EN.n6 EN 0.03675
R17556 EN.n213 EN.n212 0.0101154
R17557 EN.n181 EN.n180 0.0101154
R17558 EN.n166 EN.n165 0.0101154
R17559 EN.n196 EN.n195 0.0101154
R17560 EN.n42 EN.n31 0.0101154
R17561 EN.n30 EN.n17 0.0101154
R17562 EN EN.n216 0.00725676
R17563 EN EN.n203 0.00725676
R17564 EN EN.n171 0.00725676
R17565 EN EN.n157 0.00725676
R17566 EN EN.n114 0.00725676
R17567 EN EN.n128 0.00725676
R17568 EN EN.n141 0.00725676
R17569 EN EN.n186 0.00725676
R17570 EN EN.n106 0.00725676
R17571 EN EN.n94 0.00725676
R17572 EN.n84 EN 0.00725676
R17573 EN EN.n76 0.00725676
R17574 EN EN.n68 0.00725676
R17575 EN EN.n59 0.00725676
R17576 EN EN.n236 0.00725676
R17577 EN.n46 EN 0.00725676
R17578 EN.n32 EN 0.00725676
R17579 EN.n18 EN 0.00725676
R17580 EN EN.n10 0.00725676
R17581 EN EN.n250 0.00725676
R17582 EN.n0 EN 0.00725676
R17583 EN.n201 EN 0.00290385
R17584 EN.n169 EN 0.00290385
R17585 EN.n155 EN 0.00290385
R17586 EN.n184 EN 0.00290385
R17587 a_3210_10927.t0 a_3210_10927.t1 87.1434
R17588 a_4993_3829.n3 a_4993_3829.n2 647.119
R17589 a_4993_3829.n1 a_4993_3829.t4 350.253
R17590 a_4993_3829.n2 a_4993_3829.n0 260.339
R17591 a_4993_3829.n2 a_4993_3829.n1 246.119
R17592 a_4993_3829.n1 a_4993_3829.t5 189.588
R17593 a_4993_3829.n3 a_4993_3829.t1 89.1195
R17594 a_4993_3829.n0 a_4993_3829.t3 63.3338
R17595 a_4993_3829.t0 a_4993_3829.n3 41.0422
R17596 a_4993_3829.n0 a_4993_3829.t2 31.9797
R17597 a_4871_4233.t0 a_4871_4233.t1 198.571
R17598 a_5037_4221.t0 a_5037_4221.t1 60.0005
R17599 a_8008_10927.n3 a_8008_10927.n2 636.953
R17600 a_8008_10927.n1 a_8008_10927.t5 366.856
R17601 a_8008_10927.n2 a_8008_10927.n0 300.2
R17602 a_8008_10927.n2 a_8008_10927.n1 225.036
R17603 a_8008_10927.n1 a_8008_10927.t4 174.056
R17604 a_8008_10927.n0 a_8008_10927.t0 70.0005
R17605 a_8008_10927.n3 a_8008_10927.t3 68.0124
R17606 a_8008_10927.t1 a_8008_10927.n3 63.3219
R17607 a_8008_10927.n0 a_8008_10927.t2 61.6672
R17608 a_8183_10901.n3 a_8183_10901.n0 807.871
R17609 a_8183_10901.n4 a_8183_10901.t6 389.183
R17610 a_8183_10901.n5 a_8183_10901.n4 251.167
R17611 a_8183_10901.t0 a_8183_10901.n5 223.571
R17612 a_8183_10901.n1 a_8183_10901.t4 212.081
R17613 a_8183_10901.n2 a_8183_10901.t3 212.081
R17614 a_8183_10901.n3 a_8183_10901.n2 176.576
R17615 a_8183_10901.n4 a_8183_10901.t8 174.891
R17616 a_8183_10901.n1 a_8183_10901.t7 139.78
R17617 a_8183_10901.n2 a_8183_10901.t5 139.78
R17618 a_8183_10901.n0 a_8183_10901.t1 63.3219
R17619 a_8183_10901.n0 a_8183_10901.t2 63.3219
R17620 a_8183_10901.n2 a_8183_10901.n1 61.346
R17621 a_8183_10901.n5 a_8183_10901.n3 37.7195
R17622 CLK.n3 CLK.t6 184.768
R17623 CLK.n2 CLK.t1 184.768
R17624 CLK.n1 CLK.t0 184.768
R17625 CLK.n0 CLK.t7 184.768
R17626 CLK.n4 CLK.n3 171.375
R17627 CLK.n3 CLK.t2 146.208
R17628 CLK.n2 CLK.t5 146.208
R17629 CLK.n1 CLK.t4 146.208
R17630 CLK.n0 CLK.t3 146.208
R17631 CLK.n3 CLK.n2 40.6397
R17632 CLK.n2 CLK.n1 40.6397
R17633 CLK.n1 CLK.n0 40.6397
R17634 CLK CLK.n4 9.14336
R17635 CLK.n4 CLK 4.67352
R17636 a_6813_7093.n3 a_6813_7093.n2 330.051
R17637 a_6813_7093.n52 a_6813_7093.n51 327.253
R17638 a_6813_7093.n51 a_6813_7093.n0 217.256
R17639 a_6813_7093.n3 a_6813_7093.n1 217.256
R17640 a_6813_7093.n5 a_6813_7093.t35 212.081
R17641 a_6813_7093.n48 a_6813_7093.t31 212.081
R17642 a_6813_7093.n46 a_6813_7093.t28 212.081
R17643 a_6813_7093.n8 a_6813_7093.t24 212.081
R17644 a_6813_7093.n40 a_6813_7093.t20 212.081
R17645 a_6813_7093.n38 a_6813_7093.t29 212.081
R17646 a_6813_7093.n9 a_6813_7093.t25 212.081
R17647 a_6813_7093.n32 a_6813_7093.t22 212.081
R17648 a_6813_7093.n11 a_6813_7093.t10 212.081
R17649 a_6813_7093.n27 a_6813_7093.t9 212.081
R17650 a_6813_7093.n13 a_6813_7093.t15 212.081
R17651 a_6813_7093.n21 a_6813_7093.t12 212.081
R17652 a_6813_7093.n19 a_6813_7093.t19 212.081
R17653 a_6813_7093.n17 a_6813_7093.t38 212.081
R17654 a_6813_7093.n16 a_6813_7093.t34 212.081
R17655 a_6813_7093.n15 a_6813_7093.t33 212.081
R17656 a_6813_7093.n18 a_6813_7093.n14 169.409
R17657 a_6813_7093.n5 a_6813_7093.t27 162.274
R17658 a_6813_7093.n48 a_6813_7093.t21 162.274
R17659 a_6813_7093.n46 a_6813_7093.t17 162.274
R17660 a_6813_7093.n8 a_6813_7093.t14 162.274
R17661 a_6813_7093.n40 a_6813_7093.t11 162.274
R17662 a_6813_7093.n38 a_6813_7093.t18 162.274
R17663 a_6813_7093.n9 a_6813_7093.t16 162.274
R17664 a_6813_7093.n32 a_6813_7093.t13 162.274
R17665 a_6813_7093.n11 a_6813_7093.t36 162.274
R17666 a_6813_7093.n27 a_6813_7093.t32 162.274
R17667 a_6813_7093.n13 a_6813_7093.t39 162.274
R17668 a_6813_7093.n21 a_6813_7093.t37 162.274
R17669 a_6813_7093.n19 a_6813_7093.t8 162.274
R17670 a_6813_7093.n17 a_6813_7093.t30 162.274
R17671 a_6813_7093.n16 a_6813_7093.t26 162.274
R17672 a_6813_7093.n15 a_6813_7093.t23 162.274
R17673 a_6813_7093.n20 a_6813_7093.n14 152
R17674 a_6813_7093.n23 a_6813_7093.n22 152
R17675 a_6813_7093.n25 a_6813_7093.n24 152
R17676 a_6813_7093.n26 a_6813_7093.n12 152
R17677 a_6813_7093.n29 a_6813_7093.n28 152
R17678 a_6813_7093.n31 a_6813_7093.n30 152
R17679 a_6813_7093.n33 a_6813_7093.n10 152
R17680 a_6813_7093.n35 a_6813_7093.n34 152
R17681 a_6813_7093.n37 a_6813_7093.n36 152
R17682 a_6813_7093.n39 a_6813_7093.n7 152
R17683 a_6813_7093.n42 a_6813_7093.n41 152
R17684 a_6813_7093.n43 a_6813_7093.n6 152
R17685 a_6813_7093.n45 a_6813_7093.n44 152
R17686 a_6813_7093.n47 a_6813_7093.n4 152
R17687 a_6813_7093.n50 a_6813_7093.n49 152
R17688 a_6813_7093.n17 a_6813_7093.n16 55.2698
R17689 a_6813_7093.n16 a_6813_7093.n15 55.2698
R17690 a_6813_7093.n51 a_6813_7093.n3 44.0325
R17691 a_6813_7093.n45 a_6813_7093.n6 43.7018
R17692 a_6813_7093.n34 a_6813_7093.n33 43.7018
R17693 a_6813_7093.n26 a_6813_7093.n25 43.7018
R17694 a_6813_7093.n51 a_6813_7093.n50 43.5205
R17695 a_6813_7093.n22 a_6813_7093.n13 43.0592
R17696 a_6813_7093.n37 a_6813_7093.n9 42.4165
R17697 a_6813_7093.n0 a_6813_7093.t5 40.0005
R17698 a_6813_7093.n0 a_6813_7093.t6 40.0005
R17699 a_6813_7093.n1 a_6813_7093.t7 40.0005
R17700 a_6813_7093.n1 a_6813_7093.t4 40.0005
R17701 a_6813_7093.n47 a_6813_7093.n46 39.8458
R17702 a_6813_7093.n41 a_6813_7093.n8 35.9898
R17703 a_6813_7093.n18 a_6813_7093.n17 35.3472
R17704 a_6813_7093.n32 a_6813_7093.n31 33.4192
R17705 a_6813_7093.n28 a_6813_7093.n27 32.7765
R17706 a_6813_7093.n21 a_6813_7093.n20 31.4912
R17707 a_6813_7093.n39 a_6813_7093.n38 30.8485
R17708 a_6813_7093.n49 a_6813_7093.n48 28.2778
R17709 a_6813_7093.n2 a_6813_7093.t1 27.5805
R17710 a_6813_7093.n2 a_6813_7093.t2 27.5805
R17711 a_6813_7093.t3 a_6813_7093.n52 27.5805
R17712 a_6813_7093.n52 a_6813_7093.t0 27.5805
R17713 a_6813_7093.n49 a_6813_7093.n5 26.9925
R17714 a_6813_7093.n40 a_6813_7093.n39 24.4218
R17715 a_6813_7093.n20 a_6813_7093.n19 23.7792
R17716 a_6813_7093.n28 a_6813_7093.n11 22.4938
R17717 a_6813_7093.n31 a_6813_7093.n11 21.2085
R17718 a_6813_7093.n19 a_6813_7093.n18 19.9232
R17719 a_6813_7093.n41 a_6813_7093.n40 19.2805
R17720 a_6813_7093.n50 a_6813_7093.n4 17.4085
R17721 a_6813_7093.n44 a_6813_7093.n4 17.4085
R17722 a_6813_7093.n44 a_6813_7093.n43 17.4085
R17723 a_6813_7093.n43 a_6813_7093.n42 17.4085
R17724 a_6813_7093.n42 a_6813_7093.n7 17.4085
R17725 a_6813_7093.n36 a_6813_7093.n7 17.4085
R17726 a_6813_7093.n36 a_6813_7093.n35 17.4085
R17727 a_6813_7093.n35 a_6813_7093.n10 17.4085
R17728 a_6813_7093.n30 a_6813_7093.n10 17.4085
R17729 a_6813_7093.n30 a_6813_7093.n29 17.4085
R17730 a_6813_7093.n29 a_6813_7093.n12 17.4085
R17731 a_6813_7093.n24 a_6813_7093.n12 17.4085
R17732 a_6813_7093.n24 a_6813_7093.n23 17.4085
R17733 a_6813_7093.n23 a_6813_7093.n14 17.4085
R17734 a_6813_7093.n48 a_6813_7093.n47 15.4245
R17735 a_6813_7093.n38 a_6813_7093.n37 12.8538
R17736 a_6813_7093.n22 a_6813_7093.n21 12.2112
R17737 a_6813_7093.n27 a_6813_7093.n26 10.9258
R17738 a_6813_7093.n33 a_6813_7093.n32 10.2832
R17739 a_6813_7093.n8 a_6813_7093.n6 7.7125
R17740 a_6813_7093.n46 a_6813_7093.n45 3.8565
R17741 a_6813_7093.n34 a_6813_7093.n9 1.28583
R17742 a_6813_7093.n25 a_6813_7093.n13 0.643167
R17743 a_2584_6147.t0 a_2584_6147.n3 370.026
R17744 a_2584_6147.n0 a_2584_6147.t2 351.356
R17745 a_2584_6147.n1 a_2584_6147.t4 334.717
R17746 a_2584_6147.n3 a_2584_6147.t1 325.971
R17747 a_2584_6147.n1 a_2584_6147.t5 309.935
R17748 a_2584_6147.n0 a_2584_6147.t3 305.683
R17749 a_2584_6147.n2 a_2584_6147.n0 16.879
R17750 a_2584_6147.n3 a_2584_6147.n2 10.8867
R17751 a_2584_6147.n2 a_2584_6147.n1 9.3005
R17752 a_2306_6163.n3 a_2306_6163.n2 636.953
R17753 a_2306_6163.n1 a_2306_6163.t5 366.856
R17754 a_2306_6163.n2 a_2306_6163.n0 300.2
R17755 a_2306_6163.n2 a_2306_6163.n1 225.036
R17756 a_2306_6163.n1 a_2306_6163.t4 174.056
R17757 a_2306_6163.n0 a_2306_6163.t3 70.0005
R17758 a_2306_6163.t1 a_2306_6163.n3 68.0124
R17759 a_2306_6163.n3 a_2306_6163.t2 63.3219
R17760 a_2306_6163.n0 a_2306_6163.t0 61.6672
R17761 a_2710_6031.n3 a_2710_6031.n2 647.119
R17762 a_2710_6031.n1 a_2710_6031.t5 350.253
R17763 a_2710_6031.n2 a_2710_6031.n0 260.339
R17764 a_2710_6031.n2 a_2710_6031.n1 246.119
R17765 a_2710_6031.n1 a_2710_6031.t4 189.588
R17766 a_2710_6031.n3 a_2710_6031.t2 89.1195
R17767 a_2710_6031.n0 a_2710_6031.t3 63.3338
R17768 a_2710_6031.t0 a_2710_6031.n3 41.0422
R17769 a_2710_6031.n0 a_2710_6031.t1 31.9797
R17770 a_6942_6941.n3 a_6942_6941.n2 647.119
R17771 a_6942_6941.n1 a_6942_6941.t4 350.253
R17772 a_6942_6941.n2 a_6942_6941.n0 260.339
R17773 a_6942_6941.n2 a_6942_6941.n1 246.119
R17774 a_6942_6941.n1 a_6942_6941.t5 189.588
R17775 a_6942_6941.n3 a_6942_6941.t2 89.1195
R17776 a_6942_6941.n0 a_6942_6941.t3 63.3338
R17777 a_6942_6941.t0 a_6942_6941.n3 41.0422
R17778 a_6942_6941.n0 a_6942_6941.t1 31.9797
R17779 a_7249_6575.t0 a_7249_6575.t1 60.0005
R17780 a_7321_6575.t0 a_7321_6575.t1 198.571
R17781 a_10667_5247.n5 a_10667_5247.n4 807.871
R17782 a_10667_5247.n2 a_10667_5247.t5 389.183
R17783 a_10667_5247.n3 a_10667_5247.n2 251.167
R17784 a_10667_5247.n3 a_10667_5247.t1 223.571
R17785 a_10667_5247.n0 a_10667_5247.t7 212.081
R17786 a_10667_5247.n1 a_10667_5247.t3 212.081
R17787 a_10667_5247.n4 a_10667_5247.n1 176.576
R17788 a_10667_5247.n2 a_10667_5247.t4 174.891
R17789 a_10667_5247.n0 a_10667_5247.t6 139.78
R17790 a_10667_5247.n1 a_10667_5247.t8 139.78
R17791 a_10667_5247.n5 a_10667_5247.t2 63.3219
R17792 a_10667_5247.t0 a_10667_5247.n5 63.3219
R17793 a_10667_5247.n1 a_10667_5247.n0 61.346
R17794 a_10667_5247.n4 a_10667_5247.n3 37.7195
R17795 CF[6].n3 CF[6].n2 585
R17796 CF[6].n4 CF[6].n3 585
R17797 CF[6].n12 CF[6].t8 333.651
R17798 CF[6].n12 CF[6].t4 297.233
R17799 CF[6].n8 CF[6].t5 294.557
R17800 CF[6].n6 CF[6].t7 294.557
R17801 CF[6].n8 CF[6].t6 211.01
R17802 CF[6].n6 CF[6].t9 211.01
R17803 CF[6].n13 CF[6].n12 195.701
R17804 CF[6].n1 CF[6].n0 185
R17805 CF[6].n9 CF[6].n8 152
R17806 CF[6].n7 CF[6].n6 152
R17807 CF[6] CF[6].n1 57.7379
R17808 CF[6].n14 CF[6].n11 29.3082
R17809 CF[6].n11 CF[6].n10 27.9806
R17810 CF[6].n3 CF[6].t0 26.5955
R17811 CF[6].n3 CF[6].t1 26.5955
R17812 CF[6].n0 CF[6].t3 24.9236
R17813 CF[6].n0 CF[6].t2 24.9236
R17814 CF[6].n11 CF[6] 13.3525
R17815 CF[6].n15 CF[6].n14 11.2972
R17816 CF[6].n2 CF[6] 10.4965
R17817 CF[6].n4 CF[6] 10.4965
R17818 CF[6] CF[6].n7 10.4234
R17819 CF[6] CF[6].n5 9.4552
R17820 CF[6].n10 CF[6] 9.32621
R17821 CF[6].n14 CF[6].n13 9.3005
R17822 CF[6].n15 CF[6] 8.1504
R17823 CF[6].n2 CF[6] 6.9125
R17824 CF[6].n5 CF[6] 4.3525
R17825 CF[6] CF[6].n15 4.20667
R17826 CF[6].n5 CF[6].n4 2.5605
R17827 CF[6].n9 CF[6] 2.01193
R17828 CF[6].n7 CF[6] 2.01193
R17829 CF[6].n1 CF[6] 1.7925
R17830 CF[6].n10 CF[6].n9 1.09764
R17831 CF[6].n13 CF[6] 1.03669
R17832 a_8951_10927.n1 a_8951_10927.t2 530.01
R17833 a_8951_10927.t0 a_8951_10927.n5 421.021
R17834 a_8951_10927.n0 a_8951_10927.t3 337.142
R17835 a_8951_10927.n3 a_8951_10927.t1 280.223
R17836 a_8951_10927.n4 a_8951_10927.t7 263.173
R17837 a_8951_10927.n4 a_8951_10927.t6 227.826
R17838 a_8951_10927.n0 a_8951_10927.t4 199.762
R17839 a_8951_10927.n2 a_8951_10927.n1 170.81
R17840 a_8951_10927.n2 a_8951_10927.n0 167.321
R17841 a_8951_10927.n5 a_8951_10927.n4 152
R17842 a_8951_10927.n1 a_8951_10927.t5 141.923
R17843 a_8951_10927.n3 a_8951_10927.n2 10.8376
R17844 a_8951_10927.n5 a_8951_10927.n3 2.50485
R17845 a_2411_4917.n3 a_2411_4917.n2 674.338
R17846 a_2411_4917.n1 a_2411_4917.t5 332.58
R17847 a_2411_4917.n2 a_2411_4917.n0 284.012
R17848 a_2411_4917.n2 a_2411_4917.n1 253.648
R17849 a_2411_4917.n1 a_2411_4917.t4 168.701
R17850 a_2411_4917.n3 a_2411_4917.t3 96.1553
R17851 a_2411_4917.t1 a_2411_4917.n3 65.6672
R17852 a_2411_4917.n0 a_2411_4917.t2 65.0005
R17853 a_2411_4917.n0 a_2411_4917.t0 45.0005
R17854 a_2342_4943.n3 a_2342_4943.n2 647.119
R17855 a_2342_4943.n1 a_2342_4943.t4 350.253
R17856 a_2342_4943.n2 a_2342_4943.n0 260.339
R17857 a_2342_4943.n2 a_2342_4943.n1 246.119
R17858 a_2342_4943.n1 a_2342_4943.t5 189.588
R17859 a_2342_4943.n3 a_2342_4943.t3 89.1195
R17860 a_2342_4943.n0 a_2342_4943.t0 63.3338
R17861 a_2342_4943.t1 a_2342_4943.n3 41.0422
R17862 a_2342_4943.n0 a_2342_4943.t2 31.9797
R17863 COMP_N.n6 COMP_N.t5 235.763
R17864 COMP_N.n0 COMP_N.t2 221.72
R17865 COMP_N.n1 COMP_N.t4 221.72
R17866 COMP_N.n6 COMP_N.t1 163.464
R17867 COMP_N.n7 COMP_N.n6 152
R17868 COMP_N.n5 COMP_N.n4 152
R17869 COMP_N.n3 COMP_N.n2 152
R17870 COMP_N.n0 COMP_N.t3 149.421
R17871 COMP_N.n1 COMP_N.t0 149.421
R17872 COMP_N.n2 COMP_N.n1 58.019
R17873 COMP_N.n5 COMP_N.n0 43.7375
R17874 COMP_N.n4 COMP_N 20.8005
R17875 COMP_N.n8 COMP_N.n7 18.6384
R17876 COMP_N.n6 COMP_N.n5 17.8524
R17877 COMP_N.n2 COMP_N.n0 16.9598
R17878 COMP_N.n3 COMP_N 16.3205
R17879 COMP_N COMP_N.n3 13.1205
R17880 COMP_N.n4 COMP_N 8.6405
R17881 COMP_N COMP_N.n8 3.44845
R17882 COMP_N.n7 COMP_N 0.9605
R17883 a_7331_9269.n22 a_7331_9269.t4 286.348
R17884 a_7331_9269.n24 a_7331_9269.t0 271.051
R17885 a_7331_9269.n1 a_7331_9269.t16 221.72
R17886 a_7331_9269.n18 a_7331_9269.t10 221.72
R17887 a_7331_9269.n2 a_7331_9269.t6 221.72
R17888 a_7331_9269.n12 a_7331_9269.t12 221.72
R17889 a_7331_9269.n10 a_7331_9269.t8 221.72
R17890 a_7331_9269.n4 a_7331_9269.t14 221.72
R17891 a_7331_9269.n6 a_7331_9269.t20 221.72
R17892 a_7331_9269.n5 a_7331_9269.t15 221.72
R17893 a_7331_9269.n25 a_7331_9269.n24 206.055
R17894 a_7331_9269.n22 a_7331_9269.n21 198.177
R17895 a_7331_9269.n8 a_7331_9269.n7 177.601
R17896 a_7331_9269.n9 a_7331_9269.n8 152
R17897 a_7331_9269.n11 a_7331_9269.n3 152
R17898 a_7331_9269.n14 a_7331_9269.n13 152
R17899 a_7331_9269.n16 a_7331_9269.n15 152
R17900 a_7331_9269.n17 a_7331_9269.n0 152
R17901 a_7331_9269.n20 a_7331_9269.n19 152
R17902 a_7331_9269.n1 a_7331_9269.t7 149.421
R17903 a_7331_9269.n18 a_7331_9269.t17 149.421
R17904 a_7331_9269.n2 a_7331_9269.t11 149.421
R17905 a_7331_9269.n12 a_7331_9269.t18 149.421
R17906 a_7331_9269.n10 a_7331_9269.t13 149.421
R17907 a_7331_9269.n4 a_7331_9269.t19 149.421
R17908 a_7331_9269.n6 a_7331_9269.t9 149.421
R17909 a_7331_9269.n5 a_7331_9269.t21 149.421
R17910 a_7331_9269.n6 a_7331_9269.n5 74.9783
R17911 a_7331_9269.n7 a_7331_9269.n6 66.0523
R17912 a_7331_9269.n17 a_7331_9269.n16 60.6968
R17913 a_7331_9269.n19 a_7331_9269.n18 55.3412
R17914 a_7331_9269.n13 a_7331_9269.n2 51.7709
R17915 a_7331_9269.n9 a_7331_9269.n4 51.7709
R17916 a_7331_9269.n23 a_7331_9269.n22 48.9632
R17917 a_7331_9269.n24 a_7331_9269.n23 38.7339
R17918 a_7331_9269.n12 a_7331_9269.n11 37.4894
R17919 a_7331_9269.n11 a_7331_9269.n10 37.4894
R17920 a_7331_9269.t2 a_7331_9269.n25 26.5955
R17921 a_7331_9269.n25 a_7331_9269.t1 26.5955
R17922 a_7331_9269.n20 a_7331_9269.n0 25.6005
R17923 a_7331_9269.n15 a_7331_9269.n0 25.6005
R17924 a_7331_9269.n15 a_7331_9269.n14 25.6005
R17925 a_7331_9269.n14 a_7331_9269.n3 25.6005
R17926 a_7331_9269.n8 a_7331_9269.n3 25.6005
R17927 a_7331_9269.n21 a_7331_9269.t3 24.9236
R17928 a_7331_9269.n21 a_7331_9269.t5 24.9236
R17929 a_7331_9269.n13 a_7331_9269.n12 23.2079
R17930 a_7331_9269.n10 a_7331_9269.n9 23.2079
R17931 a_7331_9269.n19 a_7331_9269.n1 19.6375
R17932 a_7331_9269.n23 a_7331_9269.n20 18.4476
R17933 a_7331_9269.n16 a_7331_9269.n2 8.92643
R17934 a_7331_9269.n7 a_7331_9269.n4 8.92643
R17935 a_7331_9269.n18 a_7331_9269.n17 5.35606
R17936 a_4424_4667.t0 a_4424_4667.n3 370.026
R17937 a_4424_4667.n0 a_4424_4667.t4 351.356
R17938 a_4424_4667.n1 a_4424_4667.t2 334.717
R17939 a_4424_4667.n3 a_4424_4667.t1 325.971
R17940 a_4424_4667.n1 a_4424_4667.t5 309.935
R17941 a_4424_4667.n0 a_4424_4667.t3 305.683
R17942 a_4424_4667.n2 a_4424_4667.n0 16.879
R17943 a_4424_4667.n3 a_4424_4667.n2 10.8867
R17944 a_4424_4667.n2 a_4424_4667.n1 9.3005
R17945 a_4929_4399.t1 a_4929_4399.t0 198.571
R17946 a_4619_4636.n3 a_4619_4636.n2 674.338
R17947 a_4619_4636.n1 a_4619_4636.t4 332.58
R17948 a_4619_4636.n2 a_4619_4636.n0 284.012
R17949 a_4619_4636.n2 a_4619_4636.n1 253.648
R17950 a_4619_4636.n1 a_4619_4636.t5 168.701
R17951 a_4619_4636.n3 a_4619_4636.t2 96.1553
R17952 a_4619_4636.t1 a_4619_4636.n3 65.6672
R17953 a_4619_4636.n0 a_4619_4636.t3 65.0005
R17954 a_4619_4636.n0 a_4619_4636.t0 45.0005
R17955 CF[4].n11 CF[4].t7 333.651
R17956 CF[4].n11 CF[4].t9 297.233
R17957 CF[4].n5 CF[4].t6 294.557
R17958 CF[4].n8 CF[4].t4 294.557
R17959 CF[4].n1 CF[4].n0 289.096
R17960 CF[4].n5 CF[4].t8 211.01
R17961 CF[4].n8 CF[4].t5 211.01
R17962 CF[4].n12 CF[4].n11 195.701
R17963 CF[4].n3 CF[4].n2 185
R17964 CF[4].n9 CF[4].n8 153.097
R17965 CF[4].n6 CF[4].n5 152
R17966 CF[4].n3 CF[4] 49.0339
R17967 CF[4] CF[4].n7 40.9598
R17968 CF[4].n0 CF[4].t1 26.5955
R17969 CF[4].n0 CF[4].t3 26.5955
R17970 CF[4].n2 CF[4].t2 24.9236
R17971 CF[4].n2 CF[4].t0 24.9236
R17972 CF[4].n13 CF[4].n10 16.1557
R17973 CF[4].n14 CF[4].n4 15.4901
R17974 CF[4].n14 CF[4].n13 11.366
R17975 CF[4] CF[4].n1 9.48653
R17976 CF[4].n7 CF[4] 9.32621
R17977 CF[4].n13 CF[4].n12 9.3005
R17978 CF[4].n10 CF[4].n9 9.3005
R17979 CF[4].n1 CF[4] 7.7181
R17980 CF[4].n4 CF[4].n3 6.1445
R17981 CF[4] CF[4].n14 4.66911
R17982 CF[4].n4 CF[4] 4.3525
R17983 CF[4].n9 CF[4] 3.10907
R17984 CF[4].n6 CF[4] 2.01193
R17985 CF[4].n7 CF[4].n6 1.09764
R17986 CF[4].n12 CF[4] 1.03669
R17987 CF[4].n10 CF[4] 0.0991761
R17988 a_5015_3009.n1 a_5015_3009.t3 530.01
R17989 a_5015_3009.t0 a_5015_3009.n5 421.021
R17990 a_5015_3009.n0 a_5015_3009.t4 337.171
R17991 a_5015_3009.n3 a_5015_3009.t1 280.223
R17992 a_5015_3009.n4 a_5015_3009.t5 263.173
R17993 a_5015_3009.n4 a_5015_3009.t7 227.826
R17994 a_5015_3009.n0 a_5015_3009.t6 199.762
R17995 a_5015_3009.n2 a_5015_3009.n1 170.81
R17996 a_5015_3009.n2 a_5015_3009.n0 167.321
R17997 a_5015_3009.n5 a_5015_3009.n4 152
R17998 a_5015_3009.n1 a_5015_3009.t2 141.923
R17999 a_5015_3009.n3 a_5015_3009.n2 10.8376
R18000 a_5015_3009.n5 a_5015_3009.n3 2.50485
R18001 a_4463_4541.n1 a_4463_4541.t7 530.01
R18002 a_4463_4541.t0 a_4463_4541.n5 421.021
R18003 a_4463_4541.n0 a_4463_4541.t5 337.171
R18004 a_4463_4541.n3 a_4463_4541.t1 280.223
R18005 a_4463_4541.n4 a_4463_4541.t2 263.173
R18006 a_4463_4541.n4 a_4463_4541.t4 227.826
R18007 a_4463_4541.n0 a_4463_4541.t3 199.762
R18008 a_4463_4541.n2 a_4463_4541.n1 170.81
R18009 a_4463_4541.n2 a_4463_4541.n0 167.321
R18010 a_4463_4541.n5 a_4463_4541.n4 152
R18011 a_4463_4541.n1 a_4463_4541.t6 141.923
R18012 a_4463_4541.n3 a_4463_4541.n2 10.8376
R18013 a_4463_4541.n5 a_4463_4541.n3 2.50485
R18014 a_10207_10901.n5 a_10207_10901.n4 807.871
R18015 a_10207_10901.n2 a_10207_10901.t3 389.183
R18016 a_10207_10901.n3 a_10207_10901.n2 251.167
R18017 a_10207_10901.n3 a_10207_10901.t1 223.571
R18018 a_10207_10901.n0 a_10207_10901.t6 212.081
R18019 a_10207_10901.n1 a_10207_10901.t5 212.081
R18020 a_10207_10901.n4 a_10207_10901.n1 176.576
R18021 a_10207_10901.n2 a_10207_10901.t7 174.891
R18022 a_10207_10901.n0 a_10207_10901.t4 139.78
R18023 a_10207_10901.n1 a_10207_10901.t8 139.78
R18024 a_10207_10901.t0 a_10207_10901.n5 63.3219
R18025 a_10207_10901.n5 a_10207_10901.t2 63.3219
R18026 a_10207_10901.n1 a_10207_10901.n0 61.346
R18027 a_10207_10901.n4 a_10207_10901.n3 37.7195
R18028 a_10194_11293.t0 a_10194_11293.t1 126.644
R18029 a_6538_6827.n3 a_6538_6827.n2 636.953
R18030 a_6538_6827.n1 a_6538_6827.t5 366.856
R18031 a_6538_6827.n2 a_6538_6827.n0 300.2
R18032 a_6538_6827.n2 a_6538_6827.n1 225.036
R18033 a_6538_6827.n1 a_6538_6827.t4 174.056
R18034 a_6538_6827.n0 a_6538_6827.t3 70.0005
R18035 a_6538_6827.t1 a_6538_6827.n3 68.0124
R18036 a_6538_6827.n3 a_6538_6827.t2 63.3219
R18037 a_6538_6827.n0 a_6538_6827.t0 61.6672
R18038 a_6251_6549.n5 a_6251_6549.n4 807.871
R18039 a_6251_6549.n0 a_6251_6549.t5 389.183
R18040 a_6251_6549.n1 a_6251_6549.n0 251.167
R18041 a_6251_6549.n1 a_6251_6549.t1 223.571
R18042 a_6251_6549.n3 a_6251_6549.t3 212.081
R18043 a_6251_6549.n2 a_6251_6549.t8 212.081
R18044 a_6251_6549.n4 a_6251_6549.n3 176.576
R18045 a_6251_6549.n0 a_6251_6549.t7 174.891
R18046 a_6251_6549.n3 a_6251_6549.t6 139.78
R18047 a_6251_6549.n2 a_6251_6549.t4 139.78
R18048 a_6251_6549.t0 a_6251_6549.n5 63.3219
R18049 a_6251_6549.n5 a_6251_6549.t2 63.3219
R18050 a_6251_6549.n3 a_6251_6549.n2 61.346
R18051 a_6251_6549.n4 a_6251_6549.n1 37.5061
R18052 a_4424_6843.t0 a_4424_6843.n3 370.026
R18053 a_4424_6843.n0 a_4424_6843.t3 351.356
R18054 a_4424_6843.n1 a_4424_6843.t5 334.717
R18055 a_4424_6843.n3 a_4424_6843.t1 325.971
R18056 a_4424_6843.n1 a_4424_6843.t4 309.935
R18057 a_4424_6843.n0 a_4424_6843.t2 305.683
R18058 a_4424_6843.n2 a_4424_6843.n0 16.879
R18059 a_4424_6843.n3 a_4424_6843.n2 10.8867
R18060 a_4424_6843.n2 a_4424_6843.n1 9.3005
R18061 a_4380_6941.t0 a_4380_6941.t1 126.644
R18062 a_4146_6827.n3 a_4146_6827.n2 636.953
R18063 a_4146_6827.n1 a_4146_6827.t5 366.856
R18064 a_4146_6827.n2 a_4146_6827.n0 300.2
R18065 a_4146_6827.n2 a_4146_6827.n1 225.036
R18066 a_4146_6827.n1 a_4146_6827.t4 174.056
R18067 a_4146_6827.n0 a_4146_6827.t0 70.0005
R18068 a_4146_6827.n3 a_4146_6827.t2 68.0124
R18069 a_4146_6827.t1 a_4146_6827.n3 63.3219
R18070 a_4146_6827.n0 a_4146_6827.t3 61.6672
R18071 a_2526_4765.n3 a_2526_4765.n2 647.119
R18072 a_2526_4765.n1 a_2526_4765.t4 350.253
R18073 a_2526_4765.n2 a_2526_4765.n0 260.339
R18074 a_2526_4765.n2 a_2526_4765.n1 246.119
R18075 a_2526_4765.n1 a_2526_4765.t5 189.588
R18076 a_2526_4765.n3 a_2526_4765.t3 89.1195
R18077 a_2526_4765.n0 a_2526_4765.t0 63.3338
R18078 a_2526_4765.t2 a_2526_4765.n3 41.0422
R18079 a_2526_4765.n0 a_2526_4765.t1 31.9797
R18080 a_2833_4399.t0 a_2833_4399.t1 60.0005
R18081 a_2905_4399.t0 a_2905_4399.t1 198.571
R18082 CF[8].n3 CF[8].n2 585
R18083 CF[8].n4 CF[8].n3 585
R18084 CF[8].n11 CF[8].t8 333.651
R18085 CF[8].n11 CF[8].t6 297.233
R18086 CF[8].n8 CF[8].t7 294.557
R18087 CF[8].n6 CF[8].t9 294.557
R18088 CF[8].n8 CF[8].t4 211.01
R18089 CF[8].n6 CF[8].t5 211.01
R18090 CF[8].n12 CF[8].n11 195.701
R18091 CF[8].n1 CF[8].n0 185
R18092 CF[8] CF[8].n8 156.207
R18093 CF[8].n7 CF[8].n6 153.097
R18094 CF[8] CF[8].n1 57.7379
R18095 CF[8].n13 CF[8].n10 27.4732
R18096 CF[8].n3 CF[8].t2 26.5955
R18097 CF[8].n3 CF[8].t3 26.5955
R18098 CF[8].n0 CF[8].t0 24.9236
R18099 CF[8].n0 CF[8].t1 24.9236
R18100 CF[8].n10 CF[8].n7 22.5987
R18101 CF[8].n10 CF[8].n9 19.6865
R18102 CF[8].n14 CF[8].n13 11.366
R18103 CF[8].n2 CF[8] 10.4965
R18104 CF[8].n4 CF[8] 10.4965
R18105 CF[8] CF[8].n5 9.66056
R18106 CF[8].n9 CF[8] 9.32621
R18107 CF[8].n13 CF[8].n12 9.3005
R18108 CF[8].n2 CF[8] 6.9125
R18109 CF[8].n14 CF[8] 6.23127
R18110 CF[8] CF[8].n14 4.90062
R18111 CF[8].n5 CF[8] 4.3525
R18112 CF[8].n9 CF[8] 3.10907
R18113 CF[8].n7 CF[8] 3.10907
R18114 CF[8].n5 CF[8].n4 2.5605
R18115 CF[8].n1 CF[8] 1.7925
R18116 CF[8].n12 CF[8] 1.03669
R18117 a_2623_6273.n1 a_2623_6273.t6 530.01
R18118 a_2623_6273.t0 a_2623_6273.n5 421.021
R18119 a_2623_6273.n0 a_2623_6273.t5 337.171
R18120 a_2623_6273.n3 a_2623_6273.t1 280.223
R18121 a_2623_6273.n4 a_2623_6273.t4 263.173
R18122 a_2623_6273.n4 a_2623_6273.t7 227.826
R18123 a_2623_6273.n0 a_2623_6273.t3 199.762
R18124 a_2623_6273.n2 a_2623_6273.n1 170.81
R18125 a_2623_6273.n2 a_2623_6273.n0 167.321
R18126 a_2623_6273.n5 a_2623_6273.n4 152
R18127 a_2623_6273.n1 a_2623_6273.t2 141.923
R18128 a_2623_6273.n3 a_2623_6273.n2 10.8376
R18129 a_2623_6273.n5 a_2623_6273.n3 2.50485
R18130 a_3031_10901.n5 a_3031_10901.n4 807.871
R18131 a_3031_10901.n2 a_3031_10901.t5 389.183
R18132 a_3031_10901.n3 a_3031_10901.n2 251.167
R18133 a_3031_10901.n3 a_3031_10901.t1 223.571
R18134 a_3031_10901.n0 a_3031_10901.t8 212.081
R18135 a_3031_10901.n1 a_3031_10901.t4 212.081
R18136 a_3031_10901.n4 a_3031_10901.n1 176.576
R18137 a_3031_10901.n2 a_3031_10901.t3 174.891
R18138 a_3031_10901.n0 a_3031_10901.t6 139.78
R18139 a_3031_10901.n1 a_3031_10901.t7 139.78
R18140 a_3031_10901.t0 a_3031_10901.n5 63.3219
R18141 a_3031_10901.n5 a_3031_10901.t2 63.3219
R18142 a_3031_10901.n1 a_3031_10901.n0 61.346
R18143 a_3031_10901.n4 a_3031_10901.n3 37.7195
R18144 a_2965_10927.t1 a_2965_10927.t0 94.7268
R18145 a_6375_8213.n1 a_6375_8213.t7 530.01
R18146 a_6375_8213.t1 a_6375_8213.n5 421.021
R18147 a_6375_8213.n0 a_6375_8213.t4 337.142
R18148 a_6375_8213.n3 a_6375_8213.t0 280.223
R18149 a_6375_8213.n4 a_6375_8213.t5 263.173
R18150 a_6375_8213.n4 a_6375_8213.t2 227.826
R18151 a_6375_8213.n0 a_6375_8213.t6 199.762
R18152 a_6375_8213.n2 a_6375_8213.n1 170.81
R18153 a_6375_8213.n2 a_6375_8213.n0 167.321
R18154 a_6375_8213.n5 a_6375_8213.n4 152
R18155 a_6375_8213.n1 a_6375_8213.t3 141.923
R18156 a_6375_8213.n3 a_6375_8213.n2 10.8376
R18157 a_6375_8213.n5 a_6375_8213.n3 2.50485
R18158 a_6541_8213.t0 a_6541_8213.n3 370.026
R18159 a_6541_8213.n0 a_6541_8213.t5 351.356
R18160 a_6541_8213.n1 a_6541_8213.t4 334.717
R18161 a_6541_8213.n3 a_6541_8213.t1 325.971
R18162 a_6541_8213.n1 a_6541_8213.t2 309.935
R18163 a_6541_8213.n0 a_6541_8213.t3 305.683
R18164 a_6541_8213.n2 a_6541_8213.n0 16.879
R18165 a_6541_8213.n3 a_6541_8213.n2 10.8867
R18166 a_6541_8213.n2 a_6541_8213.n1 9.3005
R18167 a_10943_6549.n5 a_10943_6549.n4 807.871
R18168 a_10943_6549.n2 a_10943_6549.t6 389.183
R18169 a_10943_6549.n3 a_10943_6549.n2 251.167
R18170 a_10943_6549.n3 a_10943_6549.t2 223.571
R18171 a_10943_6549.n0 a_10943_6549.t3 212.081
R18172 a_10943_6549.n1 a_10943_6549.t7 212.081
R18173 a_10943_6549.n4 a_10943_6549.n1 176.576
R18174 a_10943_6549.n2 a_10943_6549.t8 174.891
R18175 a_10943_6549.n0 a_10943_6549.t5 139.78
R18176 a_10943_6549.n1 a_10943_6549.t4 139.78
R18177 a_10943_6549.n5 a_10943_6549.t1 63.3219
R18178 a_10943_6549.t0 a_10943_6549.n5 63.3219
R18179 a_10943_6549.n1 a_10943_6549.n0 61.346
R18180 a_10943_6549.n4 a_10943_6549.n3 37.7195
R18181 CF[9].n0 CF[9] 586.793
R18182 CF[9].n1 CF[9].n0 585
R18183 CF[9].n10 CF[9].t6 333.651
R18184 CF[9].n10 CF[9].t9 297.233
R18185 CF[9].n7 CF[9].t4 294.557
R18186 CF[9].n5 CF[9].t5 294.557
R18187 CF[9].n7 CF[9].t8 211.01
R18188 CF[9].n5 CF[9].t7 211.01
R18189 CF[9].n11 CF[9].n10 195.701
R18190 CF[9].n3 CF[9].n2 185
R18191 CF[9].n6 CF[9].n5 153.097
R18192 CF[9].n8 CF[9].n7 152
R18193 CF[9].n3 CF[9] 49.0339
R18194 CF[9].n0 CF[9].t1 26.5955
R18195 CF[9].n0 CF[9].t0 26.5955
R18196 CF[9].n2 CF[9].t2 24.9236
R18197 CF[9].n2 CF[9].t3 24.9236
R18198 CF[9].n9 CF[9].n6 21.3199
R18199 CF[9].n12 CF[9].n9 20.502
R18200 CF[9].n9 CF[9] 16.9091
R18201 CF[9].n1 CF[9] 15.6165
R18202 CF[9] CF[9].n4 14.7212
R18203 CF[9].n13 CF[9].n12 11.7768
R18204 CF[9] CF[9].n8 10.4234
R18205 CF[9].n12 CF[9].n11 9.3005
R18206 CF[9].n4 CF[9].n3 6.1445
R18207 CF[9].n4 CF[9] 4.3525
R18208 CF[9] CF[9].n13 4.06253
R18209 CF[9].n6 CF[9] 3.10907
R18210 CF[9].n8 CF[9] 2.01193
R18211 CF[9] CF[9].n1 1.7925
R18212 CF[9].n11 CF[9] 1.03669
R18213 CF[9].n13 CF[9] 0.768872
R18214 a_1835_4373.n5 a_1835_4373.n4 807.871
R18215 a_1835_4373.n0 a_1835_4373.t7 389.183
R18216 a_1835_4373.n1 a_1835_4373.n0 251.167
R18217 a_1835_4373.n1 a_1835_4373.t2 223.571
R18218 a_1835_4373.n3 a_1835_4373.t4 212.081
R18219 a_1835_4373.n2 a_1835_4373.t8 212.081
R18220 a_1835_4373.n4 a_1835_4373.n3 176.576
R18221 a_1835_4373.n0 a_1835_4373.t3 174.891
R18222 a_1835_4373.n3 a_1835_4373.t6 139.78
R18223 a_1835_4373.n2 a_1835_4373.t5 139.78
R18224 a_1835_4373.t0 a_1835_4373.n5 63.3219
R18225 a_1835_4373.n5 a_1835_4373.t1 63.3219
R18226 a_1835_4373.n3 a_1835_4373.n2 61.346
R18227 a_1835_4373.n4 a_1835_4373.n1 37.5061
R18228 a_2397_4399.n0 a_2397_4399.t1 68.3338
R18229 a_2397_4399.n0 a_2397_4399.t0 26.3935
R18230 a_2397_4399.n1 a_2397_4399.n0 14.4005
R18231 clknet_0_CLK.n31 clknet_0_CLK.n29 333.392
R18232 clknet_0_CLK.n31 clknet_0_CLK.n30 301.392
R18233 clknet_0_CLK.n33 clknet_0_CLK.n32 301.392
R18234 clknet_0_CLK.n35 clknet_0_CLK.n34 301.392
R18235 clknet_0_CLK.n39 clknet_0_CLK.n27 301.392
R18236 clknet_0_CLK.n38 clknet_0_CLK.n28 301.392
R18237 clknet_0_CLK.n37 clknet_0_CLK.n36 301.392
R18238 clknet_0_CLK clknet_0_CLK.n40 297.752
R18239 clknet_0_CLK.n2 clknet_0_CLK.n0 248.638
R18240 clknet_0_CLK.n2 clknet_0_CLK.n1 203.463
R18241 clknet_0_CLK.n4 clknet_0_CLK.n3 203.463
R18242 clknet_0_CLK.n8 clknet_0_CLK.n7 203.463
R18243 clknet_0_CLK.n24 clknet_0_CLK.n23 203.463
R18244 clknet_0_CLK.n6 clknet_0_CLK.n5 202.456
R18245 clknet_0_CLK.n26 clknet_0_CLK.n25 200.212
R18246 clknet_0_CLK.n21 clknet_0_CLK.n9 188.201
R18247 clknet_0_CLK.n13 clknet_0_CLK.t40 184.768
R18248 clknet_0_CLK.n12 clknet_0_CLK.t33 184.768
R18249 clknet_0_CLK.n11 clknet_0_CLK.t45 184.768
R18250 clknet_0_CLK.n10 clknet_0_CLK.t34 184.768
R18251 clknet_0_CLK.n15 clknet_0_CLK.t39 184.768
R18252 clknet_0_CLK.n16 clknet_0_CLK.t37 184.768
R18253 clknet_0_CLK.n17 clknet_0_CLK.t36 184.768
R18254 clknet_0_CLK.n18 clknet_0_CLK.t35 184.768
R18255 clknet_0_CLK clknet_0_CLK.n13 173.609
R18256 clknet_0_CLK.n19 clknet_0_CLK.n18 171.375
R18257 clknet_0_CLK.n13 clknet_0_CLK.t47 146.208
R18258 clknet_0_CLK.n12 clknet_0_CLK.t46 146.208
R18259 clknet_0_CLK.n11 clknet_0_CLK.t44 146.208
R18260 clknet_0_CLK.n10 clknet_0_CLK.t32 146.208
R18261 clknet_0_CLK.n15 clknet_0_CLK.t43 146.208
R18262 clknet_0_CLK.n16 clknet_0_CLK.t42 146.208
R18263 clknet_0_CLK.n17 clknet_0_CLK.t41 146.208
R18264 clknet_0_CLK.n18 clknet_0_CLK.t38 146.208
R18265 clknet_0_CLK.n4 clknet_0_CLK.n2 45.177
R18266 clknet_0_CLK.n22 clknet_0_CLK.n8 45.177
R18267 clknet_0_CLK.n24 clknet_0_CLK.n22 45.177
R18268 clknet_0_CLK.n6 clknet_0_CLK.n4 44.0476
R18269 clknet_0_CLK.n8 clknet_0_CLK.n6 44.0476
R18270 clknet_0_CLK.n13 clknet_0_CLK.n12 40.6397
R18271 clknet_0_CLK.n12 clknet_0_CLK.n11 40.6397
R18272 clknet_0_CLK.n11 clknet_0_CLK.n10 40.6397
R18273 clknet_0_CLK.n16 clknet_0_CLK.n15 40.6397
R18274 clknet_0_CLK.n17 clknet_0_CLK.n16 40.6397
R18275 clknet_0_CLK.n18 clknet_0_CLK.n17 40.6397
R18276 clknet_0_CLK.n0 clknet_0_CLK.t21 40.0005
R18277 clknet_0_CLK.n0 clknet_0_CLK.t24 40.0005
R18278 clknet_0_CLK.n1 clknet_0_CLK.t26 40.0005
R18279 clknet_0_CLK.n1 clknet_0_CLK.t28 40.0005
R18280 clknet_0_CLK.n3 clknet_0_CLK.t30 40.0005
R18281 clknet_0_CLK.n3 clknet_0_CLK.t25 40.0005
R18282 clknet_0_CLK.n5 clknet_0_CLK.t27 40.0005
R18283 clknet_0_CLK.n5 clknet_0_CLK.t29 40.0005
R18284 clknet_0_CLK.n7 clknet_0_CLK.t18 40.0005
R18285 clknet_0_CLK.n7 clknet_0_CLK.t19 40.0005
R18286 clknet_0_CLK.n9 clknet_0_CLK.t16 40.0005
R18287 clknet_0_CLK.n9 clknet_0_CLK.t17 40.0005
R18288 clknet_0_CLK.n23 clknet_0_CLK.t31 40.0005
R18289 clknet_0_CLK.n23 clknet_0_CLK.t20 40.0005
R18290 clknet_0_CLK.n25 clknet_0_CLK.t22 40.0005
R18291 clknet_0_CLK.n25 clknet_0_CLK.t23 40.0005
R18292 clknet_0_CLK.n33 clknet_0_CLK.n31 32.0005
R18293 clknet_0_CLK.n35 clknet_0_CLK.n33 32.0005
R18294 clknet_0_CLK.n39 clknet_0_CLK.n38 32.0005
R18295 clknet_0_CLK.n38 clknet_0_CLK.n37 32.0005
R18296 clknet_0_CLK.n37 clknet_0_CLK.n35 31.2005
R18297 clknet_0_CLK.n20 clknet_0_CLK 28.256
R18298 clknet_0_CLK.n29 clknet_0_CLK.t1 27.5805
R18299 clknet_0_CLK.n29 clknet_0_CLK.t4 27.5805
R18300 clknet_0_CLK.n30 clknet_0_CLK.t6 27.5805
R18301 clknet_0_CLK.n30 clknet_0_CLK.t8 27.5805
R18302 clknet_0_CLK.n32 clknet_0_CLK.t10 27.5805
R18303 clknet_0_CLK.n32 clknet_0_CLK.t5 27.5805
R18304 clknet_0_CLK.n34 clknet_0_CLK.t7 27.5805
R18305 clknet_0_CLK.n34 clknet_0_CLK.t9 27.5805
R18306 clknet_0_CLK.n27 clknet_0_CLK.t11 27.5805
R18307 clknet_0_CLK.n27 clknet_0_CLK.t0 27.5805
R18308 clknet_0_CLK.n40 clknet_0_CLK.t2 27.5805
R18309 clknet_0_CLK.n40 clknet_0_CLK.t3 27.5805
R18310 clknet_0_CLK.n28 clknet_0_CLK.t12 27.5805
R18311 clknet_0_CLK.n28 clknet_0_CLK.t13 27.5805
R18312 clknet_0_CLK.n36 clknet_0_CLK.t14 27.5805
R18313 clknet_0_CLK.n36 clknet_0_CLK.t15 27.5805
R18314 clknet_0_CLK.n20 clknet_0_CLK.n14 26.5342
R18315 clknet_0_CLK.n22 clknet_0_CLK.n21 15.262
R18316 clknet_0_CLK.n26 clknet_0_CLK.n24 13.177
R18317 clknet_0_CLK.n14 clknet_0_CLK 10.3624
R18318 clknet_0_CLK clknet_0_CLK.n39 10.2022
R18319 clknet_0_CLK.n21 clknet_0_CLK 9.4552
R18320 clknet_0_CLK clknet_0_CLK.n19 9.14336
R18321 clknet_0_CLK.n19 clknet_0_CLK 4.67352
R18322 clknet_0_CLK clknet_0_CLK.n20 4.63992
R18323 clknet_0_CLK.n14 clknet_0_CLK 3.45447
R18324 clknet_0_CLK clknet_0_CLK.n26 1.26402
R18325 a_5055_3285.n3 a_5055_3285.n0 807.871
R18326 a_5055_3285.n4 a_5055_3285.t3 389.183
R18327 a_5055_3285.n5 a_5055_3285.n4 251.167
R18328 a_5055_3285.t0 a_5055_3285.n5 223.571
R18329 a_5055_3285.n2 a_5055_3285.t5 212.081
R18330 a_5055_3285.n1 a_5055_3285.t8 212.081
R18331 a_5055_3285.n3 a_5055_3285.n2 176.576
R18332 a_5055_3285.n4 a_5055_3285.t7 174.891
R18333 a_5055_3285.n2 a_5055_3285.t6 139.78
R18334 a_5055_3285.n1 a_5055_3285.t4 139.78
R18335 a_5055_3285.n0 a_5055_3285.t2 63.3219
R18336 a_5055_3285.n0 a_5055_3285.t1 63.3219
R18337 a_5055_3285.n2 a_5055_3285.n1 61.346
R18338 a_5055_3285.n5 a_5055_3285.n3 37.5061
R18339 a_5576_3677.t0 a_5576_3677.t1 126.644
R18340 CF[2].n9 CF[2].n8 585
R18341 CF[2].n8 CF[2].n7 585
R18342 CF[2].n5 CF[2].t8 332.312
R18343 CF[2].n5 CF[2].t7 295.627
R18344 CF[2].n2 CF[2].t4 294.557
R18345 CF[2].n0 CF[2].t6 294.557
R18346 CF[2].n2 CF[2].t5 211.01
R18347 CF[2].n0 CF[2].t9 211.01
R18348 CF[2] CF[2].n5 196.004
R18349 CF[2].n11 CF[2].n10 185
R18350 CF[2] CF[2].n0 156.207
R18351 CF[2].n3 CF[2].n2 152
R18352 CF[2].n11 CF[2] 57.7379
R18353 CF[2].n8 CF[2].t2 26.5955
R18354 CF[2].n8 CF[2].t0 26.5955
R18355 CF[2].n10 CF[2].t1 24.9236
R18356 CF[2].n10 CF[2].t3 24.9236
R18357 CF[2].n4 CF[2].n1 22.9985
R18358 CF[2].n12 CF[2] 18.4466
R18359 CF[2].n4 CF[2] 16.9091
R18360 CF[2].n6 CF[2] 16.0868
R18361 CF[2] CF[2].n12 13.1329
R18362 CF[2] CF[2].n9 10.4965
R18363 CF[2].n7 CF[2] 10.4965
R18364 CF[2] CF[2].n3 10.4234
R18365 CF[2].n1 CF[2] 9.32621
R18366 CF[2].n9 CF[2] 6.9125
R18367 CF[2].n7 CF[2] 6.9125
R18368 CF[2].n6 CF[2].n4 4.11863
R18369 CF[2].n1 CF[2] 3.10907
R18370 CF[2].n12 CF[2].n6 2.2972
R18371 CF[2].n3 CF[2] 2.01193
R18372 CF[2] CF[2].n11 1.7925
R18373 a_6743_4399.n1 a_6743_4399.t6 530.01
R18374 a_6743_4399.t0 a_6743_4399.n5 421.021
R18375 a_6743_4399.n0 a_6743_4399.t2 337.142
R18376 a_6743_4399.n3 a_6743_4399.t1 280.223
R18377 a_6743_4399.n4 a_6743_4399.t3 263.173
R18378 a_6743_4399.n4 a_6743_4399.t5 227.826
R18379 a_6743_4399.n0 a_6743_4399.t7 199.762
R18380 a_6743_4399.n2 a_6743_4399.n1 170.81
R18381 a_6743_4399.n2 a_6743_4399.n0 167.321
R18382 a_6743_4399.n5 a_6743_4399.n4 152
R18383 a_6743_4399.n1 a_6743_4399.t4 141.923
R18384 a_6743_4399.n3 a_6743_4399.n2 10.8376
R18385 a_6743_4399.n5 a_6743_4399.n3 2.50485
R18386 a_4972_12015.n3 a_4972_12015.n2 636.953
R18387 a_4972_12015.n1 a_4972_12015.t4 366.856
R18388 a_4972_12015.n2 a_4972_12015.n0 300.2
R18389 a_4972_12015.n2 a_4972_12015.n1 225.036
R18390 a_4972_12015.n1 a_4972_12015.t5 174.056
R18391 a_4972_12015.n0 a_4972_12015.t1 70.0005
R18392 a_4972_12015.t2 a_4972_12015.n3 68.0124
R18393 a_4972_12015.n3 a_4972_12015.t3 63.3219
R18394 a_4972_12015.n0 a_4972_12015.t0 61.6672
R18395 a_5326_12015.t0 a_5326_12015.t1 87.1434
R18396 a_5147_11989.n5 a_5147_11989.n4 807.871
R18397 a_5147_11989.n2 a_5147_11989.t6 389.183
R18398 a_5147_11989.n3 a_5147_11989.n2 251.167
R18399 a_5147_11989.n3 a_5147_11989.t1 223.571
R18400 a_5147_11989.n0 a_5147_11989.t3 212.081
R18401 a_5147_11989.n1 a_5147_11989.t8 212.081
R18402 a_5147_11989.n4 a_5147_11989.n1 176.576
R18403 a_5147_11989.n2 a_5147_11989.t4 174.891
R18404 a_5147_11989.n0 a_5147_11989.t7 139.78
R18405 a_5147_11989.n1 a_5147_11989.t5 139.78
R18406 a_5147_11989.n5 a_5147_11989.t2 63.3219
R18407 a_5147_11989.t0 a_5147_11989.n5 63.3219
R18408 a_5147_11989.n1 a_5147_11989.n0 61.346
R18409 a_5147_11989.n4 a_5147_11989.n3 37.7195
R18410 a_4421_4399.n0 a_4421_4399.t0 68.3338
R18411 a_4421_4399.n0 a_4421_4399.t1 26.3935
R18412 a_4421_4399.n1 a_4421_4399.n0 14.4005
R18413 a_4146_4651.n3 a_4146_4651.n2 636.953
R18414 a_4146_4651.n1 a_4146_4651.t4 366.856
R18415 a_4146_4651.n2 a_4146_4651.n0 300.2
R18416 a_4146_4651.n2 a_4146_4651.n1 225.036
R18417 a_4146_4651.n1 a_4146_4651.t5 174.056
R18418 a_4146_4651.n0 a_4146_4651.t2 70.0005
R18419 a_4146_4651.t1 a_4146_4651.n3 68.0124
R18420 a_4146_4651.n3 a_4146_4651.t3 63.3219
R18421 a_4146_4651.n0 a_4146_4651.t0 61.6672
R18422 a_3583_4917.n5 a_3583_4917.n4 807.871
R18423 a_3583_4917.n0 a_3583_4917.t7 389.183
R18424 a_3583_4917.n1 a_3583_4917.n0 251.167
R18425 a_3583_4917.n1 a_3583_4917.t1 223.571
R18426 a_3583_4917.n3 a_3583_4917.t8 212.081
R18427 a_3583_4917.n2 a_3583_4917.t6 212.081
R18428 a_3583_4917.n4 a_3583_4917.n3 176.576
R18429 a_3583_4917.n0 a_3583_4917.t4 174.891
R18430 a_3583_4917.n3 a_3583_4917.t5 139.78
R18431 a_3583_4917.n2 a_3583_4917.t3 139.78
R18432 a_3583_4917.t0 a_3583_4917.n5 63.3219
R18433 a_3583_4917.n5 a_3583_4917.t2 63.3219
R18434 a_3583_4917.n3 a_3583_4917.n2 61.346
R18435 a_3583_4917.n4 a_3583_4917.n1 37.5061
R18436 SWN[9].n2 SWN[9].n1 585
R18437 SWN[9].n1 SWN[9].n0 585
R18438 SWN[9].n4 SWN[9].n3 185
R18439 SWN[9].n4 SWN[9] 57.7379
R18440 SWN[9].n1 SWN[9].t0 26.5955
R18441 SWN[9].n1 SWN[9].t1 26.5955
R18442 SWN[9].n3 SWN[9].t2 24.9236
R18443 SWN[9].n3 SWN[9].t3 24.9236
R18444 SWN[9] SWN[9].n2 10.4965
R18445 SWN[9].n0 SWN[9] 10.4965
R18446 SWN[9].n2 SWN[9] 6.9125
R18447 SWN[9].n0 SWN[9] 6.9125
R18448 SWN[9] SWN[9].n4 1.7925
R18449 a_8638_4221.t0 a_8638_4221.t1 87.1434
R18450 a_10759_6335.n5 a_10759_6335.n4 807.871
R18451 a_10759_6335.n2 a_10759_6335.t4 389.183
R18452 a_10759_6335.n3 a_10759_6335.n2 251.167
R18453 a_10759_6335.n3 a_10759_6335.t1 223.571
R18454 a_10759_6335.n0 a_10759_6335.t7 212.081
R18455 a_10759_6335.n1 a_10759_6335.t8 212.081
R18456 a_10759_6335.n4 a_10759_6335.n1 176.576
R18457 a_10759_6335.n2 a_10759_6335.t3 174.891
R18458 a_10759_6335.n0 a_10759_6335.t5 139.78
R18459 a_10759_6335.n1 a_10759_6335.t6 139.78
R18460 a_10759_6335.n5 a_10759_6335.t2 63.3219
R18461 a_10759_6335.t0 a_10759_6335.n5 63.3219
R18462 a_10759_6335.n1 a_10759_6335.n0 61.346
R18463 a_10759_6335.n4 a_10759_6335.n3 37.7195
R18464 a_4371_8449.n1 a_4371_8449.t2 530.01
R18465 a_4371_8449.t1 a_4371_8449.n5 421.021
R18466 a_4371_8449.n0 a_4371_8449.t5 337.171
R18467 a_4371_8449.n3 a_4371_8449.t0 280.223
R18468 a_4371_8449.n4 a_4371_8449.t7 263.173
R18469 a_4371_8449.n4 a_4371_8449.t4 227.826
R18470 a_4371_8449.n0 a_4371_8449.t6 199.762
R18471 a_4371_8449.n2 a_4371_8449.n1 170.81
R18472 a_4371_8449.n2 a_4371_8449.n0 167.321
R18473 a_4371_8449.n5 a_4371_8449.n4 152
R18474 a_4371_8449.n1 a_4371_8449.t3 141.923
R18475 a_4371_8449.n3 a_4371_8449.n2 10.8376
R18476 a_4371_8449.n5 a_4371_8449.n3 2.50485
R18477 a_4672_8207.t0 a_4672_8207.n0 1327.82
R18478 a_4672_8207.n0 a_4672_8207.t1 194.655
R18479 a_4672_8207.n0 a_4672_8207.t2 63.3219
R18480 a_4527_8181.n3 a_4527_8181.n2 674.338
R18481 a_4527_8181.n1 a_4527_8181.t5 332.58
R18482 a_4527_8181.n2 a_4527_8181.n0 284.012
R18483 a_4527_8181.n2 a_4527_8181.n1 253.648
R18484 a_4527_8181.n1 a_4527_8181.t4 168.701
R18485 a_4527_8181.t0 a_4527_8181.n3 96.1553
R18486 a_4527_8181.n3 a_4527_8181.t2 65.6672
R18487 a_4527_8181.n0 a_4527_8181.t1 65.0005
R18488 a_4527_8181.n0 a_4527_8181.t3 45.0005
R18489 x2/net11.n6 x2/net11.n5 585
R18490 x2/net11.n5 x2/net11.n4 585
R18491 x2/net11.n2 x2/net11.t4 230.576
R18492 x2/net11.n1 x2/net11.n0 185
R18493 x2/net11.n2 x2/net11.t5 158.275
R18494 x2/net11.n3 x2/net11.n2 153.165
R18495 x2/net11 x2/net11.n1 49.0339
R18496 x2/net11.n4 x2/net11 39.7024
R18497 x2/net11.n5 x2/net11.t0 26.5955
R18498 x2/net11.n5 x2/net11.t1 26.5955
R18499 x2/net11.n0 x2/net11.t3 24.9236
R18500 x2/net11.n0 x2/net11.t2 24.9236
R18501 x2/net11.n6 x2/net11 15.6165
R18502 x2/net11.n1 x2/net11 10.4965
R18503 x2/net11 x2/net11.n3 10.1739
R18504 x2/net11.n3 x2/net11 3.29747
R18505 x2/net11.n4 x2/net11 1.7925
R18506 x2/net11 x2/net11.n6 1.7925
R18507 clknet_1_0__leaf_CLK.n52 clknet_1_0__leaf_CLK.n50 333.392
R18508 clknet_1_0__leaf_CLK.n58 clknet_1_0__leaf_CLK.n48 301.392
R18509 clknet_1_0__leaf_CLK.n57 clknet_1_0__leaf_CLK.n49 301.392
R18510 clknet_1_0__leaf_CLK.n52 clknet_1_0__leaf_CLK.n51 301.392
R18511 clknet_1_0__leaf_CLK.n54 clknet_1_0__leaf_CLK.n53 301.392
R18512 clknet_1_0__leaf_CLK.n56 clknet_1_0__leaf_CLK.n55 301.392
R18513 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n60 297.752
R18514 clknet_1_0__leaf_CLK.n26 clknet_1_0__leaf_CLK.t37 294.557
R18515 clknet_1_0__leaf_CLK.n23 clknet_1_0__leaf_CLK.t44 294.557
R18516 clknet_1_0__leaf_CLK.n21 clknet_1_0__leaf_CLK.t40 294.557
R18517 clknet_1_0__leaf_CLK.n41 clknet_1_0__leaf_CLK.t38 294.557
R18518 clknet_1_0__leaf_CLK.n36 clknet_1_0__leaf_CLK.t45 294.557
R18519 clknet_1_0__leaf_CLK.n34 clknet_1_0__leaf_CLK.t55 294.557
R18520 clknet_1_0__leaf_CLK.n32 clknet_1_0__leaf_CLK.t50 294.557
R18521 clknet_1_0__leaf_CLK.n30 clknet_1_0__leaf_CLK.t49 294.557
R18522 clknet_1_0__leaf_CLK.n28 clknet_1_0__leaf_CLK.t46 294.557
R18523 clknet_1_0__leaf_CLK.n16 clknet_1_0__leaf_CLK.t47 294.557
R18524 clknet_1_0__leaf_CLK.n47 clknet_1_0__leaf_CLK.n46 287.303
R18525 clknet_1_0__leaf_CLK.n4 clknet_1_0__leaf_CLK.n2 248.638
R18526 clknet_1_0__leaf_CLK.n26 clknet_1_0__leaf_CLK.t43 211.01
R18527 clknet_1_0__leaf_CLK.n23 clknet_1_0__leaf_CLK.t54 211.01
R18528 clknet_1_0__leaf_CLK.n21 clknet_1_0__leaf_CLK.t41 211.01
R18529 clknet_1_0__leaf_CLK.n41 clknet_1_0__leaf_CLK.t42 211.01
R18530 clknet_1_0__leaf_CLK.n36 clknet_1_0__leaf_CLK.t52 211.01
R18531 clknet_1_0__leaf_CLK.n34 clknet_1_0__leaf_CLK.t35 211.01
R18532 clknet_1_0__leaf_CLK.n32 clknet_1_0__leaf_CLK.t34 211.01
R18533 clknet_1_0__leaf_CLK.n30 clknet_1_0__leaf_CLK.t33 211.01
R18534 clknet_1_0__leaf_CLK.n28 clknet_1_0__leaf_CLK.t32 211.01
R18535 clknet_1_0__leaf_CLK.n16 clknet_1_0__leaf_CLK.t53 211.01
R18536 clknet_1_0__leaf_CLK.n4 clknet_1_0__leaf_CLK.n3 203.463
R18537 clknet_1_0__leaf_CLK.n6 clknet_1_0__leaf_CLK.n5 203.463
R18538 clknet_1_0__leaf_CLK.n10 clknet_1_0__leaf_CLK.n9 203.463
R18539 clknet_1_0__leaf_CLK.n12 clknet_1_0__leaf_CLK.n11 203.463
R18540 clknet_1_0__leaf_CLK.n14 clknet_1_0__leaf_CLK.n13 203.463
R18541 clknet_1_0__leaf_CLK.n8 clknet_1_0__leaf_CLK.n7 202.456
R18542 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n15 200.212
R18543 clknet_1_0__leaf_CLK.n19 clknet_1_0__leaf_CLK.t39 184.768
R18544 clknet_1_0__leaf_CLK.n18 clknet_1_0__leaf_CLK.t36 184.768
R18545 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n19 173.609
R18546 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n23 156.207
R18547 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n41 156.207
R18548 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n16 156.207
R18549 clknet_1_0__leaf_CLK.n37 clknet_1_0__leaf_CLK.n36 153.097
R18550 clknet_1_0__leaf_CLK.n35 clknet_1_0__leaf_CLK.n34 153.097
R18551 clknet_1_0__leaf_CLK.n0 clknet_1_0__leaf_CLK.n26 152
R18552 clknet_1_0__leaf_CLK.n1 clknet_1_0__leaf_CLK.n21 152
R18553 clknet_1_0__leaf_CLK.n33 clknet_1_0__leaf_CLK.n32 152
R18554 clknet_1_0__leaf_CLK.n31 clknet_1_0__leaf_CLK.n30 152
R18555 clknet_1_0__leaf_CLK.n29 clknet_1_0__leaf_CLK.n28 152
R18556 clknet_1_0__leaf_CLK.n19 clknet_1_0__leaf_CLK.t51 146.208
R18557 clknet_1_0__leaf_CLK.n18 clknet_1_0__leaf_CLK.t48 146.208
R18558 clknet_1_0__leaf_CLK.n6 clknet_1_0__leaf_CLK.n4 45.177
R18559 clknet_1_0__leaf_CLK.n12 clknet_1_0__leaf_CLK.n10 45.177
R18560 clknet_1_0__leaf_CLK.n14 clknet_1_0__leaf_CLK.n12 45.177
R18561 clknet_1_0__leaf_CLK.n8 clknet_1_0__leaf_CLK.n6 44.0476
R18562 clknet_1_0__leaf_CLK.n10 clknet_1_0__leaf_CLK.n8 44.0476
R18563 clknet_1_0__leaf_CLK.n19 clknet_1_0__leaf_CLK.n18 40.6397
R18564 clknet_1_0__leaf_CLK.n2 clknet_1_0__leaf_CLK.t4 40.0005
R18565 clknet_1_0__leaf_CLK.n2 clknet_1_0__leaf_CLK.t18 40.0005
R18566 clknet_1_0__leaf_CLK.n3 clknet_1_0__leaf_CLK.t16 40.0005
R18567 clknet_1_0__leaf_CLK.n3 clknet_1_0__leaf_CLK.t23 40.0005
R18568 clknet_1_0__leaf_CLK.n5 clknet_1_0__leaf_CLK.t30 40.0005
R18569 clknet_1_0__leaf_CLK.n5 clknet_1_0__leaf_CLK.t2 40.0005
R18570 clknet_1_0__leaf_CLK.n7 clknet_1_0__leaf_CLK.t28 40.0005
R18571 clknet_1_0__leaf_CLK.n7 clknet_1_0__leaf_CLK.t25 40.0005
R18572 clknet_1_0__leaf_CLK.n9 clknet_1_0__leaf_CLK.t9 40.0005
R18573 clknet_1_0__leaf_CLK.n9 clknet_1_0__leaf_CLK.t6 40.0005
R18574 clknet_1_0__leaf_CLK.n11 clknet_1_0__leaf_CLK.t5 40.0005
R18575 clknet_1_0__leaf_CLK.n11 clknet_1_0__leaf_CLK.t27 40.0005
R18576 clknet_1_0__leaf_CLK.n13 clknet_1_0__leaf_CLK.t22 40.0005
R18577 clknet_1_0__leaf_CLK.n13 clknet_1_0__leaf_CLK.t7 40.0005
R18578 clknet_1_0__leaf_CLK.n15 clknet_1_0__leaf_CLK.t20 40.0005
R18579 clknet_1_0__leaf_CLK.n15 clknet_1_0__leaf_CLK.t14 40.0005
R18580 clknet_1_0__leaf_CLK.n59 clknet_1_0__leaf_CLK.n58 32.0005
R18581 clknet_1_0__leaf_CLK.n58 clknet_1_0__leaf_CLK.n57 32.0005
R18582 clknet_1_0__leaf_CLK.n54 clknet_1_0__leaf_CLK.n52 32.0005
R18583 clknet_1_0__leaf_CLK.n56 clknet_1_0__leaf_CLK.n54 32.0005
R18584 clknet_1_0__leaf_CLK.n57 clknet_1_0__leaf_CLK.n56 31.2005
R18585 clknet_1_0__leaf_CLK.n46 clknet_1_0__leaf_CLK.t17 27.5805
R18586 clknet_1_0__leaf_CLK.n46 clknet_1_0__leaf_CLK.t24 27.5805
R18587 clknet_1_0__leaf_CLK.n60 clknet_1_0__leaf_CLK.t10 27.5805
R18588 clknet_1_0__leaf_CLK.n60 clknet_1_0__leaf_CLK.t19 27.5805
R18589 clknet_1_0__leaf_CLK.n48 clknet_1_0__leaf_CLK.t29 27.5805
R18590 clknet_1_0__leaf_CLK.n48 clknet_1_0__leaf_CLK.t1 27.5805
R18591 clknet_1_0__leaf_CLK.n49 clknet_1_0__leaf_CLK.t26 27.5805
R18592 clknet_1_0__leaf_CLK.n49 clknet_1_0__leaf_CLK.t31 27.5805
R18593 clknet_1_0__leaf_CLK.n50 clknet_1_0__leaf_CLK.t12 27.5805
R18594 clknet_1_0__leaf_CLK.n50 clknet_1_0__leaf_CLK.t8 27.5805
R18595 clknet_1_0__leaf_CLK.n51 clknet_1_0__leaf_CLK.t21 27.5805
R18596 clknet_1_0__leaf_CLK.n51 clknet_1_0__leaf_CLK.t15 27.5805
R18597 clknet_1_0__leaf_CLK.n53 clknet_1_0__leaf_CLK.t13 27.5805
R18598 clknet_1_0__leaf_CLK.n53 clknet_1_0__leaf_CLK.t11 27.5805
R18599 clknet_1_0__leaf_CLK.n55 clknet_1_0__leaf_CLK.t3 27.5805
R18600 clknet_1_0__leaf_CLK.n55 clknet_1_0__leaf_CLK.t0 27.5805
R18601 clknet_1_0__leaf_CLK.n47 clknet_1_0__leaf_CLK.n45 25.7205
R18602 clknet_1_0__leaf_CLK.n22 clknet_1_0__leaf_CLK.n20 21.3913
R18603 clknet_1_0__leaf_CLK.n22 clknet_1_0__leaf_CLK.n1 14.5053
R18604 clknet_1_0__leaf_CLK.n27 clknet_1_0__leaf_CLK.n0 14.0946
R18605 clknet_1_0__leaf_CLK.n59 clknet_1_0__leaf_CLK.n47 14.0898
R18606 clknet_1_0__leaf_CLK.n25 clknet_1_0__leaf_CLK.n24 13.8005
R18607 clknet_1_0__leaf_CLK.n43 clknet_1_0__leaf_CLK.n42 13.8005
R18608 clknet_1_0__leaf_CLK.n38 clknet_1_0__leaf_CLK.n35 13.291
R18609 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n14 13.177
R18610 clknet_1_0__leaf_CLK.n40 clknet_1_0__leaf_CLK 12.7032
R18611 clknet_1_0__leaf_CLK.n39 clknet_1_0__leaf_CLK.n38 11.2972
R18612 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n33 10.4234
R18613 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n31 10.4234
R18614 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n29 10.4234
R18615 clknet_1_0__leaf_CLK.n20 clknet_1_0__leaf_CLK 10.3624
R18616 clknet_1_0__leaf_CLK clknet_1_0__leaf_CLK.n59 10.2022
R18617 clknet_1_0__leaf_CLK.n45 clknet_1_0__leaf_CLK.n17 9.79203
R18618 clknet_1_0__leaf_CLK.n0 clknet_1_0__leaf_CLK 9.32621
R18619 clknet_1_0__leaf_CLK.n24 clknet_1_0__leaf_CLK 9.32621
R18620 clknet_1_0__leaf_CLK.n1 clknet_1_0__leaf_CLK 9.32621
R18621 clknet_1_0__leaf_CLK.n42 clknet_1_0__leaf_CLK 9.32621
R18622 clknet_1_0__leaf_CLK.n17 clknet_1_0__leaf_CLK 9.32621
R18623 clknet_1_0__leaf_CLK.n38 clknet_1_0__leaf_CLK.n37 9.3005
R18624 clknet_1_0__leaf_CLK.n39 clknet_1_0__leaf_CLK 7.43146
R18625 clknet_1_0__leaf_CLK.n43 clknet_1_0__leaf_CLK.n40 6.49363
R18626 clknet_1_0__leaf_CLK.n45 clknet_1_0__leaf_CLK.n44 4.84528
R18627 clknet_1_0__leaf_CLK.n44 clknet_1_0__leaf_CLK.n43 4.11863
R18628 clknet_1_0__leaf_CLK.n40 clknet_1_0__leaf_CLK.n39 3.97577
R18629 clknet_1_0__leaf_CLK.n20 clknet_1_0__leaf_CLK 3.45447
R18630 clknet_1_0__leaf_CLK.n24 clknet_1_0__leaf_CLK 3.10907
R18631 clknet_1_0__leaf_CLK.n42 clknet_1_0__leaf_CLK 3.10907
R18632 clknet_1_0__leaf_CLK.n37 clknet_1_0__leaf_CLK 3.10907
R18633 clknet_1_0__leaf_CLK.n35 clknet_1_0__leaf_CLK 3.10907
R18634 clknet_1_0__leaf_CLK.n17 clknet_1_0__leaf_CLK 3.10907
R18635 clknet_1_0__leaf_CLK.n1 clknet_1_0__leaf_CLK 3.10907
R18636 clknet_1_0__leaf_CLK.n0 clknet_1_0__leaf_CLK 3.10907
R18637 clknet_1_0__leaf_CLK.n44 clknet_1_0__leaf_CLK.n27 2.90435
R18638 clknet_1_0__leaf_CLK.n25 clknet_1_0__leaf_CLK.n22 2.2972
R18639 clknet_1_0__leaf_CLK.n27 clknet_1_0__leaf_CLK.n25 2.2972
R18640 clknet_1_0__leaf_CLK.n33 clknet_1_0__leaf_CLK 2.01193
R18641 clknet_1_0__leaf_CLK.n31 clknet_1_0__leaf_CLK 2.01193
R18642 clknet_1_0__leaf_CLK.n29 clknet_1_0__leaf_CLK 2.01193
R18643 a_9595_3311.n1 a_9595_3311.t3 530.01
R18644 a_9595_3311.t0 a_9595_3311.n5 421.021
R18645 a_9595_3311.n0 a_9595_3311.t4 337.142
R18646 a_9595_3311.n3 a_9595_3311.t1 280.223
R18647 a_9595_3311.n4 a_9595_3311.t2 263.173
R18648 a_9595_3311.n4 a_9595_3311.t6 227.826
R18649 a_9595_3311.n0 a_9595_3311.t7 199.762
R18650 a_9595_3311.n2 a_9595_3311.n1 170.81
R18651 a_9595_3311.n2 a_9595_3311.n0 167.321
R18652 a_9595_3311.n5 a_9595_3311.n4 152
R18653 a_9595_3311.n1 a_9595_3311.t5 141.923
R18654 a_9595_3311.n3 a_9595_3311.n2 10.8376
R18655 a_9595_3311.n5 a_9595_3311.n3 2.50485
R18656 a_9853_6575.t0 a_9853_6575.n3 370.026
R18657 a_9853_6575.n0 a_9853_6575.t3 351.356
R18658 a_9853_6575.n1 a_9853_6575.t4 334.717
R18659 a_9853_6575.n3 a_9853_6575.t1 325.971
R18660 a_9853_6575.n1 a_9853_6575.t2 309.935
R18661 a_9853_6575.n0 a_9853_6575.t5 305.683
R18662 a_9853_6575.n2 a_9853_6575.n0 16.879
R18663 a_9853_6575.n3 a_9853_6575.n2 10.8867
R18664 a_9853_6575.n2 a_9853_6575.n1 9.3005
R18665 a_10108_6575.n1 a_10108_6575.n0 926.024
R18666 a_10108_6575.t0 a_10108_6575.n1 82.0838
R18667 a_10108_6575.n0 a_10108_6575.t1 63.3338
R18668 a_10108_6575.n1 a_10108_6575.t2 63.3219
R18669 a_10108_6575.n0 a_10108_6575.t3 29.7268
R18670 a_10203_6575.n3 a_10203_6575.n2 674.338
R18671 a_10203_6575.n1 a_10203_6575.t5 332.58
R18672 a_10203_6575.n2 a_10203_6575.n0 284.012
R18673 a_10203_6575.n2 a_10203_6575.n1 253.648
R18674 a_10203_6575.n1 a_10203_6575.t4 168.701
R18675 a_10203_6575.n3 a_10203_6575.t2 96.1553
R18676 a_10203_6575.t1 a_10203_6575.n3 65.6672
R18677 a_10203_6575.n0 a_10203_6575.t3 65.0005
R18678 a_10203_6575.n0 a_10203_6575.t0 45.0005
R18679 a_10299_7423.n4 a_10299_7423.n1 807.871
R18680 a_10299_7423.n0 a_10299_7423.t5 389.183
R18681 a_10299_7423.n5 a_10299_7423.n0 251.167
R18682 a_10299_7423.t0 a_10299_7423.n5 223.571
R18683 a_10299_7423.n2 a_10299_7423.t3 212.081
R18684 a_10299_7423.n3 a_10299_7423.t7 212.081
R18685 a_10299_7423.n4 a_10299_7423.n3 176.576
R18686 a_10299_7423.n0 a_10299_7423.t6 174.891
R18687 a_10299_7423.n2 a_10299_7423.t8 139.78
R18688 a_10299_7423.n3 a_10299_7423.t4 139.78
R18689 a_10299_7423.n1 a_10299_7423.t1 63.3219
R18690 a_10299_7423.n1 a_10299_7423.t2 63.3219
R18691 a_10299_7423.n3 a_10299_7423.n2 61.346
R18692 a_10299_7423.n5 a_10299_7423.n4 37.7195
R18693 a_7407_3009.n1 a_7407_3009.t4 530.01
R18694 a_7407_3009.t0 a_7407_3009.n5 421.021
R18695 a_7407_3009.n0 a_7407_3009.t2 337.171
R18696 a_7407_3009.n3 a_7407_3009.t1 280.223
R18697 a_7407_3009.n4 a_7407_3009.t5 263.173
R18698 a_7407_3009.n4 a_7407_3009.t6 227.826
R18699 a_7407_3009.n0 a_7407_3009.t7 199.762
R18700 a_7407_3009.n2 a_7407_3009.n1 170.81
R18701 a_7407_3009.n2 a_7407_3009.n0 167.321
R18702 a_7407_3009.n5 a_7407_3009.n4 152
R18703 a_7407_3009.n1 a_7407_3009.t3 141.923
R18704 a_7407_3009.n3 a_7407_3009.n2 10.8376
R18705 a_7407_3009.n5 a_7407_3009.n3 2.50485
R18706 a_7090_2899.n3 a_7090_2899.n2 636.953
R18707 a_7090_2899.n1 a_7090_2899.t5 366.856
R18708 a_7090_2899.n2 a_7090_2899.n0 300.2
R18709 a_7090_2899.n2 a_7090_2899.n1 225.036
R18710 a_7090_2899.n1 a_7090_2899.t4 174.056
R18711 a_7090_2899.n0 a_7090_2899.t1 70.0005
R18712 a_7090_2899.n3 a_7090_2899.t3 68.0124
R18713 a_7090_2899.t0 a_7090_2899.n3 63.3219
R18714 a_7090_2899.n0 a_7090_2899.t2 61.6672
R18715 a_7494_2767.n3 a_7494_2767.n2 647.119
R18716 a_7494_2767.n1 a_7494_2767.t4 350.253
R18717 a_7494_2767.n2 a_7494_2767.n0 260.339
R18718 a_7494_2767.n2 a_7494_2767.n1 246.119
R18719 a_7494_2767.n1 a_7494_2767.t5 189.588
R18720 a_7494_2767.n3 a_7494_2767.t2 89.1195
R18721 a_7494_2767.n0 a_7494_2767.t1 63.3338
R18722 a_7494_2767.t0 a_7494_2767.n3 41.0422
R18723 a_7494_2767.n0 a_7494_2767.t3 31.9797
R18724 a_9761_3311.t0 a_9761_3311.n3 370.026
R18725 a_9761_3311.n0 a_9761_3311.t2 351.356
R18726 a_9761_3311.n1 a_9761_3311.t3 334.717
R18727 a_9761_3311.n3 a_9761_3311.t1 325.971
R18728 a_9761_3311.n1 a_9761_3311.t5 309.935
R18729 a_9761_3311.n0 a_9761_3311.t4 305.683
R18730 a_9761_3311.n2 a_9761_3311.n0 16.879
R18731 a_9761_3311.n3 a_9761_3311.n2 10.8867
R18732 a_9761_3311.n2 a_9761_3311.n1 9.3005
R18733 a_10329_3553.n3 a_10329_3553.n2 647.119
R18734 a_10329_3553.n1 a_10329_3553.t4 350.253
R18735 a_10329_3553.n2 a_10329_3553.n0 260.339
R18736 a_10329_3553.n2 a_10329_3553.n1 246.119
R18737 a_10329_3553.n1 a_10329_3553.t5 189.588
R18738 a_10329_3553.n3 a_10329_3553.t3 89.1195
R18739 a_10329_3553.n0 a_10329_3553.t0 63.3338
R18740 a_10329_3553.t1 a_10329_3553.n3 41.0422
R18741 a_10329_3553.n0 a_10329_3553.t2 31.9797
R18742 a_10676_3311.n3 a_10676_3311.n2 636.953
R18743 a_10676_3311.n1 a_10676_3311.t4 366.856
R18744 a_10676_3311.n2 a_10676_3311.n0 300.2
R18745 a_10676_3311.n2 a_10676_3311.n1 225.036
R18746 a_10676_3311.n1 a_10676_3311.t5 174.056
R18747 a_10676_3311.n0 a_10676_3311.t1 70.0005
R18748 a_10676_3311.n3 a_10676_3311.t3 68.0124
R18749 a_10676_3311.t0 a_10676_3311.n3 63.3219
R18750 a_10676_3311.n0 a_10676_3311.t2 61.6672
R18751 a_8951_7663.n1 a_8951_7663.t6 530.01
R18752 a_8951_7663.t0 a_8951_7663.n5 421.021
R18753 a_8951_7663.n0 a_8951_7663.t3 337.142
R18754 a_8951_7663.n3 a_8951_7663.t1 280.223
R18755 a_8951_7663.n4 a_8951_7663.t2 263.173
R18756 a_8951_7663.n4 a_8951_7663.t4 227.826
R18757 a_8951_7663.n0 a_8951_7663.t5 199.762
R18758 a_8951_7663.n2 a_8951_7663.n1 170.81
R18759 a_8951_7663.n2 a_8951_7663.n0 167.321
R18760 a_8951_7663.n5 a_8951_7663.n4 152
R18761 a_8951_7663.n1 a_8951_7663.t7 141.923
R18762 a_8951_7663.n3 a_8951_7663.n2 10.8376
R18763 a_8951_7663.n5 a_8951_7663.n3 2.50485
R18764 a_9117_7663.t0 a_9117_7663.n3 370.026
R18765 a_9117_7663.n0 a_9117_7663.t4 351.356
R18766 a_9117_7663.n1 a_9117_7663.t3 334.717
R18767 a_9117_7663.n3 a_9117_7663.t1 325.971
R18768 a_9117_7663.n1 a_9117_7663.t5 309.935
R18769 a_9117_7663.n0 a_9117_7663.t2 305.683
R18770 a_9117_7663.n2 a_9117_7663.n0 16.879
R18771 a_9117_7663.n3 a_9117_7663.n2 10.8867
R18772 a_9117_7663.n2 a_9117_7663.n1 9.3005
R18773 a_2400_10107.t1 a_2400_10107.n3 370.026
R18774 a_2400_10107.n0 a_2400_10107.t4 351.356
R18775 a_2400_10107.n1 a_2400_10107.t5 334.717
R18776 a_2400_10107.n3 a_2400_10107.t0 325.971
R18777 a_2400_10107.n1 a_2400_10107.t2 309.935
R18778 a_2400_10107.n0 a_2400_10107.t3 305.683
R18779 a_2400_10107.n2 a_2400_10107.n0 16.879
R18780 a_2400_10107.n3 a_2400_10107.n2 10.8867
R18781 a_2400_10107.n2 a_2400_10107.n1 9.3005
R18782 a_2595_10076.n3 a_2595_10076.n2 674.338
R18783 a_2595_10076.n1 a_2595_10076.t4 332.58
R18784 a_2595_10076.n2 a_2595_10076.n0 284.012
R18785 a_2595_10076.n2 a_2595_10076.n1 253.648
R18786 a_2595_10076.n1 a_2595_10076.t5 168.701
R18787 a_2595_10076.n3 a_2595_10076.t3 96.1553
R18788 a_2595_10076.t1 a_2595_10076.n3 65.6672
R18789 a_2595_10076.n0 a_2595_10076.t0 65.0005
R18790 a_2595_10076.n0 a_2595_10076.t2 45.0005
R18791 a_3158_10205.n1 a_3158_10205.n0 926.024
R18792 a_3158_10205.n1 a_3158_10205.t3 82.0838
R18793 a_3158_10205.n0 a_3158_10205.t0 63.3338
R18794 a_3158_10205.t1 a_3158_10205.n1 63.3219
R18795 a_3158_10205.n0 a_3158_10205.t2 29.7268
R18796 a_7477_4641.n3 a_7477_4641.n2 647.119
R18797 a_7477_4641.n1 a_7477_4641.t5 350.253
R18798 a_7477_4641.n2 a_7477_4641.n0 260.339
R18799 a_7477_4641.n2 a_7477_4641.n1 246.119
R18800 a_7477_4641.n1 a_7477_4641.t4 189.588
R18801 a_7477_4641.n3 a_7477_4641.t3 89.1195
R18802 a_7477_4641.n0 a_7477_4641.t0 63.3338
R18803 a_7477_4641.t1 a_7477_4641.n3 41.0422
R18804 a_7477_4641.n0 a_7477_4641.t2 31.9797
R18805 a_7824_4399.n3 a_7824_4399.n2 636.953
R18806 a_7824_4399.n1 a_7824_4399.t5 366.856
R18807 a_7824_4399.n2 a_7824_4399.n0 300.2
R18808 a_7824_4399.n2 a_7824_4399.n1 225.036
R18809 a_7824_4399.n1 a_7824_4399.t4 174.056
R18810 a_7824_4399.n0 a_7824_4399.t0 70.0005
R18811 a_7824_4399.n3 a_7824_4399.t2 68.0124
R18812 a_7824_4399.t1 a_7824_4399.n3 63.3219
R18813 a_7824_4399.n0 a_7824_4399.t3 61.6672
R18814 a_8459_4159.n5 a_8459_4159.n4 807.871
R18815 a_8459_4159.n2 a_8459_4159.t7 389.183
R18816 a_8459_4159.n3 a_8459_4159.n2 251.167
R18817 a_8459_4159.n3 a_8459_4159.t1 223.571
R18818 a_8459_4159.n0 a_8459_4159.t8 212.081
R18819 a_8459_4159.n1 a_8459_4159.t3 212.081
R18820 a_8459_4159.n4 a_8459_4159.n1 176.576
R18821 a_8459_4159.n2 a_8459_4159.t6 174.891
R18822 a_8459_4159.n0 a_8459_4159.t4 139.78
R18823 a_8459_4159.n1 a_8459_4159.t5 139.78
R18824 a_8459_4159.n5 a_8459_4159.t2 63.3219
R18825 a_8459_4159.t0 a_8459_4159.n5 63.3219
R18826 a_8459_4159.n1 a_8459_4159.n0 61.346
R18827 a_8459_4159.n4 a_8459_4159.n3 37.7195
R18828 SWP[3].n5 SWP[3].n4 585
R18829 SWP[3].n6 SWP[3].n5 585
R18830 SWP[3].n0 SWP[3].t4 333.651
R18831 SWP[3].n0 SWP[3].t5 297.233
R18832 SWP[3].n1 SWP[3].n0 195.701
R18833 SWP[3].n3 SWP[3].n2 185
R18834 SWP[3] SWP[3].n3 57.7379
R18835 SWP[3].n8 SWP[3].n1 34.8582
R18836 SWP[3].n5 SWP[3].t0 26.5955
R18837 SWP[3].n5 SWP[3].t1 26.5955
R18838 SWP[3].n2 SWP[3].t3 24.9236
R18839 SWP[3].n2 SWP[3].t2 24.9236
R18840 SWP[3].n4 SWP[3] 10.4965
R18841 SWP[3].n6 SWP[3] 10.4965
R18842 SWP[3].n8 SWP[3].n7 9.3005
R18843 SWP[3].n4 SWP[3] 6.9125
R18844 SWP[3] SWP[3].n8 5.42117
R18845 SWP[3].n7 SWP[3] 4.3525
R18846 SWP[3].n7 SWP[3].n6 2.5605
R18847 SWP[3].n3 SWP[3] 1.7925
R18848 SWP[3].n1 SWP[3] 1.03669
R18849 a_3859_8725.n5 a_3859_8725.n4 807.871
R18850 a_3859_8725.n0 a_3859_8725.t8 389.183
R18851 a_3859_8725.n1 a_3859_8725.n0 251.167
R18852 a_3859_8725.n1 a_3859_8725.t2 223.571
R18853 a_3859_8725.n3 a_3859_8725.t7 212.081
R18854 a_3859_8725.n2 a_3859_8725.t3 212.081
R18855 a_3859_8725.n4 a_3859_8725.n3 176.576
R18856 a_3859_8725.n0 a_3859_8725.t5 174.891
R18857 a_3859_8725.n3 a_3859_8725.t4 139.78
R18858 a_3859_8725.n2 a_3859_8725.t6 139.78
R18859 a_3859_8725.t0 a_3859_8725.n5 63.3219
R18860 a_3859_8725.n5 a_3859_8725.t1 63.3219
R18861 a_3859_8725.n3 a_3859_8725.n2 61.346
R18862 a_3859_8725.n4 a_3859_8725.n1 37.5061
R18863 a_8275_6335.n5 a_8275_6335.n4 807.871
R18864 a_8275_6335.n2 a_8275_6335.t3 389.183
R18865 a_8275_6335.n3 a_8275_6335.n2 251.167
R18866 a_8275_6335.n3 a_8275_6335.t1 223.571
R18867 a_8275_6335.n0 a_8275_6335.t8 212.081
R18868 a_8275_6335.n1 a_8275_6335.t7 212.081
R18869 a_8275_6335.n4 a_8275_6335.n1 176.576
R18870 a_8275_6335.n2 a_8275_6335.t5 174.891
R18871 a_8275_6335.n0 a_8275_6335.t6 139.78
R18872 a_8275_6335.n1 a_8275_6335.t4 139.78
R18873 a_8275_6335.n5 a_8275_6335.t2 63.3219
R18874 a_8275_6335.t0 a_8275_6335.n5 63.3219
R18875 a_8275_6335.n1 a_8275_6335.n0 61.346
R18876 a_8275_6335.n4 a_8275_6335.n3 37.7195
R18877 a_10207_7637.n5 a_10207_7637.n4 807.871
R18878 a_10207_7637.n2 a_10207_7637.t5 389.183
R18879 a_10207_7637.n3 a_10207_7637.n2 251.167
R18880 a_10207_7637.n3 a_10207_7637.t1 223.571
R18881 a_10207_7637.n0 a_10207_7637.t7 212.081
R18882 a_10207_7637.n1 a_10207_7637.t6 212.081
R18883 a_10207_7637.n4 a_10207_7637.n1 176.576
R18884 a_10207_7637.n2 a_10207_7637.t8 174.891
R18885 a_10207_7637.n0 a_10207_7637.t4 139.78
R18886 a_10207_7637.n1 a_10207_7637.t3 139.78
R18887 a_10207_7637.t0 a_10207_7637.n5 63.3219
R18888 a_10207_7637.n5 a_10207_7637.t2 63.3219
R18889 a_10207_7637.n1 a_10207_7637.n0 61.346
R18890 a_10207_7637.n4 a_10207_7637.n3 37.7195
R18891 DOUT[4].n3 DOUT[4].n2 585
R18892 DOUT[4].n4 DOUT[4].n3 585
R18893 DOUT[4].n1 DOUT[4].n0 185
R18894 DOUT[4] DOUT[4].n1 49.0339
R18895 DOUT[4] DOUT[4].n4 45.4968
R18896 DOUT[4].n3 DOUT[4].t0 26.5955
R18897 DOUT[4].n3 DOUT[4].t1 26.5955
R18898 DOUT[4].n0 DOUT[4].t2 24.9236
R18899 DOUT[4].n0 DOUT[4].t3 24.9236
R18900 DOUT[4].n2 DOUT[4] 15.6165
R18901 DOUT[4].n1 DOUT[4] 10.4965
R18902 DOUT[4].n4 DOUT[4] 1.7925
R18903 DOUT[4].n2 DOUT[4] 1.7925
R18904 a_5502_3855.t0 a_5502_3855.t1 126.644
R18905 a_9687_6575.n1 a_9687_6575.t2 530.01
R18906 a_9687_6575.t0 a_9687_6575.n5 421.021
R18907 a_9687_6575.n0 a_9687_6575.t5 337.142
R18908 a_9687_6575.n3 a_9687_6575.t1 280.223
R18909 a_9687_6575.n4 a_9687_6575.t6 263.173
R18910 a_9687_6575.n4 a_9687_6575.t7 227.826
R18911 a_9687_6575.n0 a_9687_6575.t3 199.762
R18912 a_9687_6575.n2 a_9687_6575.n1 170.81
R18913 a_9687_6575.n2 a_9687_6575.n0 167.321
R18914 a_9687_6575.n5 a_9687_6575.n4 152
R18915 a_9687_6575.n1 a_9687_6575.t4 141.923
R18916 a_9687_6575.n3 a_9687_6575.n2 10.8376
R18917 a_9687_6575.n5 a_9687_6575.n3 2.50485
R18918 a_10311_6941.n0 a_10311_6941.t1 1327.82
R18919 a_10311_6941.t0 a_10311_6941.n0 194.655
R18920 a_10311_6941.n0 a_10311_6941.t2 63.3219
R18921 a_4043_7637.n5 a_4043_7637.n4 807.871
R18922 a_4043_7637.n0 a_4043_7637.t7 389.183
R18923 a_4043_7637.n1 a_4043_7637.n0 251.167
R18924 a_4043_7637.n1 a_4043_7637.t2 223.571
R18925 a_4043_7637.n3 a_4043_7637.t8 212.081
R18926 a_4043_7637.n2 a_4043_7637.t6 212.081
R18927 a_4043_7637.n4 a_4043_7637.n3 176.576
R18928 a_4043_7637.n0 a_4043_7637.t5 174.891
R18929 a_4043_7637.n3 a_4043_7637.t4 139.78
R18930 a_4043_7637.n2 a_4043_7637.t3 139.78
R18931 a_4043_7637.t0 a_4043_7637.n5 63.3219
R18932 a_4043_7637.n5 a_4043_7637.t1 63.3219
R18933 a_4043_7637.n3 a_4043_7637.n2 61.346
R18934 a_4043_7637.n4 a_4043_7637.n1 37.5061
R18935 SWN[4].n4 SWN[4].n3 585
R18936 SWN[4].n3 SWN[4].n2 585
R18937 SWN[4].n1 SWN[4].n0 185
R18938 SWN[4] SWN[4].n1 49.0339
R18939 SWN[4].n3 SWN[4].t0 26.5955
R18940 SWN[4].n3 SWN[4].t1 26.5955
R18941 SWN[4].n0 SWN[4].t2 24.9236
R18942 SWN[4].n0 SWN[4].t3 24.9236
R18943 SWN[4].n2 SWN[4] 19.7097
R18944 SWN[4].n4 SWN[4] 15.6165
R18945 SWN[4].n1 SWN[4] 10.4965
R18946 SWN[4].n2 SWN[4] 1.7925
R18947 SWN[4] SWN[4].n4 1.7925
R18948 a_9411_4949.n1 a_9411_4949.t5 530.01
R18949 a_9411_4949.t0 a_9411_4949.n5 421.021
R18950 a_9411_4949.n0 a_9411_4949.t7 337.142
R18951 a_9411_4949.n3 a_9411_4949.t1 280.223
R18952 a_9411_4949.n4 a_9411_4949.t2 263.173
R18953 a_9411_4949.n4 a_9411_4949.t3 227.826
R18954 a_9411_4949.n0 a_9411_4949.t4 199.762
R18955 a_9411_4949.n2 a_9411_4949.n1 170.81
R18956 a_9411_4949.n2 a_9411_4949.n0 167.321
R18957 a_9411_4949.n5 a_9411_4949.n4 152
R18958 a_9411_4949.n1 a_9411_4949.t6 141.923
R18959 a_9411_4949.n3 a_9411_4949.n2 10.8376
R18960 a_9411_4949.n5 a_9411_4949.n3 2.50485
R18961 a_9577_4949.t0 a_9577_4949.n3 370.026
R18962 a_9577_4949.n0 a_9577_4949.t4 351.356
R18963 a_9577_4949.n1 a_9577_4949.t2 334.717
R18964 a_9577_4949.n3 a_9577_4949.t1 325.971
R18965 a_9577_4949.n1 a_9577_4949.t3 309.935
R18966 a_9577_4949.n0 a_9577_4949.t5 305.683
R18967 a_9577_4949.n2 a_9577_4949.n0 16.879
R18968 a_9577_4949.n3 a_9577_4949.n2 10.8867
R18969 a_9577_4949.n2 a_9577_4949.n1 9.3005
R18970 CF[1].n12 CF[1].t8 333.651
R18971 CF[1].n12 CF[1].t6 297.233
R18972 CF[1].n3 CF[1].t7 294.557
R18973 CF[1].n0 CF[1].t4 294.557
R18974 CF[1].n8 CF[1].n7 289.096
R18975 CF[1].n3 CF[1].t9 211.01
R18976 CF[1].n0 CF[1].t5 211.01
R18977 CF[1] CF[1].n12 194.062
R18978 CF[1].n10 CF[1].n9 185
R18979 CF[1].n4 CF[1].n3 152
R18980 CF[1].n1 CF[1].n0 152
R18981 CF[1].n10 CF[1] 49.0339
R18982 CF[1].n7 CF[1].t1 26.5955
R18983 CF[1].n7 CF[1].t0 26.5955
R18984 CF[1].n13 CF[1] 25.857
R18985 CF[1].n9 CF[1].t2 24.9236
R18986 CF[1].n9 CF[1].t3 24.9236
R18987 CF[1].n6 CF[1].n2 23.3403
R18988 CF[1].n6 CF[1].n5 22.5189
R18989 CF[1].n13 CF[1].n11 18.7661
R18990 CF[1] CF[1].n14 17.6077
R18991 CF[1].n14 CF[1].n6 16.6667
R18992 CF[1] CF[1].n8 9.48653
R18993 CF[1].n5 CF[1] 9.32621
R18994 CF[1].n2 CF[1] 9.32621
R18995 CF[1].n8 CF[1] 7.7181
R18996 CF[1].n11 CF[1].n10 6.1445
R18997 CF[1].n14 CF[1].n13 5.18792
R18998 CF[1].n11 CF[1] 4.3525
R18999 CF[1].n4 CF[1] 2.01193
R19000 CF[1].n1 CF[1] 2.01193
R19001 CF[1].n5 CF[1].n4 1.09764
R19002 CF[1].n2 CF[1].n1 1.09764
R19003 a_6855_6717.n1 a_6855_6717.t2 530.01
R19004 a_6855_6717.t0 a_6855_6717.n5 421.021
R19005 a_6855_6717.n0 a_6855_6717.t6 337.171
R19006 a_6855_6717.n3 a_6855_6717.t1 280.223
R19007 a_6855_6717.n4 a_6855_6717.t4 263.173
R19008 a_6855_6717.n4 a_6855_6717.t5 227.826
R19009 a_6855_6717.n0 a_6855_6717.t3 199.762
R19010 a_6855_6717.n2 a_6855_6717.n1 170.81
R19011 a_6855_6717.n2 a_6855_6717.n0 167.321
R19012 a_6855_6717.n5 a_6855_6717.n4 152
R19013 a_6855_6717.n1 a_6855_6717.t7 141.923
R19014 a_6855_6717.n3 a_6855_6717.n2 10.8376
R19015 a_6855_6717.n5 a_6855_6717.n3 2.50485
R19016 a_8435_8181.n22 a_8435_8181.t4 286.348
R19017 a_8435_8181.n24 a_8435_8181.t1 271.051
R19018 a_8435_8181.n1 a_8435_8181.t13 221.72
R19019 a_8435_8181.n18 a_8435_8181.t15 221.72
R19020 a_8435_8181.n2 a_8435_8181.t9 221.72
R19021 a_8435_8181.n12 a_8435_8181.t20 221.72
R19022 a_8435_8181.n10 a_8435_8181.t10 221.72
R19023 a_8435_8181.n4 a_8435_8181.t16 221.72
R19024 a_8435_8181.n6 a_8435_8181.t7 221.72
R19025 a_8435_8181.n5 a_8435_8181.t18 221.72
R19026 a_8435_8181.n25 a_8435_8181.n24 206.055
R19027 a_8435_8181.n22 a_8435_8181.n21 198.177
R19028 a_8435_8181.n8 a_8435_8181.n7 177.601
R19029 a_8435_8181.n9 a_8435_8181.n8 152
R19030 a_8435_8181.n11 a_8435_8181.n3 152
R19031 a_8435_8181.n14 a_8435_8181.n13 152
R19032 a_8435_8181.n16 a_8435_8181.n15 152
R19033 a_8435_8181.n17 a_8435_8181.n0 152
R19034 a_8435_8181.n20 a_8435_8181.n19 152
R19035 a_8435_8181.n1 a_8435_8181.t6 149.421
R19036 a_8435_8181.n18 a_8435_8181.t8 149.421
R19037 a_8435_8181.n2 a_8435_8181.t19 149.421
R19038 a_8435_8181.n12 a_8435_8181.t14 149.421
R19039 a_8435_8181.n10 a_8435_8181.t21 149.421
R19040 a_8435_8181.n4 a_8435_8181.t11 149.421
R19041 a_8435_8181.n6 a_8435_8181.t17 149.421
R19042 a_8435_8181.n5 a_8435_8181.t12 149.421
R19043 a_8435_8181.n6 a_8435_8181.n5 74.9783
R19044 a_8435_8181.n7 a_8435_8181.n6 66.0523
R19045 a_8435_8181.n17 a_8435_8181.n16 60.6968
R19046 a_8435_8181.n19 a_8435_8181.n18 55.3412
R19047 a_8435_8181.n13 a_8435_8181.n2 51.7709
R19048 a_8435_8181.n9 a_8435_8181.n4 51.7709
R19049 a_8435_8181.n23 a_8435_8181.n22 48.9632
R19050 a_8435_8181.n24 a_8435_8181.n23 38.7339
R19051 a_8435_8181.n12 a_8435_8181.n11 37.4894
R19052 a_8435_8181.n11 a_8435_8181.n10 37.4894
R19053 a_8435_8181.n25 a_8435_8181.t5 26.5955
R19054 a_8435_8181.t0 a_8435_8181.n25 26.5955
R19055 a_8435_8181.n20 a_8435_8181.n0 25.6005
R19056 a_8435_8181.n15 a_8435_8181.n0 25.6005
R19057 a_8435_8181.n15 a_8435_8181.n14 25.6005
R19058 a_8435_8181.n14 a_8435_8181.n3 25.6005
R19059 a_8435_8181.n8 a_8435_8181.n3 25.6005
R19060 a_8435_8181.n21 a_8435_8181.t2 24.9236
R19061 a_8435_8181.n21 a_8435_8181.t3 24.9236
R19062 a_8435_8181.n13 a_8435_8181.n12 23.2079
R19063 a_8435_8181.n10 a_8435_8181.n9 23.2079
R19064 a_8435_8181.n19 a_8435_8181.n1 19.6375
R19065 a_8435_8181.n23 a_8435_8181.n20 18.4476
R19066 a_8435_8181.n16 a_8435_8181.n2 8.92643
R19067 a_8435_8181.n7 a_8435_8181.n4 8.92643
R19068 a_8435_8181.n18 a_8435_8181.n17 5.35606
R19069 x3/COMP_BUF_P.n3 x3/COMP_BUF_P.n2 374.966
R19070 x3/COMP_BUF_P.n31 x3/COMP_BUF_P.t34 333.651
R19071 x3/COMP_BUF_P.n28 x3/COMP_BUF_P.t17 333.651
R19072 x3/COMP_BUF_P.n24 x3/COMP_BUF_P.t31 333.651
R19073 x3/COMP_BUF_P.n18 x3/COMP_BUF_P.t35 333.651
R19074 x3/COMP_BUF_P.n12 x3/COMP_BUF_P.t30 333.651
R19075 x3/COMP_BUF_P.n29 x3/COMP_BUF_P.t23 332.312
R19076 x3/COMP_BUF_P.n22 x3/COMP_BUF_P.t26 332.312
R19077 x3/COMP_BUF_P.n17 x3/COMP_BUF_P.t25 332.312
R19078 x3/COMP_BUF_P.n15 x3/COMP_BUF_P.t21 332.312
R19079 x3/COMP_BUF_P.n14 x3/COMP_BUF_P.t32 332.312
R19080 x3/COMP_BUF_P.n4 x3/COMP_BUF_P.n0 311.719
R19081 x3/COMP_BUF_P.n3 x3/COMP_BUF_P.n1 311.719
R19082 x3/COMP_BUF_P x3/COMP_BUF_P.n34 311.719
R19083 x3/COMP_BUF_P.n31 x3/COMP_BUF_P.t29 297.233
R19084 x3/COMP_BUF_P.n28 x3/COMP_BUF_P.t33 297.233
R19085 x3/COMP_BUF_P.n24 x3/COMP_BUF_P.t18 297.233
R19086 x3/COMP_BUF_P.n18 x3/COMP_BUF_P.t28 297.233
R19087 x3/COMP_BUF_P.n12 x3/COMP_BUF_P.t19 297.233
R19088 x3/COMP_BUF_P.n29 x3/COMP_BUF_P.t24 295.627
R19089 x3/COMP_BUF_P.n22 x3/COMP_BUF_P.t27 295.627
R19090 x3/COMP_BUF_P.n17 x3/COMP_BUF_P.t16 295.627
R19091 x3/COMP_BUF_P.n15 x3/COMP_BUF_P.t22 295.627
R19092 x3/COMP_BUF_P.n14 x3/COMP_BUF_P.t20 295.627
R19093 x3/COMP_BUF_P.n8 x3/COMP_BUF_P.n7 261.425
R19094 x3/COMP_BUF_P.n11 x3/COMP_BUF_P.n10 202.444
R19095 x3/COMP_BUF_P.n8 x3/COMP_BUF_P.n6 198.177
R19096 x3/COMP_BUF_P.n9 x3/COMP_BUF_P.n5 198.177
R19097 x3/COMP_BUF_P.n25 x3/COMP_BUF_P.n24 196.493
R19098 x3/COMP_BUF_P x3/COMP_BUF_P.n22 196.004
R19099 x3/COMP_BUF_P x3/COMP_BUF_P.n17 196.004
R19100 x3/COMP_BUF_P x3/COMP_BUF_P.n15 196.004
R19101 x3/COMP_BUF_P x3/COMP_BUF_P.n14 196.004
R19102 x3/COMP_BUF_P x3/COMP_BUF_P.n29 195.401
R19103 x3/COMP_BUF_P x3/COMP_BUF_P.n28 194.062
R19104 x3/COMP_BUF_P.n32 x3/COMP_BUF_P.n31 193.506
R19105 x3/COMP_BUF_P.n19 x3/COMP_BUF_P.n18 193.506
R19106 x3/COMP_BUF_P.n13 x3/COMP_BUF_P.n12 193.506
R19107 x3/COMP_BUF_P.n4 x3/COMP_BUF_P.n3 63.2476
R19108 x3/COMP_BUF_P.n9 x3/COMP_BUF_P.n8 63.2476
R19109 x3/COMP_BUF_P.n33 x3/COMP_BUF_P.n4 50.4476
R19110 x3/COMP_BUF_P.n11 x3/COMP_BUF_P.n9 50.4476
R19111 x3/COMP_BUF_P.n27 x3/COMP_BUF_P.n13 33.5138
R19112 x3/COMP_BUF_P.n23 x3/COMP_BUF_P 32.5327
R19113 x3/COMP_BUF_P.n33 x3/COMP_BUF_P 32.2272
R19114 x3/COMP_BUF_P.n20 x3/COMP_BUF_P.n19 31.2077
R19115 x3/COMP_BUF_P.n26 x3/COMP_BUF_P.n25 30.7651
R19116 x3/COMP_BUF_P.n30 x3/COMP_BUF_P 29.8476
R19117 x3/COMP_BUF_P.n0 x3/COMP_BUF_P.t5 26.5955
R19118 x3/COMP_BUF_P.n0 x3/COMP_BUF_P.t2 26.5955
R19119 x3/COMP_BUF_P.n1 x3/COMP_BUF_P.t6 26.5955
R19120 x3/COMP_BUF_P.n1 x3/COMP_BUF_P.t0 26.5955
R19121 x3/COMP_BUF_P.n2 x3/COMP_BUF_P.t4 26.5955
R19122 x3/COMP_BUF_P.n2 x3/COMP_BUF_P.t3 26.5955
R19123 x3/COMP_BUF_P.n34 x3/COMP_BUF_P.t7 26.5955
R19124 x3/COMP_BUF_P.n34 x3/COMP_BUF_P.t1 26.5955
R19125 x3/COMP_BUF_P x3/COMP_BUF_P.n32 26.4135
R19126 x3/COMP_BUF_P.n30 x3/COMP_BUF_P 25.857
R19127 x3/COMP_BUF_P.n20 x3/COMP_BUF_P 25.8025
R19128 x3/COMP_BUF_P.n7 x3/COMP_BUF_P.t15 24.9236
R19129 x3/COMP_BUF_P.n7 x3/COMP_BUF_P.t14 24.9236
R19130 x3/COMP_BUF_P.n6 x3/COMP_BUF_P.t9 24.9236
R19131 x3/COMP_BUF_P.n6 x3/COMP_BUF_P.t11 24.9236
R19132 x3/COMP_BUF_P.n5 x3/COMP_BUF_P.t8 24.9236
R19133 x3/COMP_BUF_P.n5 x3/COMP_BUF_P.t13 24.9236
R19134 x3/COMP_BUF_P.n10 x3/COMP_BUF_P.t10 24.9236
R19135 x3/COMP_BUF_P.n10 x3/COMP_BUF_P.t12 24.9236
R19136 x3/COMP_BUF_P.n16 x3/COMP_BUF_P 22.4782
R19137 x3/COMP_BUF_P.n33 x3/COMP_BUF_P 12.8005
R19138 x3/COMP_BUF_P x3/COMP_BUF_P.n30 12.6567
R19139 x3/COMP_BUF_P.n16 x3/COMP_BUF_P 11.286
R19140 x3/COMP_BUF_P.n30 x3/COMP_BUF_P.n27 9.11176
R19141 x3/COMP_BUF_P.n26 x3/COMP_BUF_P.n23 7.15364
R19142 x3/COMP_BUF_P.n21 x3/COMP_BUF_P.n20 7.10077
R19143 x3/COMP_BUF_P.n27 x3/COMP_BUF_P.n26 6.49551
R19144 x3/COMP_BUF_P x3/COMP_BUF_P.n11 5.77305
R19145 x3/COMP_BUF_P.n21 x3/COMP_BUF_P.n16 5.04171
R19146 x3/COMP_BUF_P x3/COMP_BUF_P.n33 4.26717
R19147 x3/COMP_BUF_P.n32 x3/COMP_BUF_P 4.17441
R19148 x3/COMP_BUF_P.n19 x3/COMP_BUF_P 4.17441
R19149 x3/COMP_BUF_P.n13 x3/COMP_BUF_P 4.17441
R19150 x3/COMP_BUF_P.n23 x3/COMP_BUF_P.n21 3.24998
R19151 x3/COMP_BUF_P.n25 x3/COMP_BUF_P 0.24431
R19152 a_7563_2741.n3 a_7563_2741.n2 674.338
R19153 a_7563_2741.n1 a_7563_2741.t4 332.58
R19154 a_7563_2741.n2 a_7563_2741.n0 284.012
R19155 a_7563_2741.n2 a_7563_2741.n1 253.648
R19156 a_7563_2741.n1 a_7563_2741.t5 168.701
R19157 a_7563_2741.n3 a_7563_2741.t3 96.1553
R19158 a_7563_2741.t0 a_7563_2741.n3 65.6672
R19159 a_7563_2741.n0 a_7563_2741.t2 65.0005
R19160 a_7563_2741.n0 a_7563_2741.t1 45.0005
R19161 a_10032_7663.n3 a_10032_7663.n2 636.953
R19162 a_10032_7663.n1 a_10032_7663.t5 366.856
R19163 a_10032_7663.n2 a_10032_7663.n0 300.2
R19164 a_10032_7663.n2 a_10032_7663.n1 225.036
R19165 a_10032_7663.n1 a_10032_7663.t4 174.056
R19166 a_10032_7663.n0 a_10032_7663.t0 70.0005
R19167 a_10032_7663.n3 a_10032_7663.t2 68.0124
R19168 a_10032_7663.t1 a_10032_7663.n3 63.3219
R19169 a_10032_7663.n0 a_10032_7663.t3 61.6672
R19170 a_2032_8323.t1 a_2032_8323.n3 370.026
R19171 a_2032_8323.n0 a_2032_8323.t2 351.356
R19172 a_2032_8323.n1 a_2032_8323.t3 334.717
R19173 a_2032_8323.n3 a_2032_8323.t0 325.971
R19174 a_2032_8323.n1 a_2032_8323.t5 309.935
R19175 a_2032_8323.n0 a_2032_8323.t4 305.683
R19176 a_2032_8323.n2 a_2032_8323.n0 16.879
R19177 a_2032_8323.n3 a_2032_8323.n2 10.8867
R19178 a_2032_8323.n2 a_2032_8323.n1 9.3005
R19179 a_1754_8339.n3 a_1754_8339.n2 636.953
R19180 a_1754_8339.n1 a_1754_8339.t5 366.856
R19181 a_1754_8339.n2 a_1754_8339.n0 300.2
R19182 a_1754_8339.n2 a_1754_8339.n1 225.036
R19183 a_1754_8339.n1 a_1754_8339.t4 174.056
R19184 a_1754_8339.n0 a_1754_8339.t2 70.0005
R19185 a_1754_8339.t0 a_1754_8339.n3 68.0124
R19186 a_1754_8339.n3 a_1754_8339.t1 63.3219
R19187 a_1754_8339.n0 a_1754_8339.t3 61.6672
R19188 a_2158_8207.n3 a_2158_8207.n2 647.119
R19189 a_2158_8207.n1 a_2158_8207.t4 350.253
R19190 a_2158_8207.n2 a_2158_8207.n0 260.339
R19191 a_2158_8207.n2 a_2158_8207.n1 246.119
R19192 a_2158_8207.n1 a_2158_8207.t5 189.588
R19193 a_2158_8207.n3 a_2158_8207.t0 89.1195
R19194 a_2158_8207.n0 a_2158_8207.t1 63.3338
R19195 a_2158_8207.t2 a_2158_8207.n3 41.0422
R19196 a_2158_8207.n0 a_2158_8207.t3 31.9797
R19197 a_7654_4943.n52 a_7654_4943.n51 330.308
R19198 a_7654_4943.n50 a_7654_4943.n2 327.253
R19199 a_7654_4943.n50 a_7654_4943.n1 217.256
R19200 a_7654_4943.n51 a_7654_4943.n0 217.256
R19201 a_7654_4943.n12 a_7654_4943.t22 212.081
R19202 a_7654_4943.n13 a_7654_4943.t25 212.081
R19203 a_7654_4943.n14 a_7654_4943.t23 212.081
R19204 a_7654_4943.n16 a_7654_4943.t12 212.081
R19205 a_7654_4943.n18 a_7654_4943.t8 212.081
R19206 a_7654_4943.n10 a_7654_4943.t36 212.081
R19207 a_7654_4943.n24 a_7654_4943.t14 212.081
R19208 a_7654_4943.n8 a_7654_4943.t10 212.081
R19209 a_7654_4943.n29 a_7654_4943.t38 212.081
R19210 a_7654_4943.n6 a_7654_4943.t35 212.081
R19211 a_7654_4943.n35 a_7654_4943.t31 212.081
R19212 a_7654_4943.n37 a_7654_4943.t29 212.081
R19213 a_7654_4943.n38 a_7654_4943.t27 212.081
R19214 a_7654_4943.n44 a_7654_4943.t33 212.081
R19215 a_7654_4943.n46 a_7654_4943.t30 212.081
R19216 a_7654_4943.n47 a_7654_4943.t20 212.081
R19217 a_7654_4943.n15 a_7654_4943.n11 169.409
R19218 a_7654_4943.n12 a_7654_4943.t26 162.274
R19219 a_7654_4943.n13 a_7654_4943.t32 162.274
R19220 a_7654_4943.n14 a_7654_4943.t28 162.274
R19221 a_7654_4943.n16 a_7654_4943.t19 162.274
R19222 a_7654_4943.n18 a_7654_4943.t17 162.274
R19223 a_7654_4943.n10 a_7654_4943.t15 162.274
R19224 a_7654_4943.n24 a_7654_4943.t21 162.274
R19225 a_7654_4943.n8 a_7654_4943.t18 162.274
R19226 a_7654_4943.n29 a_7654_4943.t16 162.274
R19227 a_7654_4943.n6 a_7654_4943.t13 162.274
R19228 a_7654_4943.n35 a_7654_4943.t9 162.274
R19229 a_7654_4943.n37 a_7654_4943.t37 162.274
R19230 a_7654_4943.n38 a_7654_4943.t34 162.274
R19231 a_7654_4943.n44 a_7654_4943.t11 162.274
R19232 a_7654_4943.n46 a_7654_4943.t39 162.274
R19233 a_7654_4943.n47 a_7654_4943.t24 162.274
R19234 a_7654_4943.n49 a_7654_4943.n48 152
R19235 a_7654_4943.n45 a_7654_4943.n3 152
R19236 a_7654_4943.n43 a_7654_4943.n42 152
R19237 a_7654_4943.n41 a_7654_4943.n4 152
R19238 a_7654_4943.n40 a_7654_4943.n39 152
R19239 a_7654_4943.n36 a_7654_4943.n5 152
R19240 a_7654_4943.n34 a_7654_4943.n33 152
R19241 a_7654_4943.n32 a_7654_4943.n31 152
R19242 a_7654_4943.n30 a_7654_4943.n7 152
R19243 a_7654_4943.n28 a_7654_4943.n27 152
R19244 a_7654_4943.n26 a_7654_4943.n25 152
R19245 a_7654_4943.n23 a_7654_4943.n9 152
R19246 a_7654_4943.n22 a_7654_4943.n21 152
R19247 a_7654_4943.n20 a_7654_4943.n19 152
R19248 a_7654_4943.n17 a_7654_4943.n11 152
R19249 a_7654_4943.n13 a_7654_4943.n12 55.2698
R19250 a_7654_4943.n14 a_7654_4943.n13 55.2698
R19251 a_7654_4943.n51 a_7654_4943.n50 44.0325
R19252 a_7654_4943.n23 a_7654_4943.n22 43.7018
R19253 a_7654_4943.n31 a_7654_4943.n30 43.7018
R19254 a_7654_4943.n43 a_7654_4943.n4 43.7018
R19255 a_7654_4943.n50 a_7654_4943.n49 43.5205
R19256 a_7654_4943.n19 a_7654_4943.n10 43.0592
R19257 a_7654_4943.n34 a_7654_4943.n6 42.4165
R19258 a_7654_4943.n1 a_7654_4943.t4 40.0005
R19259 a_7654_4943.n1 a_7654_4943.t5 40.0005
R19260 a_7654_4943.n0 a_7654_4943.t6 40.0005
R19261 a_7654_4943.n0 a_7654_4943.t7 40.0005
R19262 a_7654_4943.n45 a_7654_4943.n44 39.8458
R19263 a_7654_4943.n39 a_7654_4943.n38 35.9898
R19264 a_7654_4943.n15 a_7654_4943.n14 35.3472
R19265 a_7654_4943.n29 a_7654_4943.n28 33.4192
R19266 a_7654_4943.n25 a_7654_4943.n24 32.7765
R19267 a_7654_4943.n18 a_7654_4943.n17 31.4912
R19268 a_7654_4943.n36 a_7654_4943.n35 30.8485
R19269 a_7654_4943.n48 a_7654_4943.n46 28.2778
R19270 a_7654_4943.n2 a_7654_4943.t0 27.5805
R19271 a_7654_4943.n2 a_7654_4943.t1 27.5805
R19272 a_7654_4943.n52 a_7654_4943.t2 27.5805
R19273 a_7654_4943.t3 a_7654_4943.n52 27.5805
R19274 a_7654_4943.n48 a_7654_4943.n47 26.9925
R19275 a_7654_4943.n37 a_7654_4943.n36 24.4218
R19276 a_7654_4943.n17 a_7654_4943.n16 23.7792
R19277 a_7654_4943.n25 a_7654_4943.n8 22.4938
R19278 a_7654_4943.n28 a_7654_4943.n8 21.2085
R19279 a_7654_4943.n16 a_7654_4943.n15 19.9232
R19280 a_7654_4943.n39 a_7654_4943.n37 19.2805
R19281 a_7654_4943.n20 a_7654_4943.n11 17.4085
R19282 a_7654_4943.n21 a_7654_4943.n20 17.4085
R19283 a_7654_4943.n21 a_7654_4943.n9 17.4085
R19284 a_7654_4943.n26 a_7654_4943.n9 17.4085
R19285 a_7654_4943.n27 a_7654_4943.n26 17.4085
R19286 a_7654_4943.n27 a_7654_4943.n7 17.4085
R19287 a_7654_4943.n32 a_7654_4943.n7 17.4085
R19288 a_7654_4943.n33 a_7654_4943.n32 17.4085
R19289 a_7654_4943.n33 a_7654_4943.n5 17.4085
R19290 a_7654_4943.n40 a_7654_4943.n5 17.4085
R19291 a_7654_4943.n41 a_7654_4943.n40 17.4085
R19292 a_7654_4943.n42 a_7654_4943.n41 17.4085
R19293 a_7654_4943.n42 a_7654_4943.n3 17.4085
R19294 a_7654_4943.n49 a_7654_4943.n3 17.4085
R19295 a_7654_4943.n46 a_7654_4943.n45 15.4245
R19296 a_7654_4943.n35 a_7654_4943.n34 12.8538
R19297 a_7654_4943.n19 a_7654_4943.n18 12.2112
R19298 a_7654_4943.n24 a_7654_4943.n23 10.9258
R19299 a_7654_4943.n30 a_7654_4943.n29 10.2832
R19300 a_7654_4943.n38 a_7654_4943.n4 7.7125
R19301 a_7654_4943.n44 a_7654_4943.n43 3.8565
R19302 a_7654_4943.n31 a_7654_4943.n6 1.28583
R19303 a_7654_4943.n22 a_7654_4943.n10 0.643167
R19304 a_3859_6549.n5 a_3859_6549.n4 807.871
R19305 a_3859_6549.n0 a_3859_6549.t8 389.183
R19306 a_3859_6549.n1 a_3859_6549.n0 251.167
R19307 a_3859_6549.n1 a_3859_6549.t1 223.571
R19308 a_3859_6549.n3 a_3859_6549.t5 212.081
R19309 a_3859_6549.n2 a_3859_6549.t6 212.081
R19310 a_3859_6549.n4 a_3859_6549.n3 176.576
R19311 a_3859_6549.n0 a_3859_6549.t3 174.891
R19312 a_3859_6549.n3 a_3859_6549.t7 139.78
R19313 a_3859_6549.n2 a_3859_6549.t4 139.78
R19314 a_3859_6549.t0 a_3859_6549.n5 63.3219
R19315 a_3859_6549.n5 a_3859_6549.t2 63.3219
R19316 a_3859_6549.n3 a_3859_6549.n2 61.346
R19317 a_3859_6549.n4 a_3859_6549.n1 37.5061
R19318 a_4421_6575.n0 a_4421_6575.t1 68.3338
R19319 a_4421_6575.n0 a_4421_6575.t0 26.3935
R19320 a_4421_6575.n1 a_4421_6575.n0 14.4005
R19321 a_6796_8573.n1 a_6796_8573.n0 926.024
R19322 a_6796_8573.t1 a_6796_8573.n1 82.0838
R19323 a_6796_8573.n0 a_6796_8573.t0 63.3338
R19324 a_6796_8573.n1 a_6796_8573.t2 63.3219
R19325 a_6796_8573.n0 a_6796_8573.t3 29.7268
R19326 a_6891_8585.n3 a_6891_8585.n2 674.338
R19327 a_6891_8585.n1 a_6891_8585.t5 332.58
R19328 a_6891_8585.n2 a_6891_8585.n0 284.012
R19329 a_6891_8585.n2 a_6891_8585.n1 253.648
R19330 a_6891_8585.n1 a_6891_8585.t4 168.701
R19331 a_6891_8585.t1 a_6891_8585.n3 96.1553
R19332 a_6891_8585.n3 a_6891_8585.t2 65.6672
R19333 a_6891_8585.n0 a_6891_8585.t0 65.0005
R19334 a_6891_8585.n0 a_6891_8585.t3 45.0005
R19335 a_7090_9003.n3 a_7090_9003.n2 636.953
R19336 a_7090_9003.n1 a_7090_9003.t4 366.856
R19337 a_7090_9003.n2 a_7090_9003.n0 300.2
R19338 a_7090_9003.n2 a_7090_9003.n1 225.036
R19339 a_7090_9003.n1 a_7090_9003.t5 174.056
R19340 a_7090_9003.n0 a_7090_9003.t2 70.0005
R19341 a_7090_9003.t0 a_7090_9003.n3 68.0124
R19342 a_7090_9003.n3 a_7090_9003.t1 63.3219
R19343 a_7090_9003.n0 a_7090_9003.t3 61.6672
R19344 a_6803_8725.n3 a_6803_8725.n0 807.871
R19345 a_6803_8725.n4 a_6803_8725.t6 389.183
R19346 a_6803_8725.n5 a_6803_8725.n4 251.167
R19347 a_6803_8725.t0 a_6803_8725.n5 223.571
R19348 a_6803_8725.n2 a_6803_8725.t5 212.081
R19349 a_6803_8725.n1 a_6803_8725.t7 212.081
R19350 a_6803_8725.n3 a_6803_8725.n2 176.576
R19351 a_6803_8725.n4 a_6803_8725.t3 174.891
R19352 a_6803_8725.n2 a_6803_8725.t8 139.78
R19353 a_6803_8725.n1 a_6803_8725.t4 139.78
R19354 a_6803_8725.n0 a_6803_8725.t2 63.3219
R19355 a_6803_8725.n0 a_6803_8725.t1 63.3219
R19356 a_6803_8725.n2 a_6803_8725.n1 61.346
R19357 a_6803_8725.n5 a_6803_8725.n3 37.5061
R19358 a_7125_8751.t0 a_7125_8751.t1 87.1434
R19359 a_2143_10389.n1 a_2143_10389.t3 530.01
R19360 a_2143_10389.t0 a_2143_10389.n5 421.021
R19361 a_2143_10389.n0 a_2143_10389.t6 337.142
R19362 a_2143_10389.n3 a_2143_10389.t1 280.223
R19363 a_2143_10389.n4 a_2143_10389.t2 263.173
R19364 a_2143_10389.n4 a_2143_10389.t4 227.826
R19365 a_2143_10389.n0 a_2143_10389.t5 199.762
R19366 a_2143_10389.n2 a_2143_10389.n1 170.81
R19367 a_2143_10389.n2 a_2143_10389.n0 167.321
R19368 a_2143_10389.n5 a_2143_10389.n4 152
R19369 a_2143_10389.n1 a_2143_10389.t7 141.923
R19370 a_2143_10389.n3 a_2143_10389.n2 10.8376
R19371 a_2143_10389.n5 a_2143_10389.n3 2.50485
R19372 a_2309_10389.t0 a_2309_10389.n3 370.026
R19373 a_2309_10389.n0 a_2309_10389.t5 351.356
R19374 a_2309_10389.n1 a_2309_10389.t3 334.717
R19375 a_2309_10389.n3 a_2309_10389.t1 325.971
R19376 a_2309_10389.n1 a_2309_10389.t4 309.935
R19377 a_2309_10389.n0 a_2309_10389.t2 305.683
R19378 a_2309_10389.n2 a_2309_10389.n0 16.879
R19379 a_2309_10389.n3 a_2309_10389.n2 10.8867
R19380 a_2309_10389.n2 a_2309_10389.n1 9.3005
R19381 CF[3].n11 CF[3].n10 585
R19382 CF[3].n10 CF[3].n9 585
R19383 CF[3].n6 CF[3].t9 332.312
R19384 CF[3].n6 CF[3].t4 295.627
R19385 CF[3].n3 CF[3].t5 294.557
R19386 CF[3].n0 CF[3].t6 294.557
R19387 CF[3].n3 CF[3].t7 211.01
R19388 CF[3].n0 CF[3].t8 211.01
R19389 CF[3].n7 CF[3].n6 194.845
R19390 CF[3].n13 CF[3].n12 185
R19391 CF[3] CF[3].n3 156.207
R19392 CF[3].n1 CF[3].n0 152
R19393 CF[3].n13 CF[3] 57.7379
R19394 CF[3].n5 CF[3].n2 36.8378
R19395 CF[3].n8 CF[3].n7 28.3505
R19396 CF[3].n10 CF[3].t1 26.5955
R19397 CF[3].n10 CF[3].t2 26.5955
R19398 CF[3].n12 CF[3].t3 24.9236
R19399 CF[3].n12 CF[3].t0 24.9236
R19400 CF[3].n5 CF[3].n4 21.2082
R19401 CF[3].n14 CF[3] 13.6525
R19402 CF[3] CF[3].n14 13.4644
R19403 CF[3].n14 CF[3].n8 11.1641
R19404 CF[3] CF[3].n11 10.4965
R19405 CF[3].n9 CF[3] 10.4965
R19406 CF[3].n4 CF[3] 9.32621
R19407 CF[3].n2 CF[3] 9.32621
R19408 CF[3].n8 CF[3].n5 8.01149
R19409 CF[3].n11 CF[3] 6.9125
R19410 CF[3].n9 CF[3] 6.9125
R19411 CF[3].n7 CF[3] 4.17441
R19412 CF[3].n4 CF[3] 3.10907
R19413 CF[3].n1 CF[3] 2.01193
R19414 CF[3] CF[3].n13 1.7925
R19415 CF[3].n2 CF[3].n1 1.09764
R19416 a_8126_2767.n1 a_8126_2767.n0 926.024
R19417 a_8126_2767.n1 a_8126_2767.t2 82.0838
R19418 a_8126_2767.n0 a_8126_2767.t3 63.3338
R19419 a_8126_2767.t0 a_8126_2767.n1 63.3219
R19420 a_8126_2767.n0 a_8126_2767.t1 29.7268
R19421 x2/net3.n3 x2/net3.n2 585
R19422 x2/net3.n4 x2/net3.n3 585
R19423 x2/net3.n5 x2/net3.t4 333.651
R19424 x2/net3.n5 x2/net3.t5 297.233
R19425 x2/net3 x2/net3.n5 194.062
R19426 x2/net3.n1 x2/net3.n0 185
R19427 x2/net3 x2/net3.n1 57.7379
R19428 x2/net3.n3 x2/net3.t0 26.5955
R19429 x2/net3.n3 x2/net3.t1 26.5955
R19430 x2/net3.n0 x2/net3.t3 24.9236
R19431 x2/net3.n0 x2/net3.t2 24.9236
R19432 x2/net3.n6 x2/net3 19.1983
R19433 x2/net3.n2 x2/net3 10.4965
R19434 x2/net3.n4 x2/net3 10.4965
R19435 x2/net3.n2 x2/net3 6.9125
R19436 x2/net3 x2/net3.n6 4.3525
R19437 x2/net3.n6 x2/net3.n4 2.5605
R19438 x2/net3.n1 x2/net3 1.7925
R19439 a_7348_10927.n1 a_7348_10927.n0 926.024
R19440 a_7348_10927.n1 a_7348_10927.t2 82.0838
R19441 a_7348_10927.n0 a_7348_10927.t3 63.3338
R19442 a_7348_10927.t0 a_7348_10927.n1 63.3219
R19443 a_7348_10927.n0 a_7348_10927.t1 29.7268
R19444 x2/net9.n5 x2/net9.n4 585
R19445 x2/net9.n6 x2/net9.n5 585
R19446 x2/net9.n2 x2/net9.t5 333.651
R19447 x2/net9.n2 x2/net9.t4 297.233
R19448 x2/net9.n3 x2/net9.n2 195.701
R19449 x2/net9.n1 x2/net9.n0 185
R19450 x2/net9 x2/net9.n1 49.0339
R19451 x2/net9.n5 x2/net9.t0 26.5955
R19452 x2/net9.n5 x2/net9.t1 26.5955
R19453 x2/net9.n0 x2/net9.t3 24.9236
R19454 x2/net9.n0 x2/net9.t2 24.9236
R19455 x2/net9.n4 x2/net9 20.6333
R19456 x2/net9.n6 x2/net9 15.6165
R19457 x2/net9 x2/net9.n3 14.4935
R19458 x2/net9.n1 x2/net9 10.4965
R19459 x2/net9.n4 x2/net9 1.7925
R19460 x2/net9 x2/net9.n6 1.7925
R19461 x2/net9.n3 x2/net9 1.03669
R19462 a_4411_6005.n5 a_4411_6005.n4 807.871
R19463 a_4411_6005.n0 a_4411_6005.t6 389.183
R19464 a_4411_6005.n1 a_4411_6005.n0 251.167
R19465 a_4411_6005.n1 a_4411_6005.t1 223.571
R19466 a_4411_6005.n3 a_4411_6005.t3 212.081
R19467 a_4411_6005.n2 a_4411_6005.t7 212.081
R19468 a_4411_6005.n4 a_4411_6005.n3 176.576
R19469 a_4411_6005.n0 a_4411_6005.t5 174.891
R19470 a_4411_6005.n3 a_4411_6005.t8 139.78
R19471 a_4411_6005.n2 a_4411_6005.t4 139.78
R19472 a_4411_6005.t0 a_4411_6005.n5 63.3219
R19473 a_4411_6005.n5 a_4411_6005.t2 63.3219
R19474 a_4411_6005.n3 a_4411_6005.n2 61.346
R19475 a_4411_6005.n4 a_4411_6005.n1 37.5061
R19476 SWN[2].n2 SWN[2].n1 585
R19477 SWN[2].n1 SWN[2].n0 585
R19478 SWN[2].n4 SWN[2].n3 185
R19479 SWN[2].n4 SWN[2] 57.7379
R19480 SWN[2].n1 SWN[2].t1 26.5955
R19481 SWN[2].n1 SWN[2].t0 26.5955
R19482 SWN[2].n3 SWN[2].t2 24.9236
R19483 SWN[2].n3 SWN[2].t3 24.9236
R19484 SWN[2] SWN[2].n2 10.4965
R19485 SWN[2].n0 SWN[2] 10.4965
R19486 SWN[2].n2 SWN[2] 6.9125
R19487 SWN[2].n0 SWN[2] 6.9125
R19488 SWN[2] SWN[2].n4 1.7925
R19489 a_1775_10927.n1 a_1775_10927.t3 530.01
R19490 a_1775_10927.t0 a_1775_10927.n5 421.021
R19491 a_1775_10927.n0 a_1775_10927.t4 337.142
R19492 a_1775_10927.n3 a_1775_10927.t1 280.223
R19493 a_1775_10927.n4 a_1775_10927.t7 263.173
R19494 a_1775_10927.n4 a_1775_10927.t6 227.826
R19495 a_1775_10927.n0 a_1775_10927.t2 199.762
R19496 a_1775_10927.n2 a_1775_10927.n1 170.81
R19497 a_1775_10927.n2 a_1775_10927.n0 167.321
R19498 a_1775_10927.n5 a_1775_10927.n4 152
R19499 a_1775_10927.n1 a_1775_10927.t5 141.923
R19500 a_1775_10927.n3 a_1775_10927.n2 10.8376
R19501 a_1775_10927.n5 a_1775_10927.n3 2.50485
R19502 a_2856_10927.n3 a_2856_10927.n2 636.953
R19503 a_2856_10927.n1 a_2856_10927.t5 366.856
R19504 a_2856_10927.n2 a_2856_10927.n0 300.2
R19505 a_2856_10927.n2 a_2856_10927.n1 225.036
R19506 a_2856_10927.n1 a_2856_10927.t4 174.056
R19507 a_2856_10927.n0 a_2856_10927.t0 70.0005
R19508 a_2856_10927.n3 a_2856_10927.t2 68.0124
R19509 a_2856_10927.t1 a_2856_10927.n3 63.3219
R19510 a_2856_10927.n0 a_2856_10927.t3 61.6672
R19511 a_2840_11837.n1 a_2840_11837.n0 926.024
R19512 a_2840_11837.t0 a_2840_11837.n1 82.0838
R19513 a_2840_11837.n0 a_2840_11837.t3 63.3338
R19514 a_2840_11837.n1 a_2840_11837.t1 63.3219
R19515 a_2840_11837.n0 a_2840_11837.t2 29.7268
R19516 a_4274_4943.n3 a_4274_4943.n2 647.119
R19517 a_4274_4943.n1 a_4274_4943.t4 350.253
R19518 a_4274_4943.n2 a_4274_4943.n0 260.339
R19519 a_4274_4943.n2 a_4274_4943.n1 246.119
R19520 a_4274_4943.n1 a_4274_4943.t5 189.588
R19521 a_4274_4943.n3 a_4274_4943.t3 89.1195
R19522 a_4274_4943.n0 a_4274_4943.t2 63.3338
R19523 a_4274_4943.t0 a_4274_4943.n3 41.0422
R19524 a_4274_4943.n0 a_4274_4943.t1 31.9797
R19525 a_4581_5309.t0 a_4581_5309.t1 60.0005
R19526 a_4653_5309.t0 a_4653_5309.t1 198.571
R19527 a_1651_4917.n5 a_1651_4917.n4 807.871
R19528 a_1651_4917.n0 a_1651_4917.t8 389.183
R19529 a_1651_4917.n1 a_1651_4917.n0 251.167
R19530 a_1651_4917.n1 a_1651_4917.t2 223.571
R19531 a_1651_4917.n3 a_1651_4917.t3 212.081
R19532 a_1651_4917.n2 a_1651_4917.t7 212.081
R19533 a_1651_4917.n4 a_1651_4917.n3 176.576
R19534 a_1651_4917.n0 a_1651_4917.t5 174.891
R19535 a_1651_4917.n3 a_1651_4917.t6 139.78
R19536 a_1651_4917.n2 a_1651_4917.t4 139.78
R19537 a_1651_4917.t0 a_1651_4917.n5 63.3219
R19538 a_1651_4917.n5 a_1651_4917.t1 63.3219
R19539 a_1651_4917.n3 a_1651_4917.n2 61.346
R19540 a_1651_4917.n4 a_1651_4917.n1 37.5061
R19541 SWP[8].n4 SWP[8].n3 585
R19542 SWP[8].n5 SWP[8].n4 585
R19543 SWP[8].n0 SWP[8].t5 332.312
R19544 SWP[8].n0 SWP[8].t4 295.627
R19545 SWP[8] SWP[8].n0 195.401
R19546 SWP[8].n2 SWP[8].n1 185
R19547 SWP[8] SWP[8].n2 57.7379
R19548 SWP[8] SWP[8].n7 47.8228
R19549 SWP[8].n4 SWP[8].t1 26.5955
R19550 SWP[8].n4 SWP[8].t0 26.5955
R19551 SWP[8].n7 SWP[8] 26.4614
R19552 SWP[8].n1 SWP[8].t2 24.9236
R19553 SWP[8].n1 SWP[8].t3 24.9236
R19554 SWP[8].n7 SWP[8].n6 19.8446
R19555 SWP[8].n3 SWP[8] 10.4965
R19556 SWP[8].n5 SWP[8] 10.4965
R19557 SWP[8].n3 SWP[8] 6.9125
R19558 SWP[8].n6 SWP[8] 4.3525
R19559 SWP[8].n6 SWP[8].n5 2.5605
R19560 SWP[8].n2 SWP[8] 1.7925
R19561 CKO.n42 CKO.n38 588.617
R19562 CKO CKO.n35 586.253
R19563 CKO.n35 CKO.n34 585
R19564 CKO.n41 CKO.n38 585
R19565 CKO.n28 CKO.t14 294.557
R19566 CKO.n22 CKO.t18 294.557
R19567 CKO.n19 CKO.t8 294.557
R19568 CKO.n16 CKO.t13 294.557
R19569 CKO.n13 CKO.t20 294.557
R19570 CKO.n11 CKO.t4 294.557
R19571 CKO.n8 CKO.t16 294.557
R19572 CKO.n5 CKO.t22 294.557
R19573 CKO.n2 CKO.t23 294.557
R19574 CKO.n0 CKO.t21 294.557
R19575 CKO CKO.t2 269.426
R19576 CKO CKO.t3 269.426
R19577 CKO.n28 CKO.t17 211.01
R19578 CKO.n22 CKO.t7 211.01
R19579 CKO.n19 CKO.t15 211.01
R19580 CKO.n16 CKO.t19 211.01
R19581 CKO.n13 CKO.t6 211.01
R19582 CKO.n11 CKO.t12 211.01
R19583 CKO.n8 CKO.t5 211.01
R19584 CKO.n5 CKO.t10 211.01
R19585 CKO.n2 CKO.t11 211.01
R19586 CKO.n0 CKO.t9 211.01
R19587 CKO CKO.n16 156.207
R19588 CKO CKO.n11 156.207
R19589 CKO CKO.n5 156.207
R19590 CKO CKO.n0 156.207
R19591 CKO.n29 CKO.n28 152
R19592 CKO.n23 CKO.n22 152
R19593 CKO.n20 CKO.n19 152
R19594 CKO.n14 CKO.n13 152
R19595 CKO.n9 CKO.n8 152
R19596 CKO.n3 CKO.n2 152
R19597 CKO.n35 CKO.t0 46.2955
R19598 CKO.n38 CKO.t1 46.2955
R19599 CKO.n21 CKO 22.7951
R19600 CKO.n18 CKO.n15 21.1854
R19601 CKO.n7 CKO.n4 20.5972
R19602 CKO.n25 CKO.n24 19.9901
R19603 CKO.n10 CKO 18.0246
R19604 CKO.n33 CKO 15.3605
R19605 CKO.n31 CKO.n30 14.916
R19606 CKO.n43 CKO.n42 14.916
R19607 CKO.n27 CKO.n26 14.2917
R19608 CKO CKO.n39 11.2645
R19609 CKO CKO.n20 10.4234
R19610 CKO CKO.n9 10.4234
R19611 CKO.n26 CKO.n12 10.1427
R19612 CKO.n25 CKO.n21 10.1365
R19613 CKO.n32 CKO.n1 9.66056
R19614 CKO.n10 CKO.n7 9.64748
R19615 CKO.n30 CKO 9.32621
R19616 CKO.n24 CKO 9.32621
R19617 CKO.n17 CKO 9.32621
R19618 CKO.n15 CKO 9.32621
R19619 CKO.n12 CKO 9.32621
R19620 CKO.n6 CKO 9.32621
R19621 CKO.n4 CKO 9.32621
R19622 CKO.n1 CKO 9.32621
R19623 CKO.n18 CKO.n17 9.3005
R19624 CKO.n7 CKO.n6 9.3005
R19625 CKO.n37 CKO.n36 9.3005
R19626 CKO.n32 CKO.n31 7.96341
R19627 CKO.n40 CKO 6.6565
R19628 CKO CKO.n43 6.23928
R19629 CKO.n39 CKO 6.1445
R19630 CKO.n36 CKO.n34 5.84398
R19631 CKO CKO.n37 5.1176
R19632 CKO.n39 CKO 4.63498
R19633 CKO.n40 CKO 3.61789
R19634 CKO CKO.n41 3.47876
R19635 CKO.n27 CKO.n10 3.20792
R19636 CKO.n17 CKO 3.10907
R19637 CKO.n12 CKO 3.10907
R19638 CKO.n6 CKO 3.10907
R19639 CKO.n1 CKO 3.10907
R19640 CKO.n26 CKO.n25 2.39885
R19641 CKO.n36 CKO 2.36572
R19642 CKO.n42 CKO 2.36572
R19643 CKO.n41 CKO.n40 2.36572
R19644 CKO.n33 CKO 2.0485
R19645 CKO.n21 CKO.n18 2.01939
R19646 CKO.n29 CKO 2.01193
R19647 CKO.n23 CKO 2.01193
R19648 CKO.n20 CKO 2.01193
R19649 CKO.n14 CKO 2.01193
R19650 CKO.n9 CKO 2.01193
R19651 CKO.n3 CKO 2.01193
R19652 CKO.n31 CKO.n27 1.69006
R19653 CKO.n34 CKO 1.25267
R19654 CKO CKO.n33 1.11354
R19655 CKO.n30 CKO.n29 1.09764
R19656 CKO.n24 CKO.n23 1.09764
R19657 CKO.n15 CKO.n14 1.09764
R19658 CKO.n4 CKO.n3 1.09764
R19659 CKO.n37 CKO.n32 0.479853
R19660 CKO.n43 CKO 0.162245
R19661 a_2255_5185.n1 a_2255_5185.t5 530.01
R19662 a_2255_5185.t0 a_2255_5185.n5 421.021
R19663 a_2255_5185.n0 a_2255_5185.t3 337.171
R19664 a_2255_5185.n3 a_2255_5185.t1 280.223
R19665 a_2255_5185.n4 a_2255_5185.t2 263.173
R19666 a_2255_5185.n4 a_2255_5185.t6 227.826
R19667 a_2255_5185.n0 a_2255_5185.t7 199.762
R19668 a_2255_5185.n2 a_2255_5185.n1 170.81
R19669 a_2255_5185.n2 a_2255_5185.n0 167.321
R19670 a_2255_5185.n5 a_2255_5185.n4 152
R19671 a_2255_5185.n1 a_2255_5185.t4 141.923
R19672 a_2255_5185.n3 a_2255_5185.n2 10.8376
R19673 a_2255_5185.n5 a_2255_5185.n3 2.50485
R19674 a_4145_5309.t0 a_4145_5309.t1 94.7268
R19675 a_2877_10357.n3 a_2877_10357.n2 647.119
R19676 a_2877_10357.n1 a_2877_10357.t5 350.253
R19677 a_2877_10357.n2 a_2877_10357.n0 260.339
R19678 a_2877_10357.n2 a_2877_10357.n1 246.119
R19679 a_2877_10357.n1 a_2877_10357.t4 189.588
R19680 a_2877_10357.n3 a_2877_10357.t1 89.1195
R19681 a_2877_10357.n0 a_2877_10357.t2 63.3338
R19682 a_2877_10357.t3 a_2877_10357.n3 41.0422
R19683 a_2877_10357.n0 a_2877_10357.t0 31.9797
R19684 a_2767_10383.n0 a_2767_10383.t2 1327.82
R19685 a_2767_10383.n0 a_2767_10383.t1 194.655
R19686 a_2767_10383.t0 a_2767_10383.n0 63.3219
R19687 a_1835_5461.n5 a_1835_5461.n4 807.871
R19688 a_1835_5461.n0 a_1835_5461.t8 389.183
R19689 a_1835_5461.n1 a_1835_5461.n0 251.167
R19690 a_1835_5461.n1 a_1835_5461.t2 223.571
R19691 a_1835_5461.n3 a_1835_5461.t5 212.081
R19692 a_1835_5461.n2 a_1835_5461.t3 212.081
R19693 a_1835_5461.n4 a_1835_5461.n3 176.576
R19694 a_1835_5461.n0 a_1835_5461.t4 174.891
R19695 a_1835_5461.n3 a_1835_5461.t7 139.78
R19696 a_1835_5461.n2 a_1835_5461.t6 139.78
R19697 a_1835_5461.t0 a_1835_5461.n5 63.3219
R19698 a_1835_5461.n5 a_1835_5461.t1 63.3219
R19699 a_1835_5461.n3 a_1835_5461.n2 61.346
R19700 a_1835_5461.n4 a_1835_5461.n1 37.5061
R19701 SWN[7].n4 SWN[7].n3 585
R19702 SWN[7].n3 SWN[7].n2 585
R19703 SWN[7].n1 SWN[7].n0 185
R19704 SWN[7] SWN[7].n1 49.0339
R19705 SWN[7].n3 SWN[7].t0 26.5955
R19706 SWN[7].n3 SWN[7].t1 26.5955
R19707 SWN[7].n0 SWN[7].t2 24.9236
R19708 SWN[7].n0 SWN[7].t3 24.9236
R19709 SWN[7].n2 SWN[7] 24.0039
R19710 SWN[7].n4 SWN[7] 15.6165
R19711 SWN[7].n1 SWN[7] 10.4965
R19712 SWN[7].n2 SWN[7] 1.7925
R19713 SWN[7] SWN[7].n4 1.7925
R19714 a_1467_8181.n4 a_1467_8181.n1 807.871
R19715 a_1467_8181.n0 a_1467_8181.t7 389.183
R19716 a_1467_8181.n5 a_1467_8181.n0 251.167
R19717 a_1467_8181.t0 a_1467_8181.n5 223.571
R19718 a_1467_8181.n3 a_1467_8181.t5 212.081
R19719 a_1467_8181.n2 a_1467_8181.t8 212.081
R19720 a_1467_8181.n4 a_1467_8181.n3 176.576
R19721 a_1467_8181.n0 a_1467_8181.t3 174.891
R19722 a_1467_8181.n3 a_1467_8181.t4 139.78
R19723 a_1467_8181.n2 a_1467_8181.t6 139.78
R19724 a_1467_8181.n1 a_1467_8181.t2 63.3219
R19725 a_1467_8181.n1 a_1467_8181.t1 63.3219
R19726 a_1467_8181.n3 a_1467_8181.n2 61.346
R19727 a_1467_8181.n5 a_1467_8181.n4 37.5061
R19728 a_2029_8573.t1 a_2029_8573.t0 94.7268
R19729 a_1754_9003.n3 a_1754_9003.n2 636.953
R19730 a_1754_9003.n1 a_1754_9003.t4 366.856
R19731 a_1754_9003.n2 a_1754_9003.n0 300.2
R19732 a_1754_9003.n2 a_1754_9003.n1 225.036
R19733 a_1754_9003.n1 a_1754_9003.t5 174.056
R19734 a_1754_9003.n0 a_1754_9003.t3 70.0005
R19735 a_1754_9003.t0 a_1754_9003.n3 68.0124
R19736 a_1754_9003.n3 a_1754_9003.t1 63.3219
R19737 a_1754_9003.n0 a_1754_9003.t2 61.6672
R19738 a_1467_8725.n3 a_1467_8725.n0 807.871
R19739 a_1467_8725.n4 a_1467_8725.t7 389.183
R19740 a_1467_8725.n5 a_1467_8725.n4 251.167
R19741 a_1467_8725.t0 a_1467_8725.n5 223.571
R19742 a_1467_8725.n2 a_1467_8725.t3 212.081
R19743 a_1467_8725.n1 a_1467_8725.t5 212.081
R19744 a_1467_8725.n3 a_1467_8725.n2 176.576
R19745 a_1467_8725.n4 a_1467_8725.t4 174.891
R19746 a_1467_8725.n2 a_1467_8725.t6 139.78
R19747 a_1467_8725.n1 a_1467_8725.t8 139.78
R19748 a_1467_8725.n0 a_1467_8725.t2 63.3219
R19749 a_1467_8725.n0 a_1467_8725.t1 63.3219
R19750 a_1467_8725.n2 a_1467_8725.n1 61.346
R19751 a_1467_8725.n5 a_1467_8725.n3 37.5061
R19752 a_1789_8751.t0 a_1789_8751.t1 87.1434
R19753 x3/COMP_BUF_N.n30 x3/COMP_BUF_N.t24 332.312
R19754 x3/COMP_BUF_N.n27 x3/COMP_BUF_N.t30 332.312
R19755 x3/COMP_BUF_N.n11 x3/COMP_BUF_N.t28 332.312
R19756 x3/COMP_BUF_N.n12 x3/COMP_BUF_N.t33 332.312
R19757 x3/COMP_BUF_N.n24 x3/COMP_BUF_N.t17 332.312
R19758 x3/COMP_BUF_N.n18 x3/COMP_BUF_N.t29 332.312
R19759 x3/COMP_BUF_N.n20 x3/COMP_BUF_N.t26 332.312
R19760 x3/COMP_BUF_N.n17 x3/COMP_BUF_N.t22 332.312
R19761 x3/COMP_BUF_N.n15 x3/COMP_BUF_N.t21 332.312
R19762 x3/COMP_BUF_N.n10 x3/COMP_BUF_N.t31 332.312
R19763 x3/COMP_BUF_N.n32 x3/COMP_BUF_N.n9 321.507
R19764 x3/COMP_BUF_N x3/COMP_BUF_N.n0 311.719
R19765 x3/COMP_BUF_N.n35 x3/COMP_BUF_N.n8 311.719
R19766 x3/COMP_BUF_N.n34 x3/COMP_BUF_N.n33 311.719
R19767 x3/COMP_BUF_N.n30 x3/COMP_BUF_N.t19 295.627
R19768 x3/COMP_BUF_N.n27 x3/COMP_BUF_N.t20 295.627
R19769 x3/COMP_BUF_N.n11 x3/COMP_BUF_N.t23 295.627
R19770 x3/COMP_BUF_N.n12 x3/COMP_BUF_N.t34 295.627
R19771 x3/COMP_BUF_N.n24 x3/COMP_BUF_N.t18 295.627
R19772 x3/COMP_BUF_N.n18 x3/COMP_BUF_N.t16 295.627
R19773 x3/COMP_BUF_N.n20 x3/COMP_BUF_N.t27 295.627
R19774 x3/COMP_BUF_N.n17 x3/COMP_BUF_N.t35 295.627
R19775 x3/COMP_BUF_N.n15 x3/COMP_BUF_N.t25 295.627
R19776 x3/COMP_BUF_N.n10 x3/COMP_BUF_N.t32 295.627
R19777 x3/COMP_BUF_N.n4 x3/COMP_BUF_N.n3 261.425
R19778 x3/COMP_BUF_N.n7 x3/COMP_BUF_N.n6 202.444
R19779 x3/COMP_BUF_N.n4 x3/COMP_BUF_N.n2 198.177
R19780 x3/COMP_BUF_N.n5 x3/COMP_BUF_N.n1 198.177
R19781 x3/COMP_BUF_N x3/COMP_BUF_N.n30 196.004
R19782 x3/COMP_BUF_N x3/COMP_BUF_N.n20 196.004
R19783 x3/COMP_BUF_N x3/COMP_BUF_N.n17 196.004
R19784 x3/COMP_BUF_N x3/COMP_BUF_N.n10 196.004
R19785 x3/COMP_BUF_N x3/COMP_BUF_N.n27 195.401
R19786 x3/COMP_BUF_N x3/COMP_BUF_N.n11 195.401
R19787 x3/COMP_BUF_N x3/COMP_BUF_N.n24 195.401
R19788 x3/COMP_BUF_N.n13 x3/COMP_BUF_N.n12 194.845
R19789 x3/COMP_BUF_N.n19 x3/COMP_BUF_N.n18 194.845
R19790 x3/COMP_BUF_N.n16 x3/COMP_BUF_N.n15 194.845
R19791 x3/COMP_BUF_N.n5 x3/COMP_BUF_N.n4 63.2476
R19792 x3/COMP_BUF_N.n35 x3/COMP_BUF_N.n34 63.2476
R19793 x3/COMP_BUF_N.n34 x3/COMP_BUF_N.n32 53.4593
R19794 x3/COMP_BUF_N.n7 x3/COMP_BUF_N.n5 50.4476
R19795 x3/COMP_BUF_N.n36 x3/COMP_BUF_N.n35 50.4476
R19796 x3/COMP_BUF_N.n29 x3/COMP_BUF_N 40.4559
R19797 x3/COMP_BUF_N.n23 x3/COMP_BUF_N.n16 36.5579
R19798 x3/COMP_BUF_N.n14 x3/COMP_BUF_N 32.0406
R19799 x3/COMP_BUF_N.n14 x3/COMP_BUF_N.n13 31.5531
R19800 x3/COMP_BUF_N.n21 x3/COMP_BUF_N.n19 31.4165
R19801 x3/COMP_BUF_N.n25 x3/COMP_BUF_N 30.6511
R19802 x3/COMP_BUF_N.n21 x3/COMP_BUF_N 27.2668
R19803 x3/COMP_BUF_N.n0 x3/COMP_BUF_N.t0 26.5955
R19804 x3/COMP_BUF_N.n0 x3/COMP_BUF_N.t2 26.5955
R19805 x3/COMP_BUF_N.n8 x3/COMP_BUF_N.t6 26.5955
R19806 x3/COMP_BUF_N.n8 x3/COMP_BUF_N.t3 26.5955
R19807 x3/COMP_BUF_N.n9 x3/COMP_BUF_N.t1 26.5955
R19808 x3/COMP_BUF_N.n9 x3/COMP_BUF_N.t5 26.5955
R19809 x3/COMP_BUF_N.n33 x3/COMP_BUF_N.t7 26.5955
R19810 x3/COMP_BUF_N.n33 x3/COMP_BUF_N.t4 26.5955
R19811 x3/COMP_BUF_N.n28 x3/COMP_BUF_N 25.857
R19812 x3/COMP_BUF_N.n3 x3/COMP_BUF_N.t15 24.9236
R19813 x3/COMP_BUF_N.n3 x3/COMP_BUF_N.t11 24.9236
R19814 x3/COMP_BUF_N.n2 x3/COMP_BUF_N.t13 24.9236
R19815 x3/COMP_BUF_N.n2 x3/COMP_BUF_N.t10 24.9236
R19816 x3/COMP_BUF_N.n1 x3/COMP_BUF_N.t12 24.9236
R19817 x3/COMP_BUF_N.n1 x3/COMP_BUF_N.t9 24.9236
R19818 x3/COMP_BUF_N.n6 x3/COMP_BUF_N.t14 24.9236
R19819 x3/COMP_BUF_N.n6 x3/COMP_BUF_N.t8 24.9236
R19820 x3/COMP_BUF_N.n31 x3/COMP_BUF_N 16.7737
R19821 x3/COMP_BUF_N.n29 x3/COMP_BUF_N.n28 14.8303
R19822 x3/COMP_BUF_N.n32 x3/COMP_BUF_N 14.7971
R19823 x3/COMP_BUF_N.n36 x3/COMP_BUF_N 12.8005
R19824 x3/COMP_BUF_N.n22 x3/COMP_BUF_N 12.2737
R19825 x3/COMP_BUF_N x3/COMP_BUF_N.n7 5.77305
R19826 x3/COMP_BUF_N.n31 x3/COMP_BUF_N.n29 5.63649
R19827 x3/COMP_BUF_N.n28 x3/COMP_BUF_N.n26 4.79462
R19828 x3/COMP_BUF_N.n26 x3/COMP_BUF_N.n25 4.72577
R19829 x3/COMP_BUF_N.n23 x3/COMP_BUF_N.n22 4.5005
R19830 x3/COMP_BUF_N x3/COMP_BUF_N.n36 4.26717
R19831 x3/COMP_BUF_N.n13 x3/COMP_BUF_N 4.17441
R19832 x3/COMP_BUF_N.n19 x3/COMP_BUF_N 4.17441
R19833 x3/COMP_BUF_N.n16 x3/COMP_BUF_N 4.17441
R19834 x3/COMP_BUF_N.n22 x3/COMP_BUF_N.n21 3.74363
R19835 x3/COMP_BUF_N.n26 x3/COMP_BUF_N.n14 3.21135
R19836 x3/COMP_BUF_N.n25 x3/COMP_BUF_N.n23 1.99363
R19837 x3/COMP_BUF_N x3/COMP_BUF_N.n31 0.997066
R19838 a_4779_5461.n5 a_4779_5461.n4 807.871
R19839 a_4779_5461.n0 a_4779_5461.t8 389.183
R19840 a_4779_5461.n1 a_4779_5461.n0 251.167
R19841 a_4779_5461.n1 a_4779_5461.t2 223.571
R19842 a_4779_5461.n3 a_4779_5461.t5 212.081
R19843 a_4779_5461.n2 a_4779_5461.t6 212.081
R19844 a_4779_5461.n4 a_4779_5461.n3 176.576
R19845 a_4779_5461.n0 a_4779_5461.t3 174.891
R19846 a_4779_5461.n3 a_4779_5461.t7 139.78
R19847 a_4779_5461.n2 a_4779_5461.t4 139.78
R19848 a_4779_5461.t0 a_4779_5461.n5 63.3219
R19849 a_4779_5461.n5 a_4779_5461.t1 63.3219
R19850 a_4779_5461.n3 a_4779_5461.n2 61.346
R19851 a_4779_5461.n4 a_4779_5461.n1 37.5061
R19852 a_5341_5487.n0 a_5341_5487.t0 68.3338
R19853 a_5341_5487.n0 a_5341_5487.t1 26.3935
R19854 a_5341_5487.n1 a_5341_5487.n0 14.4005
R19855 a_5040_10383.n0 a_5040_10383.t2 1327.82
R19856 a_5040_10383.n0 a_5040_10383.t1 194.655
R19857 a_5040_10383.t0 a_5040_10383.n0 63.3219
R19858 a_4895_10357.n3 a_4895_10357.n2 674.338
R19859 a_4895_10357.n1 a_4895_10357.t4 332.58
R19860 a_4895_10357.n2 a_4895_10357.n0 284.012
R19861 a_4895_10357.n2 a_4895_10357.n1 253.648
R19862 a_4895_10357.n1 a_4895_10357.t5 168.701
R19863 a_4895_10357.t0 a_4895_10357.n3 96.1553
R19864 a_4895_10357.n3 a_4895_10357.t3 65.6672
R19865 a_4895_10357.n0 a_4895_10357.t1 65.0005
R19866 a_4895_10357.n0 a_4895_10357.t2 45.0005
R19867 a_10281_4221.t0 a_10281_4221.t1 60.0005
R19868 a_6803_2741.n5 a_6803_2741.n4 807.871
R19869 a_6803_2741.n0 a_6803_2741.t6 389.183
R19870 a_6803_2741.n1 a_6803_2741.n0 251.167
R19871 a_6803_2741.n1 a_6803_2741.t1 223.571
R19872 a_6803_2741.n3 a_6803_2741.t7 212.081
R19873 a_6803_2741.n2 a_6803_2741.t3 212.081
R19874 a_6803_2741.n4 a_6803_2741.n3 176.576
R19875 a_6803_2741.n0 a_6803_2741.t4 174.891
R19876 a_6803_2741.n3 a_6803_2741.t5 139.78
R19877 a_6803_2741.n2 a_6803_2741.t8 139.78
R19878 a_6803_2741.t0 a_6803_2741.n5 63.3219
R19879 a_6803_2741.n5 a_6803_2741.t2 63.3219
R19880 a_6803_2741.n3 a_6803_2741.n2 61.346
R19881 a_6803_2741.n4 a_6803_2741.n1 37.5061
R19882 a_8951_8751.n1 a_8951_8751.t2 530.01
R19883 a_8951_8751.t0 a_8951_8751.n5 421.021
R19884 a_8951_8751.n0 a_8951_8751.t4 337.142
R19885 a_8951_8751.n3 a_8951_8751.t1 280.223
R19886 a_8951_8751.n4 a_8951_8751.t5 263.173
R19887 a_8951_8751.n4 a_8951_8751.t6 227.826
R19888 a_8951_8751.n0 a_8951_8751.t7 199.762
R19889 a_8951_8751.n2 a_8951_8751.n1 170.81
R19890 a_8951_8751.n2 a_8951_8751.n0 167.321
R19891 a_8951_8751.n5 a_8951_8751.n4 152
R19892 a_8951_8751.n1 a_8951_8751.t3 141.923
R19893 a_8951_8751.n3 a_8951_8751.n2 10.8376
R19894 a_8951_8751.n5 a_8951_8751.n3 2.50485
R19895 a_4515_12381.n0 a_4515_12381.t2 1327.82
R19896 a_4515_12381.t0 a_4515_12381.n0 194.655
R19897 a_4515_12381.n0 a_4515_12381.t1 63.3219
R19898 a_5307_7093.n22 a_5307_7093.t5 286.348
R19899 a_5307_7093.n24 a_5307_7093.t0 271.051
R19900 a_5307_7093.n1 a_5307_7093.t20 221.72
R19901 a_5307_7093.n18 a_5307_7093.t10 221.72
R19902 a_5307_7093.n2 a_5307_7093.t16 221.72
R19903 a_5307_7093.n12 a_5307_7093.t12 221.72
R19904 a_5307_7093.n10 a_5307_7093.t18 221.72
R19905 a_5307_7093.n4 a_5307_7093.t14 221.72
R19906 a_5307_7093.n6 a_5307_7093.t8 221.72
R19907 a_5307_7093.n5 a_5307_7093.t9 221.72
R19908 a_5307_7093.n25 a_5307_7093.n24 206.055
R19909 a_5307_7093.n22 a_5307_7093.n21 198.177
R19910 a_5307_7093.n8 a_5307_7093.n7 177.601
R19911 a_5307_7093.n9 a_5307_7093.n8 152
R19912 a_5307_7093.n11 a_5307_7093.n3 152
R19913 a_5307_7093.n14 a_5307_7093.n13 152
R19914 a_5307_7093.n16 a_5307_7093.n15 152
R19915 a_5307_7093.n17 a_5307_7093.n0 152
R19916 a_5307_7093.n20 a_5307_7093.n19 152
R19917 a_5307_7093.n1 a_5307_7093.t15 149.421
R19918 a_5307_7093.n18 a_5307_7093.t21 149.421
R19919 a_5307_7093.n2 a_5307_7093.t11 149.421
R19920 a_5307_7093.n12 a_5307_7093.t6 149.421
R19921 a_5307_7093.n10 a_5307_7093.t13 149.421
R19922 a_5307_7093.n4 a_5307_7093.t7 149.421
R19923 a_5307_7093.n6 a_5307_7093.t17 149.421
R19924 a_5307_7093.n5 a_5307_7093.t19 149.421
R19925 a_5307_7093.n6 a_5307_7093.n5 74.9783
R19926 a_5307_7093.n7 a_5307_7093.n6 66.0523
R19927 a_5307_7093.n17 a_5307_7093.n16 60.6968
R19928 a_5307_7093.n19 a_5307_7093.n18 55.3412
R19929 a_5307_7093.n13 a_5307_7093.n2 51.7709
R19930 a_5307_7093.n9 a_5307_7093.n4 51.7709
R19931 a_5307_7093.n23 a_5307_7093.n22 48.9632
R19932 a_5307_7093.n24 a_5307_7093.n23 38.7339
R19933 a_5307_7093.n12 a_5307_7093.n11 37.4894
R19934 a_5307_7093.n11 a_5307_7093.n10 37.4894
R19935 a_5307_7093.t2 a_5307_7093.n25 26.5955
R19936 a_5307_7093.n25 a_5307_7093.t1 26.5955
R19937 a_5307_7093.n20 a_5307_7093.n0 25.6005
R19938 a_5307_7093.n15 a_5307_7093.n0 25.6005
R19939 a_5307_7093.n15 a_5307_7093.n14 25.6005
R19940 a_5307_7093.n14 a_5307_7093.n3 25.6005
R19941 a_5307_7093.n8 a_5307_7093.n3 25.6005
R19942 a_5307_7093.n21 a_5307_7093.t4 24.9236
R19943 a_5307_7093.n21 a_5307_7093.t3 24.9236
R19944 a_5307_7093.n13 a_5307_7093.n12 23.2079
R19945 a_5307_7093.n10 a_5307_7093.n9 23.2079
R19946 a_5307_7093.n19 a_5307_7093.n1 19.6375
R19947 a_5307_7093.n23 a_5307_7093.n20 18.4476
R19948 a_5307_7093.n16 a_5307_7093.n2 8.92643
R19949 a_5307_7093.n7 a_5307_7093.n4 8.92643
R19950 a_5307_7093.n18 a_5307_7093.n17 5.35606
R19951 FINAL.n9 FINAL.n2 321.507
R19952 FINAL.n11 FINAL.n0 311.719
R19953 FINAL.n10 FINAL.n1 311.719
R19954 FINAL FINAL.n20 311.719
R19955 FINAL.n15 FINAL.n14 261.425
R19956 FINAL.n6 FINAL.t18 256.07
R19957 FINAL.n3 FINAL.t17 256.07
R19958 FINAL.n18 FINAL.n17 202.444
R19959 FINAL.n15 FINAL.n13 198.177
R19960 FINAL.n16 FINAL.n12 198.177
R19961 FINAL.n7 FINAL.n6 152
R19962 FINAL.n4 FINAL.n3 152
R19963 FINAL.n6 FINAL.t16 150.03
R19964 FINAL.n3 FINAL.t19 150.03
R19965 FINAL.n16 FINAL.n15 63.2476
R19966 FINAL.n11 FINAL.n10 63.2476
R19967 FINAL.n10 FINAL.n9 53.4593
R19968 FINAL.n18 FINAL.n16 50.4476
R19969 FINAL.n19 FINAL.n11 50.4476
R19970 FINAL.n8 FINAL.n5 37.3488
R19971 FINAL.n0 FINAL.t1 26.5955
R19972 FINAL.n0 FINAL.t3 26.5955
R19973 FINAL.n1 FINAL.t2 26.5955
R19974 FINAL.n1 FINAL.t4 26.5955
R19975 FINAL.n2 FINAL.t0 26.5955
R19976 FINAL.n2 FINAL.t5 26.5955
R19977 FINAL.n20 FINAL.t7 26.5955
R19978 FINAL.n20 FINAL.t6 26.5955
R19979 FINAL.n14 FINAL.t11 24.9236
R19980 FINAL.n14 FINAL.t8 24.9236
R19981 FINAL.n13 FINAL.t13 24.9236
R19982 FINAL.n13 FINAL.t15 24.9236
R19983 FINAL.n12 FINAL.t12 24.9236
R19984 FINAL.n12 FINAL.t14 24.9236
R19985 FINAL.n17 FINAL.t10 24.9236
R19986 FINAL.n17 FINAL.t9 24.9236
R19987 FINAL.n8 FINAL 21.6175
R19988 FINAL.n9 FINAL 15.4106
R19989 FINAL.n19 FINAL 12.8005
R19990 FINAL FINAL.n7 8.23114
R19991 FINAL.n7 FINAL 7.6805
R19992 FINAL.n4 FINAL 7.6805
R19993 FINAL FINAL.n8 6.09528
R19994 FINAL FINAL.n18 5.77305
R19995 FINAL.n5 FINAL.n4 4.6085
R19996 FINAL.n5 FINAL 4.58918
R19997 FINAL FINAL.n19 4.26717
R19998 SWP[0].n4 SWP[0].n3 585
R19999 SWP[0].n5 SWP[0].n4 585
R20000 SWP[0].n0 SWP[0].t5 333.651
R20001 SWP[0].n0 SWP[0].t4 297.233
R20002 SWP[0].n8 SWP[0].n0 195.701
R20003 SWP[0].n2 SWP[0].n1 185
R20004 SWP[0] SWP[0].n2 57.7379
R20005 SWP[0].n8 SWP[0].n7 38.0426
R20006 SWP[0].n4 SWP[0].t0 26.5955
R20007 SWP[0].n4 SWP[0].t1 26.5955
R20008 SWP[0].n1 SWP[0].t2 24.9236
R20009 SWP[0].n1 SWP[0].t3 24.9236
R20010 SWP[0].n7 SWP[0] 17.8184
R20011 SWP[0].n3 SWP[0] 10.4965
R20012 SWP[0].n5 SWP[0] 10.4965
R20013 SWP[0].n7 SWP[0].n6 9.3005
R20014 SWP[0].n3 SWP[0] 6.9125
R20015 SWP[0].n6 SWP[0] 4.3525
R20016 SWP[0].n6 SWP[0].n5 2.5605
R20017 SWP[0].n2 SWP[0] 1.7925
R20018 SWP[0] SWP[0].n8 1.03669
R20019 a_9832_9661.n1 a_9832_9661.n0 926.024
R20020 a_9832_9661.t0 a_9832_9661.n1 82.0838
R20021 a_9832_9661.n0 a_9832_9661.t1 63.3338
R20022 a_9832_9661.n1 a_9832_9661.t2 63.3219
R20023 a_9832_9661.n0 a_9832_9661.t3 29.7268
R20024 a_5960_3677.t0 a_5960_3677.n0 1327.82
R20025 a_5960_3677.n0 a_5960_3677.t1 194.655
R20026 a_5960_3677.n0 a_5960_3677.t2 63.3219
R20027 a_8262_6031.t0 a_8262_6031.t1 126.644
R20028 a_3767_8181.n5 a_3767_8181.n4 807.871
R20029 a_3767_8181.n0 a_3767_8181.t4 389.183
R20030 a_3767_8181.n1 a_3767_8181.n0 251.167
R20031 a_3767_8181.n1 a_3767_8181.t1 223.571
R20032 a_3767_8181.n3 a_3767_8181.t7 212.081
R20033 a_3767_8181.n2 a_3767_8181.t3 212.081
R20034 a_3767_8181.n4 a_3767_8181.n3 176.576
R20035 a_3767_8181.n0 a_3767_8181.t6 174.891
R20036 a_3767_8181.n3 a_3767_8181.t5 139.78
R20037 a_3767_8181.n2 a_3767_8181.t8 139.78
R20038 a_3767_8181.t0 a_3767_8181.n5 63.3219
R20039 a_3767_8181.n5 a_3767_8181.t2 63.3219
R20040 a_3767_8181.n3 a_3767_8181.n2 61.346
R20041 a_3767_8181.n4 a_3767_8181.n1 37.5061
R20042 SWN[5].n2 SWN[5].n1 585
R20043 SWN[5].n1 SWN[5].n0 585
R20044 SWN[5].n4 SWN[5].n3 185
R20045 SWN[5].n4 SWN[5] 57.7379
R20046 SWN[5].n1 SWN[5].t0 26.5955
R20047 SWN[5].n1 SWN[5].t1 26.5955
R20048 SWN[5].n3 SWN[5].t3 24.9236
R20049 SWN[5].n3 SWN[5].t2 24.9236
R20050 SWN[5] SWN[5].n2 10.4965
R20051 SWN[5].n0 SWN[5] 10.4965
R20052 SWN[5].n2 SWN[5] 6.9125
R20053 SWN[5].n0 SWN[5] 6.9125
R20054 SWN[5] SWN[5].n4 1.7925
R20055 x2/net5.n5 x2/net5.n4 585
R20056 x2/net5.n4 x2/net5.n3 585
R20057 x2/net5.n0 x2/net5.t4 333.651
R20058 x2/net5.n0 x2/net5.t5 297.233
R20059 x2/net5 x2/net5.n0 195.701
R20060 x2/net5.n2 x2/net5.n1 185
R20061 x2/net5 x2/net5.n2 57.7379
R20062 x2/net5.n4 x2/net5.t1 26.5955
R20063 x2/net5.n4 x2/net5.t0 26.5955
R20064 x2/net5.n1 x2/net5.t3 24.9236
R20065 x2/net5.n1 x2/net5.t2 24.9236
R20066 x2/net5 x2/net5.n5 10.4965
R20067 x2/net5.n3 x2/net5 10.4965
R20068 x2/net5.n5 x2/net5 6.9125
R20069 x2/net5.n3 x2/net5 6.9125
R20070 x2/net5.n2 x2/net5 1.7925
R20071 a_9372_10927.n1 a_9372_10927.n0 926.024
R20072 a_9372_10927.t0 a_9372_10927.n1 82.0838
R20073 a_9372_10927.n0 a_9372_10927.t3 63.3338
R20074 a_9372_10927.n1 a_9372_10927.t1 63.3219
R20075 a_9372_10927.n0 a_9372_10927.t2 29.7268
R20076 SWN[6].n2 SWN[6] 586.793
R20077 SWN[6].n3 SWN[6].n2 585
R20078 SWN[6].n1 SWN[6].n0 185
R20079 SWN[6] SWN[6].n1 49.0339
R20080 SWN[6].n2 SWN[6].t1 26.5955
R20081 SWN[6].n2 SWN[6].t0 26.5955
R20082 SWN[6].n0 SWN[6].t2 24.9236
R20083 SWN[6].n0 SWN[6].t3 24.9236
R20084 SWN[6].n4 SWN[6] 16.8462
R20085 SWN[6].n3 SWN[6] 15.6165
R20086 SWN[6].n4 SWN[6] 13.0565
R20087 SWN[6].n1 SWN[6] 10.4965
R20088 SWN[6] SWN[6].n4 4.3525
R20089 SWN[6] SWN[6].n3 1.7925
R20090 a_9117_8751.t0 a_9117_8751.n3 370.026
R20091 a_9117_8751.n0 a_9117_8751.t2 351.356
R20092 a_9117_8751.n1 a_9117_8751.t5 334.717
R20093 a_9117_8751.n3 a_9117_8751.t1 325.971
R20094 a_9117_8751.n1 a_9117_8751.t3 309.935
R20095 a_9117_8751.n0 a_9117_8751.t4 305.683
R20096 a_9117_8751.n2 a_9117_8751.n0 16.879
R20097 a_9117_8751.n3 a_9117_8751.n2 10.8867
R20098 a_9117_8751.n2 a_9117_8751.n1 9.3005
R20099 a_9685_8993.n3 a_9685_8993.n2 647.119
R20100 a_9685_8993.n1 a_9685_8993.t4 350.253
R20101 a_9685_8993.n2 a_9685_8993.n0 260.339
R20102 a_9685_8993.n2 a_9685_8993.n1 246.119
R20103 a_9685_8993.n1 a_9685_8993.t5 189.588
R20104 a_9685_8993.n3 a_9685_8993.t2 89.1195
R20105 a_9685_8993.n0 a_9685_8993.t0 63.3338
R20106 a_9685_8993.t1 a_9685_8993.n3 41.0422
R20107 a_9685_8993.n0 a_9685_8993.t3 31.9797
R20108 a_10032_8751.n3 a_10032_8751.n2 636.953
R20109 a_10032_8751.n1 a_10032_8751.t5 366.856
R20110 a_10032_8751.n2 a_10032_8751.n0 300.2
R20111 a_10032_8751.n2 a_10032_8751.n1 225.036
R20112 a_10032_8751.n1 a_10032_8751.t4 174.056
R20113 a_10032_8751.n0 a_10032_8751.t1 70.0005
R20114 a_10032_8751.n3 a_10032_8751.t3 68.0124
R20115 a_10032_8751.t0 a_10032_8751.n3 63.3219
R20116 a_10032_8751.n0 a_10032_8751.t2 61.6672
R20117 a_9685_7905.n3 a_9685_7905.n2 647.119
R20118 a_9685_7905.n1 a_9685_7905.t4 350.253
R20119 a_9685_7905.n2 a_9685_7905.n0 260.339
R20120 a_9685_7905.n2 a_9685_7905.n1 246.119
R20121 a_9685_7905.n1 a_9685_7905.t5 189.588
R20122 a_9685_7905.n3 a_9685_7905.t1 89.1195
R20123 a_9685_7905.n0 a_9685_7905.t0 63.3338
R20124 a_9685_7905.t2 a_9685_7905.n3 41.0422
R20125 a_9685_7905.n0 a_9685_7905.t3 31.9797
R20126 a_2779_6005.n3 a_2779_6005.n2 674.338
R20127 a_2779_6005.n1 a_2779_6005.t4 332.58
R20128 a_2779_6005.n2 a_2779_6005.n0 284.012
R20129 a_2779_6005.n2 a_2779_6005.n1 253.648
R20130 a_2779_6005.n1 a_2779_6005.t5 168.701
R20131 a_2779_6005.t0 a_2779_6005.n3 96.1553
R20132 a_2779_6005.n3 a_2779_6005.t3 65.6672
R20133 a_2779_6005.n0 a_2779_6005.t1 65.0005
R20134 a_2779_6005.n0 a_2779_6005.t2 45.0005
R20135 a_3342_6031.n1 a_3342_6031.n0 926.024
R20136 a_3342_6031.n1 a_3342_6031.t3 82.0838
R20137 a_3342_6031.n0 a_3342_6031.t0 63.3338
R20138 a_3342_6031.t1 a_3342_6031.n1 63.3219
R20139 a_3342_6031.n0 a_3342_6031.t2 29.7268
R20140 a_5915_7663.n1 a_5915_7663.t3 530.01
R20141 a_5915_7663.t0 a_5915_7663.n5 421.021
R20142 a_5915_7663.n0 a_5915_7663.t7 337.142
R20143 a_5915_7663.n3 a_5915_7663.t1 280.223
R20144 a_5915_7663.n4 a_5915_7663.t6 263.173
R20145 a_5915_7663.n4 a_5915_7663.t2 227.826
R20146 a_5915_7663.n0 a_5915_7663.t4 199.762
R20147 a_5915_7663.n2 a_5915_7663.n1 170.81
R20148 a_5915_7663.n2 a_5915_7663.n0 167.321
R20149 a_5915_7663.n5 a_5915_7663.n4 152
R20150 a_5915_7663.n1 a_5915_7663.t5 141.923
R20151 a_5915_7663.n3 a_5915_7663.n2 10.8376
R20152 a_5915_7663.n5 a_5915_7663.n3 2.50485
R20153 a_6081_7663.t0 a_6081_7663.n3 370.026
R20154 a_6081_7663.n0 a_6081_7663.t2 351.356
R20155 a_6081_7663.n1 a_6081_7663.t3 334.717
R20156 a_6081_7663.n3 a_6081_7663.t1 325.971
R20157 a_6081_7663.n1 a_6081_7663.t4 309.935
R20158 a_6081_7663.n0 a_6081_7663.t5 305.683
R20159 a_6081_7663.n2 a_6081_7663.n0 16.879
R20160 a_6081_7663.n3 a_6081_7663.n2 10.8867
R20161 a_6081_7663.n2 a_6081_7663.n1 9.3005
R20162 a_7093_10927.t1 a_7093_10927.n3 370.026
R20163 a_7093_10927.n0 a_7093_10927.t2 351.356
R20164 a_7093_10927.n1 a_7093_10927.t4 334.717
R20165 a_7093_10927.n3 a_7093_10927.t0 325.971
R20166 a_7093_10927.n1 a_7093_10927.t5 309.935
R20167 a_7093_10927.n0 a_7093_10927.t3 305.683
R20168 a_7093_10927.n2 a_7093_10927.n0 16.879
R20169 a_7093_10927.n3 a_7093_10927.n2 10.8867
R20170 a_7093_10927.n2 a_7093_10927.n1 9.3005
R20171 a_7661_11169.n3 a_7661_11169.n2 647.119
R20172 a_7661_11169.n1 a_7661_11169.t5 350.253
R20173 a_7661_11169.n2 a_7661_11169.n0 260.339
R20174 a_7661_11169.n2 a_7661_11169.n1 246.119
R20175 a_7661_11169.n1 a_7661_11169.t4 189.588
R20176 a_7661_11169.n3 a_7661_11169.t2 89.1195
R20177 a_7661_11169.n0 a_7661_11169.t3 63.3338
R20178 a_7661_11169.t0 a_7661_11169.n3 41.0422
R20179 a_7661_11169.n0 a_7661_11169.t1 31.9797
R20180 a_9372_8751.n1 a_9372_8751.n0 926.024
R20181 a_9372_8751.t0 a_9372_8751.n1 82.0838
R20182 a_9372_8751.n0 a_9372_8751.t1 63.3338
R20183 a_9372_8751.n1 a_9372_8751.t3 63.3219
R20184 a_9372_8751.n0 a_9372_8751.t2 29.7268
R20185 a_9467_8751.n3 a_9467_8751.n2 674.338
R20186 a_9467_8751.n1 a_9467_8751.t4 332.58
R20187 a_9467_8751.n2 a_9467_8751.n0 284.012
R20188 a_9467_8751.n2 a_9467_8751.n1 253.648
R20189 a_9467_8751.n1 a_9467_8751.t5 168.701
R20190 a_9467_8751.n3 a_9467_8751.t2 96.1553
R20191 a_9467_8751.t1 a_9467_8751.n3 65.6672
R20192 a_9467_8751.n0 a_9467_8751.t3 65.0005
R20193 a_9467_8751.n0 a_9467_8751.t0 45.0005
R20194 a_4407_12015.n3 a_4407_12015.n2 674.338
R20195 a_4407_12015.n1 a_4407_12015.t4 332.58
R20196 a_4407_12015.n2 a_4407_12015.n0 284.012
R20197 a_4407_12015.n2 a_4407_12015.n1 253.648
R20198 a_4407_12015.n1 a_4407_12015.t5 168.701
R20199 a_4407_12015.t0 a_4407_12015.n3 96.1553
R20200 a_4407_12015.n3 a_4407_12015.t1 65.6672
R20201 a_4407_12015.n0 a_4407_12015.t2 65.0005
R20202 a_4407_12015.n0 a_4407_12015.t3 45.0005
R20203 a_4625_12257.n3 a_4625_12257.n2 647.119
R20204 a_4625_12257.n1 a_4625_12257.t5 350.253
R20205 a_4625_12257.n2 a_4625_12257.n0 260.339
R20206 a_4625_12257.n2 a_4625_12257.n1 246.119
R20207 a_4625_12257.n1 a_4625_12257.t4 189.588
R20208 a_4625_12257.n3 a_4625_12257.t1 89.1195
R20209 a_4625_12257.n0 a_4625_12257.t0 63.3338
R20210 a_4625_12257.t2 a_4625_12257.n3 41.0422
R20211 a_4625_12257.n0 a_4625_12257.t3 31.9797
R20212 a_3399_10687.n5 a_3399_10687.n4 807.871
R20213 a_3399_10687.n2 a_3399_10687.t5 389.183
R20214 a_3399_10687.n3 a_3399_10687.n2 251.167
R20215 a_3399_10687.n3 a_3399_10687.t1 223.571
R20216 a_3399_10687.n0 a_3399_10687.t7 212.081
R20217 a_3399_10687.n1 a_3399_10687.t8 212.081
R20218 a_3399_10687.n4 a_3399_10687.n1 176.576
R20219 a_3399_10687.n2 a_3399_10687.t6 174.891
R20220 a_3399_10687.n0 a_3399_10687.t3 139.78
R20221 a_3399_10687.n1 a_3399_10687.t4 139.78
R20222 a_3399_10687.t0 a_3399_10687.n5 63.3219
R20223 a_3399_10687.n5 a_3399_10687.t2 63.3219
R20224 a_3399_10687.n1 a_3399_10687.n0 61.346
R20225 a_3399_10687.n4 a_3399_10687.n3 37.7195
R20226 x2/net6.n9 x2/net6.n8 585
R20227 x2/net6.n10 x2/net6.n9 585
R20228 x2/net6.n2 x2/net6.t9 332.312
R20229 x2/net6.n2 x2/net6.t6 295.627
R20230 x2/net6.n4 x2/net6.t4 212.081
R20231 x2/net6.n3 x2/net6.t5 212.081
R20232 x2/net6 x2/net6.n2 196.004
R20233 x2/net6.n1 x2/net6.n0 185
R20234 x2/net6.n5 x2/net6.n4 182.673
R20235 x2/net6.n4 x2/net6.t7 139.78
R20236 x2/net6.n3 x2/net6.t8 139.78
R20237 x2/net6.n4 x2/net6.n3 61.346
R20238 x2/net6.n7 x2/net6.n1 53.3859
R20239 x2/net6.n9 x2/net6.t1 26.5955
R20240 x2/net6.n9 x2/net6.t0 26.5955
R20241 x2/net6.n0 x2/net6.t3 24.9236
R20242 x2/net6.n0 x2/net6.t2 24.9236
R20243 x2/net6.n6 x2/net6.n5 22.6452
R20244 x2/net6.n7 x2/net6 13.1516
R20245 x2/net6.n6 x2/net6 12.6844
R20246 x2/net6.n8 x2/net6 10.4965
R20247 x2/net6.n10 x2/net6 10.4965
R20248 x2/net6.n8 x2/net6 6.9125
R20249 x2/net6 x2/net6.n10 6.9125
R20250 x2/net6 x2/net6.n7 4.3525
R20251 x2/net6.n5 x2/net6 2.3045
R20252 x2/net6.n1 x2/net6 1.7925
R20253 x2/net6 x2/net6.n6 1.37207
R20254 a_5734_2767.n1 a_5734_2767.n0 926.024
R20255 a_5734_2767.n1 a_5734_2767.t3 82.0838
R20256 a_5734_2767.n0 a_5734_2767.t2 63.3338
R20257 a_5734_2767.t0 a_5734_2767.n1 63.3219
R20258 a_5734_2767.n0 a_5734_2767.t1 29.7268
R20259 a_4187_5185.n1 a_4187_5185.t2 530.01
R20260 a_4187_5185.t0 a_4187_5185.n5 421.021
R20261 a_4187_5185.n0 a_4187_5185.t6 337.171
R20262 a_4187_5185.n3 a_4187_5185.t1 280.223
R20263 a_4187_5185.n4 a_4187_5185.t5 263.173
R20264 a_4187_5185.n4 a_4187_5185.t3 227.826
R20265 a_4187_5185.n0 a_4187_5185.t4 199.762
R20266 a_4187_5185.n2 a_4187_5185.n1 170.81
R20267 a_4187_5185.n2 a_4187_5185.n0 167.321
R20268 a_4187_5185.n5 a_4187_5185.n4 152
R20269 a_4187_5185.n1 a_4187_5185.t7 141.923
R20270 a_4187_5185.n3 a_4187_5185.n2 10.8376
R20271 a_4187_5185.n5 a_4187_5185.n3 2.50485
R20272 a_4488_4943.t0 a_4488_4943.n0 1327.82
R20273 a_4488_4943.n0 a_4488_4943.t2 194.655
R20274 a_4488_4943.n0 a_4488_4943.t1 63.3219
R20275 a_4343_4917.n3 a_4343_4917.n2 674.338
R20276 a_4343_4917.n1 a_4343_4917.t5 332.58
R20277 a_4343_4917.n2 a_4343_4917.n0 284.012
R20278 a_4343_4917.n2 a_4343_4917.n1 253.648
R20279 a_4343_4917.n1 a_4343_4917.t4 168.701
R20280 a_4343_4917.n3 a_4343_4917.t1 96.1553
R20281 a_4343_4917.t0 a_4343_4917.n3 65.6672
R20282 a_4343_4917.n0 a_4343_4917.t2 65.0005
R20283 a_4343_4917.n0 a_4343_4917.t3 45.0005
R20284 a_8197_10389.t0 a_8197_10389.n3 370.026
R20285 a_8197_10389.n0 a_8197_10389.t5 351.356
R20286 a_8197_10389.n1 a_8197_10389.t3 334.717
R20287 a_8197_10389.n3 a_8197_10389.t1 325.971
R20288 a_8197_10389.n1 a_8197_10389.t4 309.935
R20289 a_8197_10389.n0 a_8197_10389.t2 305.683
R20290 a_8197_10389.n2 a_8197_10389.n0 16.879
R20291 a_8197_10389.n3 a_8197_10389.n2 10.8867
R20292 a_8197_10389.n2 a_8197_10389.n1 9.3005
R20293 a_9112_10761.n3 a_9112_10761.n2 636.953
R20294 a_9112_10761.n1 a_9112_10761.t5 366.856
R20295 a_9112_10761.n2 a_9112_10761.n0 300.2
R20296 a_9112_10761.n2 a_9112_10761.n1 225.036
R20297 a_9112_10761.n1 a_9112_10761.t4 174.056
R20298 a_9112_10761.n0 a_9112_10761.t2 70.0005
R20299 a_9112_10761.t1 a_9112_10761.n3 68.0124
R20300 a_9112_10761.n3 a_9112_10761.t3 63.3219
R20301 a_9112_10761.n0 a_9112_10761.t0 61.6672
R20302 a_9274_10383.t0 a_9274_10383.t1 126.644
R20303 a_8284_4233.n3 a_8284_4233.n2 636.953
R20304 a_8284_4233.n1 a_8284_4233.t4 366.856
R20305 a_8284_4233.n2 a_8284_4233.n0 300.2
R20306 a_8284_4233.n2 a_8284_4233.n1 225.036
R20307 a_8284_4233.n1 a_8284_4233.t5 174.056
R20308 a_8284_4233.n0 a_8284_4233.t0 70.0005
R20309 a_8284_4233.n3 a_8284_4233.t3 68.0124
R20310 a_8284_4233.t2 a_8284_4233.n3 63.3219
R20311 a_8284_4233.n0 a_8284_4233.t1 61.6672
R20312 a_9595_5487.n1 a_9595_5487.t7 530.01
R20313 a_9595_5487.t0 a_9595_5487.n5 421.021
R20314 a_9595_5487.n0 a_9595_5487.t3 337.142
R20315 a_9595_5487.n3 a_9595_5487.t1 280.223
R20316 a_9595_5487.n4 a_9595_5487.t6 263.173
R20317 a_9595_5487.n4 a_9595_5487.t4 227.826
R20318 a_9595_5487.n0 a_9595_5487.t5 199.762
R20319 a_9595_5487.n2 a_9595_5487.n1 170.81
R20320 a_9595_5487.n2 a_9595_5487.n0 167.321
R20321 a_9595_5487.n5 a_9595_5487.n4 152
R20322 a_9595_5487.n1 a_9595_5487.t2 141.923
R20323 a_9595_5487.n3 a_9595_5487.n2 10.8376
R20324 a_9595_5487.n5 a_9595_5487.n3 2.50485
R20325 a_10016_5487.n1 a_10016_5487.n0 926.024
R20326 a_10016_5487.t0 a_10016_5487.n1 82.0838
R20327 a_10016_5487.n0 a_10016_5487.t3 63.3338
R20328 a_10016_5487.n1 a_10016_5487.t1 63.3219
R20329 a_10016_5487.n0 a_10016_5487.t2 29.7268
R20330 a_10111_5487.n3 a_10111_5487.n2 674.338
R20331 a_10111_5487.n1 a_10111_5487.t4 332.58
R20332 a_10111_5487.n2 a_10111_5487.n0 284.012
R20333 a_10111_5487.n2 a_10111_5487.n1 253.648
R20334 a_10111_5487.n1 a_10111_5487.t5 168.701
R20335 a_10111_5487.n3 a_10111_5487.t2 96.1553
R20336 a_10111_5487.t1 a_10111_5487.n3 65.6672
R20337 a_10111_5487.n0 a_10111_5487.t3 65.0005
R20338 a_10111_5487.n0 a_10111_5487.t0 45.0005
R20339 a_10676_5487.n3 a_10676_5487.n2 636.953
R20340 a_10676_5487.n1 a_10676_5487.t5 366.856
R20341 a_10676_5487.n2 a_10676_5487.n0 300.2
R20342 a_10676_5487.n2 a_10676_5487.n1 225.036
R20343 a_10676_5487.n1 a_10676_5487.t4 174.056
R20344 a_10676_5487.n0 a_10676_5487.t1 70.0005
R20345 a_10676_5487.n3 a_10676_5487.t2 68.0124
R20346 a_10676_5487.t0 a_10676_5487.n3 63.3219
R20347 a_10676_5487.n0 a_10676_5487.t3 61.6672
R20348 a_10768_6575.n3 a_10768_6575.n2 636.953
R20349 a_10768_6575.n1 a_10768_6575.t5 366.856
R20350 a_10768_6575.n2 a_10768_6575.n0 300.2
R20351 a_10768_6575.n2 a_10768_6575.n1 225.036
R20352 a_10768_6575.n1 a_10768_6575.t4 174.056
R20353 a_10768_6575.n0 a_10768_6575.t2 70.0005
R20354 a_10768_6575.t1 a_10768_6575.n3 68.0124
R20355 a_10768_6575.n3 a_10768_6575.t3 63.3219
R20356 a_10768_6575.n0 a_10768_6575.t0 61.6672
R20357 a_10877_6575.t1 a_10877_6575.t0 94.7268
R20358 a_10667_9599.n4 a_10667_9599.n1 807.871
R20359 a_10667_9599.n0 a_10667_9599.t5 389.183
R20360 a_10667_9599.n5 a_10667_9599.n0 251.167
R20361 a_10667_9599.t0 a_10667_9599.n5 223.571
R20362 a_10667_9599.n2 a_10667_9599.t8 212.081
R20363 a_10667_9599.n3 a_10667_9599.t4 212.081
R20364 a_10667_9599.n4 a_10667_9599.n3 176.576
R20365 a_10667_9599.n0 a_10667_9599.t6 174.891
R20366 a_10667_9599.n2 a_10667_9599.t3 139.78
R20367 a_10667_9599.n3 a_10667_9599.t7 139.78
R20368 a_10667_9599.n1 a_10667_9599.t1 63.3219
R20369 a_10667_9599.n1 a_10667_9599.t2 63.3219
R20370 a_10667_9599.n3 a_10667_9599.n2 61.346
R20371 a_10667_9599.n5 a_10667_9599.n4 37.7195
R20372 DOUT[0].n4 DOUT[0].n3 585
R20373 DOUT[0].n3 DOUT[0].n2 585
R20374 DOUT[0].n1 DOUT[0].n0 185
R20375 DOUT[0].n5 DOUT[0].n1 53.3859
R20376 DOUT[0].n3 DOUT[0].t0 26.5955
R20377 DOUT[0].n3 DOUT[0].t1 26.5955
R20378 DOUT[0].n0 DOUT[0].t3 24.9236
R20379 DOUT[0].n0 DOUT[0].t2 24.9236
R20380 DOUT[0] DOUT[0].n4 10.4965
R20381 DOUT[0].n2 DOUT[0] 10.4965
R20382 DOUT[0] DOUT[0].n5 9.66056
R20383 DOUT[0].n4 DOUT[0] 6.9125
R20384 DOUT[0].n2 DOUT[0] 6.9125
R20385 DOUT[0].n5 DOUT[0] 4.3525
R20386 DOUT[0].n1 DOUT[0] 1.7925
R20387 a_7999_4373.n3 a_7999_4373.n0 807.871
R20388 a_7999_4373.n4 a_7999_4373.t6 389.183
R20389 a_7999_4373.n5 a_7999_4373.n4 251.167
R20390 a_7999_4373.t0 a_7999_4373.n5 223.571
R20391 a_7999_4373.n1 a_7999_4373.t8 212.081
R20392 a_7999_4373.n2 a_7999_4373.t3 212.081
R20393 a_7999_4373.n3 a_7999_4373.n2 176.576
R20394 a_7999_4373.n4 a_7999_4373.t5 174.891
R20395 a_7999_4373.n1 a_7999_4373.t4 139.78
R20396 a_7999_4373.n2 a_7999_4373.t7 139.78
R20397 a_7999_4373.n0 a_7999_4373.t1 63.3219
R20398 a_7999_4373.n0 a_7999_4373.t2 63.3219
R20399 a_7999_4373.n2 a_7999_4373.n1 61.346
R20400 a_7999_4373.n5 a_7999_4373.n3 37.7195
R20401 a_9575_9117.n0 a_9575_9117.t1 1327.82
R20402 a_9575_9117.t0 a_9575_9117.n0 194.655
R20403 a_9575_9117.n0 a_9575_9117.t2 63.3219
R20404 a_10237_6005.n3 a_10237_6005.n2 647.119
R20405 a_10237_6005.n1 a_10237_6005.t5 350.253
R20406 a_10237_6005.n2 a_10237_6005.n0 260.339
R20407 a_10237_6005.n2 a_10237_6005.n1 246.119
R20408 a_10237_6005.n1 a_10237_6005.t4 189.588
R20409 a_10237_6005.n3 a_10237_6005.t1 89.1195
R20410 a_10237_6005.n0 a_10237_6005.t0 63.3338
R20411 a_10237_6005.t2 a_10237_6005.n3 41.0422
R20412 a_10237_6005.n0 a_10237_6005.t3 31.9797
R20413 a_10127_6031.t0 a_10127_6031.n0 1327.82
R20414 a_10127_6031.n0 a_10127_6031.t1 194.655
R20415 a_10127_6031.n0 a_10127_6031.t2 63.3219
R20416 a_7631_8511.n5 a_7631_8511.n4 807.871
R20417 a_7631_8511.n2 a_7631_8511.t8 389.183
R20418 a_7631_8511.n3 a_7631_8511.n2 251.167
R20419 a_7631_8511.n3 a_7631_8511.t1 223.571
R20420 a_7631_8511.n0 a_7631_8511.t4 212.081
R20421 a_7631_8511.n1 a_7631_8511.t6 212.081
R20422 a_7631_8511.n4 a_7631_8511.n1 176.576
R20423 a_7631_8511.n2 a_7631_8511.t3 174.891
R20424 a_7631_8511.n0 a_7631_8511.t7 139.78
R20425 a_7631_8511.n1 a_7631_8511.t5 139.78
R20426 a_7631_8511.t0 a_7631_8511.n5 63.3219
R20427 a_7631_8511.n5 a_7631_8511.t2 63.3219
R20428 a_7631_8511.n1 a_7631_8511.n0 61.346
R20429 a_7631_8511.n4 a_7631_8511.n3 37.7195
R20430 a_7565_8585.n0 a_7565_8585.t0 68.3338
R20431 a_7565_8585.n0 a_7565_8585.t1 26.3935
R20432 a_7565_8585.n1 a_7565_8585.n0 14.4005
R20433 a_7368_9019.t1 a_7368_9019.n3 370.026
R20434 a_7368_9019.n0 a_7368_9019.t3 351.356
R20435 a_7368_9019.n1 a_7368_9019.t5 334.717
R20436 a_7368_9019.n3 a_7368_9019.t0 325.971
R20437 a_7368_9019.n1 a_7368_9019.t4 309.935
R20438 a_7368_9019.n0 a_7368_9019.t2 305.683
R20439 a_7368_9019.n2 a_7368_9019.n0 16.879
R20440 a_7368_9019.n3 a_7368_9019.n2 10.8867
R20441 a_7368_9019.n2 a_7368_9019.n1 9.3005
R20442 a_7324_9117.t0 a_7324_9117.t1 126.644
R20443 a_4148_5059.t0 a_4148_5059.n3 370.026
R20444 a_4148_5059.n0 a_4148_5059.t4 351.356
R20445 a_4148_5059.n1 a_4148_5059.t3 334.717
R20446 a_4148_5059.n3 a_4148_5059.t1 325.971
R20447 a_4148_5059.n1 a_4148_5059.t2 309.935
R20448 a_4148_5059.n0 a_4148_5059.t5 305.683
R20449 a_4148_5059.n2 a_4148_5059.n0 16.879
R20450 a_4148_5059.n3 a_4148_5059.n2 10.8867
R20451 a_4148_5059.n2 a_4148_5059.n1 9.3005
R20452 a_4906_4943.n1 a_4906_4943.n0 926.024
R20453 a_4906_4943.n1 a_4906_4943.t3 82.0838
R20454 a_4906_4943.n0 a_4906_4943.t0 63.3338
R20455 a_4906_4943.t1 a_4906_4943.n1 63.3219
R20456 a_4906_4943.n0 a_4906_4943.t2 29.7268
R20457 a_1941_10927.t0 a_1941_10927.n3 370.026
R20458 a_1941_10927.n0 a_1941_10927.t2 351.356
R20459 a_1941_10927.n1 a_1941_10927.t4 334.717
R20460 a_1941_10927.n3 a_1941_10927.t1 325.971
R20461 a_1941_10927.n1 a_1941_10927.t5 309.935
R20462 a_1941_10927.n0 a_1941_10927.t3 305.683
R20463 a_1941_10927.n2 a_1941_10927.n0 16.879
R20464 a_1941_10927.n3 a_1941_10927.n2 10.8867
R20465 a_1941_10927.n2 a_1941_10927.n1 9.3005
R20466 a_2509_11169.n3 a_2509_11169.n2 647.119
R20467 a_2509_11169.n1 a_2509_11169.t4 350.253
R20468 a_2509_11169.n2 a_2509_11169.n0 260.339
R20469 a_2509_11169.n2 a_2509_11169.n1 246.119
R20470 a_2509_11169.n1 a_2509_11169.t5 189.588
R20471 a_2509_11169.n3 a_2509_11169.t2 89.1195
R20472 a_2509_11169.n0 a_2509_11169.t3 63.3338
R20473 a_2509_11169.t0 a_2509_11169.n3 41.0422
R20474 a_2509_11169.n0 a_2509_11169.t1 31.9797
R20475 a_2439_4541.n1 a_2439_4541.t5 530.01
R20476 a_2439_4541.t0 a_2439_4541.n5 421.021
R20477 a_2439_4541.n0 a_2439_4541.t3 337.171
R20478 a_2439_4541.n3 a_2439_4541.t1 280.223
R20479 a_2439_4541.n4 a_2439_4541.t6 263.173
R20480 a_2439_4541.n4 a_2439_4541.t2 227.826
R20481 a_2439_4541.n0 a_2439_4541.t7 199.762
R20482 a_2439_4541.n2 a_2439_4541.n1 170.81
R20483 a_2439_4541.n2 a_2439_4541.n0 167.321
R20484 a_2439_4541.n5 a_2439_4541.n4 152
R20485 a_2439_4541.n1 a_2439_4541.t4 141.923
R20486 a_2439_4541.n3 a_2439_4541.n2 10.8376
R20487 a_2439_4541.n5 a_2439_4541.n3 2.50485
R20488 a_2400_4667.t0 a_2400_4667.n3 370.026
R20489 a_2400_4667.n0 a_2400_4667.t3 351.356
R20490 a_2400_4667.n1 a_2400_4667.t5 334.717
R20491 a_2400_4667.n3 a_2400_4667.t1 325.971
R20492 a_2400_4667.n1 a_2400_4667.t4 309.935
R20493 a_2400_4667.n0 a_2400_4667.t2 305.683
R20494 a_2400_4667.n2 a_2400_4667.n0 16.879
R20495 a_2400_4667.n3 a_2400_4667.n2 10.8867
R20496 a_2400_4667.n2 a_2400_4667.n1 9.3005
R20497 a_7109_8181.n3 a_7109_8181.n2 647.119
R20498 a_7109_8181.n1 a_7109_8181.t4 350.253
R20499 a_7109_8181.n2 a_7109_8181.n0 260.339
R20500 a_7109_8181.n2 a_7109_8181.n1 246.119
R20501 a_7109_8181.n1 a_7109_8181.t5 189.588
R20502 a_7109_8181.n3 a_7109_8181.t2 89.1195
R20503 a_7109_8181.n0 a_7109_8181.t3 63.3338
R20504 a_7109_8181.t0 a_7109_8181.n3 41.0422
R20505 a_7109_8181.n0 a_7109_8181.t1 31.9797
R20506 a_6987_8585.t1 a_6987_8585.t0 198.571
R20507 a_7153_8573.t0 a_7153_8573.t1 60.0005
R20508 a_4550_4765.n3 a_4550_4765.n2 647.119
R20509 a_4550_4765.n1 a_4550_4765.t5 350.253
R20510 a_4550_4765.n2 a_4550_4765.n0 260.339
R20511 a_4550_4765.n2 a_4550_4765.n1 246.119
R20512 a_4550_4765.n1 a_4550_4765.t4 189.588
R20513 a_4550_4765.n3 a_4550_4765.t2 89.1195
R20514 a_4550_4765.n0 a_4550_4765.t3 63.3338
R20515 a_4550_4765.t0 a_4550_4765.n3 41.0422
R20516 a_4550_4765.n0 a_4550_4765.t1 31.9797
R20517 a_4764_4765.t0 a_4764_4765.n0 1327.82
R20518 a_4764_4765.n0 a_4764_4765.t1 194.655
R20519 a_4764_4765.n0 a_4764_4765.t2 63.3219
R20520 a_7348_5487.n1 a_7348_5487.n0 926.024
R20521 a_7348_5487.n1 a_7348_5487.t2 82.0838
R20522 a_7348_5487.n0 a_7348_5487.t3 63.3338
R20523 a_7348_5487.t0 a_7348_5487.n1 63.3219
R20524 a_7348_5487.n0 a_7348_5487.t1 29.7268
R20525 a_7948_7637.n21 a_7948_7637.n20 316.591
R20526 a_7948_7637.n20 a_7948_7637.n0 217.256
R20527 a_7948_7637.n2 a_7948_7637.t10 212.081
R20528 a_7948_7637.n17 a_7948_7637.t9 212.081
R20529 a_7948_7637.n15 a_7948_7637.t6 212.081
R20530 a_7948_7637.n8 a_7948_7637.t11 212.081
R20531 a_7948_7637.n9 a_7948_7637.t4 212.081
R20532 a_7948_7637.n6 a_7948_7637.t7 212.081
R20533 a_7948_7637.n5 a_7948_7637.t5 212.081
R20534 a_7948_7637.n4 a_7948_7637.t15 212.081
R20535 a_7948_7637.n11 a_7948_7637.n7 169.409
R20536 a_7948_7637.n2 a_7948_7637.t18 162.274
R20537 a_7948_7637.n17 a_7948_7637.t17 162.274
R20538 a_7948_7637.n15 a_7948_7637.t14 162.274
R20539 a_7948_7637.n8 a_7948_7637.t19 162.274
R20540 a_7948_7637.n9 a_7948_7637.t12 162.274
R20541 a_7948_7637.n6 a_7948_7637.t16 162.274
R20542 a_7948_7637.n5 a_7948_7637.t13 162.274
R20543 a_7948_7637.n4 a_7948_7637.t8 162.274
R20544 a_7948_7637.n11 a_7948_7637.n10 152
R20545 a_7948_7637.n12 a_7948_7637.n3 152
R20546 a_7948_7637.n14 a_7948_7637.n13 152
R20547 a_7948_7637.n16 a_7948_7637.n1 152
R20548 a_7948_7637.n19 a_7948_7637.n18 152
R20549 a_7948_7637.n6 a_7948_7637.n5 55.2698
R20550 a_7948_7637.n5 a_7948_7637.n4 55.2698
R20551 a_7948_7637.n14 a_7948_7637.n3 43.7018
R20552 a_7948_7637.n20 a_7948_7637.n19 43.5205
R20553 a_7948_7637.n0 a_7948_7637.t2 40.0005
R20554 a_7948_7637.n0 a_7948_7637.t3 40.0005
R20555 a_7948_7637.n16 a_7948_7637.n15 39.8458
R20556 a_7948_7637.n10 a_7948_7637.n8 35.9898
R20557 a_7948_7637.n7 a_7948_7637.n6 30.8485
R20558 a_7948_7637.n18 a_7948_7637.n17 28.2778
R20559 a_7948_7637.n21 a_7948_7637.t0 27.5805
R20560 a_7948_7637.t1 a_7948_7637.n21 27.5805
R20561 a_7948_7637.n18 a_7948_7637.n2 26.9925
R20562 a_7948_7637.n9 a_7948_7637.n7 24.4218
R20563 a_7948_7637.n10 a_7948_7637.n9 19.2805
R20564 a_7948_7637.n19 a_7948_7637.n1 17.4085
R20565 a_7948_7637.n13 a_7948_7637.n1 17.4085
R20566 a_7948_7637.n13 a_7948_7637.n12 17.4085
R20567 a_7948_7637.n12 a_7948_7637.n11 17.4085
R20568 a_7948_7637.n17 a_7948_7637.n16 15.4245
R20569 a_7948_7637.n8 a_7948_7637.n3 7.7125
R20570 a_7948_7637.n15 a_7948_7637.n14 3.8565
R20571 clkload0.X.n8 clkload0.X.n6 333.392
R20572 clkload0.X.n8 clkload0.X.n7 301.392
R20573 clkload0.X.n10 clkload0.X.n9 301.392
R20574 clkload0.X.n11 clkload0.X.n5 298.296
R20575 clkload0.X.n2 clkload0.X.n0 248.638
R20576 clkload0.X.n2 clkload0.X.n1 203.463
R20577 clkload0.X.n4 clkload0.X.n3 203.463
R20578 clkload0.X clkload0.X.n13 199.673
R20579 clkload0.X.n4 clkload0.X.n2 45.177
R20580 clkload0.X.n0 clkload0.X.t9 40.0005
R20581 clkload0.X.n0 clkload0.X.t10 40.0005
R20582 clkload0.X.n1 clkload0.X.t12 40.0005
R20583 clkload0.X.n1 clkload0.X.t8 40.0005
R20584 clkload0.X.n3 clkload0.X.t14 40.0005
R20585 clkload0.X.n3 clkload0.X.t11 40.0005
R20586 clkload0.X.n13 clkload0.X.t13 40.0005
R20587 clkload0.X.n13 clkload0.X.t15 40.0005
R20588 clkload0.X.n10 clkload0.X.n8 32.0005
R20589 clkload0.X.n6 clkload0.X.t2 27.5805
R20590 clkload0.X.n6 clkload0.X.t3 27.5805
R20591 clkload0.X.n7 clkload0.X.t5 27.5805
R20592 clkload0.X.n7 clkload0.X.t1 27.5805
R20593 clkload0.X.n5 clkload0.X.t6 27.5805
R20594 clkload0.X.n5 clkload0.X.t0 27.5805
R20595 clkload0.X.n9 clkload0.X.t7 27.5805
R20596 clkload0.X.n9 clkload0.X.t4 27.5805
R20597 clkload0.X.n12 clkload0.X.n4 27.1064
R20598 clkload0.X.n11 clkload0.X.n10 19.2005
R20599 clkload0.X.n12 clkload0.X 3.76132
R20600 clkload0.X clkload0.X.n11 2.2438
R20601 clkload0.X clkload0.X.n12 0.726273
R20602 a_5102_11471.n3 a_5102_11471.n2 647.119
R20603 a_5102_11471.n1 a_5102_11471.t4 350.253
R20604 a_5102_11471.n2 a_5102_11471.n0 260.339
R20605 a_5102_11471.n2 a_5102_11471.n1 246.119
R20606 a_5102_11471.n1 a_5102_11471.t5 189.588
R20607 a_5102_11471.n3 a_5102_11471.t1 89.1195
R20608 a_5102_11471.n0 a_5102_11471.t0 63.3338
R20609 a_5102_11471.t2 a_5102_11471.n3 41.0422
R20610 a_5102_11471.n0 a_5102_11471.t3 31.9797
R20611 a_5409_11837.t0 a_5409_11837.t1 60.0005
R20612 a_5481_11837.t1 a_5481_11837.t0 198.571
R20613 a_7827_3855.n0 a_7827_3855.t1 1327.82
R20614 a_7827_3855.t0 a_7827_3855.n0 194.655
R20615 a_7827_3855.n0 a_7827_3855.t2 63.3219
R20616 a_6927_3311.n1 a_6927_3311.t6 530.01
R20617 a_6927_3311.t0 a_6927_3311.n5 421.021
R20618 a_6927_3311.n0 a_6927_3311.t3 337.142
R20619 a_6927_3311.n3 a_6927_3311.t1 280.223
R20620 a_6927_3311.n4 a_6927_3311.t7 263.173
R20621 a_6927_3311.n4 a_6927_3311.t2 227.826
R20622 a_6927_3311.n0 a_6927_3311.t4 199.762
R20623 a_6927_3311.n2 a_6927_3311.n1 170.81
R20624 a_6927_3311.n2 a_6927_3311.n0 167.321
R20625 a_6927_3311.n5 a_6927_3311.n4 152
R20626 a_6927_3311.n1 a_6927_3311.t5 141.923
R20627 a_6927_3311.n3 a_6927_3311.n2 10.8376
R20628 a_6927_3311.n5 a_6927_3311.n3 2.50485
R20629 a_7093_3311.t0 a_7093_3311.n3 370.026
R20630 a_7093_3311.n0 a_7093_3311.t4 351.356
R20631 a_7093_3311.n1 a_7093_3311.t2 334.717
R20632 a_7093_3311.n3 a_7093_3311.t1 325.971
R20633 a_7093_3311.n1 a_7093_3311.t5 309.935
R20634 a_7093_3311.n0 a_7093_3311.t3 305.683
R20635 a_7093_3311.n2 a_7093_3311.n0 16.879
R20636 a_7093_3311.n3 a_7093_3311.n2 10.8867
R20637 a_7093_3311.n2 a_7093_3311.n1 9.3005
R20638 a_10111_3311.n3 a_10111_3311.n2 674.338
R20639 a_10111_3311.n1 a_10111_3311.t4 332.58
R20640 a_10111_3311.n2 a_10111_3311.n0 284.012
R20641 a_10111_3311.n2 a_10111_3311.n1 253.648
R20642 a_10111_3311.n1 a_10111_3311.t5 168.701
R20643 a_10111_3311.n3 a_10111_3311.t2 96.1553
R20644 a_10111_3311.t1 a_10111_3311.n3 65.6672
R20645 a_10111_3311.n0 a_10111_3311.t3 65.0005
R20646 a_10111_3311.n0 a_10111_3311.t0 45.0005
R20647 a_10207_3311.t1 a_10207_3311.t0 198.571
R20648 a_4765_8573.t0 a_4765_8573.t1 60.0005
R20649 a_4698_2899.n3 a_4698_2899.n2 636.953
R20650 a_4698_2899.n1 a_4698_2899.t5 366.856
R20651 a_4698_2899.n2 a_4698_2899.n0 300.2
R20652 a_4698_2899.n2 a_4698_2899.n1 225.036
R20653 a_4698_2899.n1 a_4698_2899.t4 174.056
R20654 a_4698_2899.n0 a_4698_2899.t2 70.0005
R20655 a_4698_2899.t0 a_4698_2899.n3 68.0124
R20656 a_4698_2899.n3 a_4698_2899.t3 63.3219
R20657 a_4698_2899.n0 a_4698_2899.t1 61.6672
R20658 a_4411_2741.n5 a_4411_2741.n4 807.871
R20659 a_4411_2741.n0 a_4411_2741.t5 389.183
R20660 a_4411_2741.n1 a_4411_2741.n0 251.167
R20661 a_4411_2741.n1 a_4411_2741.t1 223.571
R20662 a_4411_2741.n3 a_4411_2741.t3 212.081
R20663 a_4411_2741.n2 a_4411_2741.t7 212.081
R20664 a_4411_2741.n4 a_4411_2741.n3 176.576
R20665 a_4411_2741.n0 a_4411_2741.t6 174.891
R20666 a_4411_2741.n3 a_4411_2741.t8 139.78
R20667 a_4411_2741.n2 a_4411_2741.t4 139.78
R20668 a_4411_2741.t0 a_4411_2741.n5 63.3219
R20669 a_4411_2741.n5 a_4411_2741.t2 63.3219
R20670 a_4411_2741.n3 a_4411_2741.n2 61.346
R20671 a_4411_2741.n4 a_4411_2741.n1 37.5061
R20672 a_3859_4373.n3 a_3859_4373.n0 807.871
R20673 a_3859_4373.n4 a_3859_4373.t4 389.183
R20674 a_3859_4373.n5 a_3859_4373.n4 251.167
R20675 a_3859_4373.t0 a_3859_4373.n5 223.571
R20676 a_3859_4373.n2 a_3859_4373.t7 212.081
R20677 a_3859_4373.n1 a_3859_4373.t8 212.081
R20678 a_3859_4373.n3 a_3859_4373.n2 176.576
R20679 a_3859_4373.n4 a_3859_4373.t5 174.891
R20680 a_3859_4373.n2 a_3859_4373.t3 139.78
R20681 a_3859_4373.n1 a_3859_4373.t6 139.78
R20682 a_3859_4373.n0 a_3859_4373.t2 63.3219
R20683 a_3859_4373.n0 a_3859_4373.t1 63.3219
R20684 a_3859_4373.n2 a_3859_4373.n1 61.346
R20685 a_3859_4373.n5 a_3859_4373.n3 37.5061
R20686 SWP[6].n5 SWP[6].n4 585
R20687 SWP[6].n4 SWP[6].n3 585
R20688 SWP[6].n0 SWP[6].t4 333.651
R20689 SWP[6].n0 SWP[6].t5 297.233
R20690 SWP[6].n7 SWP[6].n0 195.701
R20691 SWP[6].n2 SWP[6].n1 185
R20692 SWP[6] SWP[6].n2 49.0339
R20693 SWP[6].n7 SWP[6].n6 42.1523
R20694 SWP[6].n4 SWP[6].t1 26.5955
R20695 SWP[6].n4 SWP[6].t0 26.5955
R20696 SWP[6].n1 SWP[6].t3 24.9236
R20697 SWP[6].n1 SWP[6].t2 24.9236
R20698 SWP[6].n6 SWP[6] 24.0538
R20699 SWP[6].n3 SWP[6] 15.6165
R20700 SWP[6].n6 SWP[6].n5 11.8605
R20701 SWP[6].n2 SWP[6] 10.4965
R20702 SWP[6].n5 SWP[6] 1.7925
R20703 SWP[6].n3 SWP[6] 1.7925
R20704 SWP[6] SWP[6].n7 1.03669
R20705 a_4181_8751.t0 a_4181_8751.t1 87.1434
R20706 a_9669_6037.t0 a_9669_6037.n3 370.026
R20707 a_9669_6037.n0 a_9669_6037.t2 351.356
R20708 a_9669_6037.n1 a_9669_6037.t3 334.717
R20709 a_9669_6037.n3 a_9669_6037.t1 325.971
R20710 a_9669_6037.n1 a_9669_6037.t4 309.935
R20711 a_9669_6037.n0 a_9669_6037.t5 305.683
R20712 a_9669_6037.n2 a_9669_6037.n0 16.879
R20713 a_9669_6037.n3 a_9669_6037.n2 10.8867
R20714 a_9669_6037.n2 a_9669_6037.n1 9.3005
R20715 a_10584_6409.n3 a_10584_6409.n2 636.953
R20716 a_10584_6409.n1 a_10584_6409.t4 366.856
R20717 a_10584_6409.n2 a_10584_6409.n0 300.2
R20718 a_10584_6409.n2 a_10584_6409.n1 225.036
R20719 a_10584_6409.n1 a_10584_6409.t5 174.056
R20720 a_10584_6409.n0 a_10584_6409.t1 70.0005
R20721 a_10584_6409.n3 a_10584_6409.t3 68.0124
R20722 a_10584_6409.t0 a_10584_6409.n3 63.3219
R20723 a_10584_6409.n0 a_10584_6409.t2 61.6672
R20724 DOUT[5].n2 DOUT[5].n1 585
R20725 DOUT[5].n1 DOUT[5].n0 585
R20726 DOUT[5].n4 DOUT[5].n3 185
R20727 DOUT[5].n4 DOUT[5] 57.7379
R20728 DOUT[5].n1 DOUT[5].t1 26.5955
R20729 DOUT[5].n1 DOUT[5].t0 26.5955
R20730 DOUT[5].n3 DOUT[5].t2 24.9236
R20731 DOUT[5].n3 DOUT[5].t3 24.9236
R20732 DOUT[5] DOUT[5].n2 10.4965
R20733 DOUT[5].n0 DOUT[5] 10.4965
R20734 DOUT[5].n2 DOUT[5] 6.9125
R20735 DOUT[5].n0 DOUT[5] 6.9125
R20736 DOUT[5] DOUT[5].n4 1.7925
R20737 a_6251_10901.n3 a_6251_10901.n0 807.871
R20738 a_6251_10901.n4 a_6251_10901.t6 389.183
R20739 a_6251_10901.n5 a_6251_10901.n4 251.167
R20740 a_6251_10901.t0 a_6251_10901.n5 223.571
R20741 a_6251_10901.n1 a_6251_10901.t3 212.081
R20742 a_6251_10901.n2 a_6251_10901.t5 212.081
R20743 a_6251_10901.n3 a_6251_10901.n2 176.576
R20744 a_6251_10901.n4 a_6251_10901.t4 174.891
R20745 a_6251_10901.n1 a_6251_10901.t7 139.78
R20746 a_6251_10901.n2 a_6251_10901.t8 139.78
R20747 a_6251_10901.n0 a_6251_10901.t1 63.3219
R20748 a_6251_10901.n0 a_6251_10901.t2 63.3219
R20749 a_6251_10901.n2 a_6251_10901.n1 61.346
R20750 a_6251_10901.n5 a_6251_10901.n3 37.7195
R20751 a_7164_4399.n1 a_7164_4399.n0 926.024
R20752 a_7164_4399.n1 a_7164_4399.t2 82.0838
R20753 a_7164_4399.n0 a_7164_4399.t3 63.3338
R20754 a_7164_4399.t0 a_7164_4399.n1 63.3219
R20755 a_7164_4399.n0 a_7164_4399.t1 29.7268
R20756 a_2439_5629.n1 a_2439_5629.t7 530.01
R20757 a_2439_5629.t1 a_2439_5629.n5 421.021
R20758 a_2439_5629.n0 a_2439_5629.t5 337.171
R20759 a_2439_5629.n3 a_2439_5629.t0 280.223
R20760 a_2439_5629.n4 a_2439_5629.t2 263.173
R20761 a_2439_5629.n4 a_2439_5629.t4 227.826
R20762 a_2439_5629.n0 a_2439_5629.t3 199.762
R20763 a_2439_5629.n2 a_2439_5629.n1 170.81
R20764 a_2439_5629.n2 a_2439_5629.n0 167.321
R20765 a_2439_5629.n5 a_2439_5629.n4 152
R20766 a_2439_5629.n1 a_2439_5629.t6 141.923
R20767 a_2439_5629.n3 a_2439_5629.n2 10.8376
R20768 a_2439_5629.n5 a_2439_5629.n3 2.50485
R20769 a_2400_5755.t0 a_2400_5755.n3 370.026
R20770 a_2400_5755.n0 a_2400_5755.t4 351.356
R20771 a_2400_5755.n1 a_2400_5755.t2 334.717
R20772 a_2400_5755.n3 a_2400_5755.t1 325.971
R20773 a_2400_5755.n1 a_2400_5755.t5 309.935
R20774 a_2400_5755.n0 a_2400_5755.t3 305.683
R20775 a_2400_5755.n2 a_2400_5755.n0 16.879
R20776 a_2400_5755.n3 a_2400_5755.n2 10.8867
R20777 a_2400_5755.n2 a_2400_5755.n1 9.3005
R20778 a_5659_3453.n1 a_5659_3453.t6 530.01
R20779 a_5659_3453.t0 a_5659_3453.n5 421.021
R20780 a_5659_3453.n0 a_5659_3453.t4 337.171
R20781 a_5659_3453.n3 a_5659_3453.t1 280.223
R20782 a_5659_3453.n4 a_5659_3453.t7 263.173
R20783 a_5659_3453.n4 a_5659_3453.t3 227.826
R20784 a_5659_3453.n0 a_5659_3453.t2 199.762
R20785 a_5659_3453.n2 a_5659_3453.n1 170.81
R20786 a_5659_3453.n2 a_5659_3453.n0 167.321
R20787 a_5659_3453.n5 a_5659_3453.n4 152
R20788 a_5659_3453.n1 a_5659_3453.t5 141.923
R20789 a_5659_3453.n3 a_5659_3453.n2 10.8376
R20790 a_5659_3453.n5 a_5659_3453.n3 2.50485
R20791 a_9563_7663.t1 a_9563_7663.t0 198.571
R20792 a_9729_7663.t0 a_9729_7663.t1 60.0005
R20793 x2/net13.n27 x2/net13.n26 244.069
R20794 x2/net13.n24 x2/net13.n0 236.589
R20795 x2/net13.n5 x2/net13.t18 212.081
R20796 x2/net13.n7 x2/net13.t10 212.081
R20797 x2/net13.n4 x2/net13.t15 212.081
R20798 x2/net13.n11 x2/net13.t20 212.081
R20799 x2/net13.n3 x2/net13.t12 212.081
R20800 x2/net13.n16 x2/net13.t22 212.081
R20801 x2/net13.n18 x2/net13.t16 212.081
R20802 x2/net13.n19 x2/net13.t19 212.081
R20803 x2/net13.n27 x2/net13.n25 204.893
R20804 x2/net13.n23 x2/net13.n1 188.492
R20805 x2/net13.n6 x2/net13 171.969
R20806 x2/net13.n21 x2/net13.n20 152
R20807 x2/net13.n17 x2/net13.n2 152
R20808 x2/net13.n15 x2/net13.n14 152
R20809 x2/net13.n13 x2/net13.n12 152
R20810 x2/net13.n10 x2/net13 152
R20811 x2/net13.n9 x2/net13.n8 152
R20812 x2/net13.n5 x2/net13.t8 139.78
R20813 x2/net13.n7 x2/net13.t14 139.78
R20814 x2/net13.n4 x2/net13.t21 139.78
R20815 x2/net13.n11 x2/net13.t11 139.78
R20816 x2/net13.n3 x2/net13.t17 139.78
R20817 x2/net13.n16 x2/net13.t13 139.78
R20818 x2/net13.n18 x2/net13.t23 139.78
R20819 x2/net13.n19 x2/net13.t9 139.78
R20820 x2/net13.n6 x2/net13.n5 30.6732
R20821 x2/net13.n7 x2/net13.n6 30.6732
R20822 x2/net13.n8 x2/net13.n7 30.6732
R20823 x2/net13.n8 x2/net13.n4 30.6732
R20824 x2/net13.n10 x2/net13.n4 30.6732
R20825 x2/net13.n11 x2/net13.n10 30.6732
R20826 x2/net13.n12 x2/net13.n11 30.6732
R20827 x2/net13.n12 x2/net13.n3 30.6732
R20828 x2/net13.n15 x2/net13.n3 30.6732
R20829 x2/net13.n16 x2/net13.n15 30.6732
R20830 x2/net13.n17 x2/net13.n16 30.6732
R20831 x2/net13.n18 x2/net13.n17 30.6732
R20832 x2/net13.n20 x2/net13.n18 30.6732
R20833 x2/net13.n20 x2/net13.n19 30.6732
R20834 x2/net13.n25 x2/net13.t1 26.5955
R20835 x2/net13.n25 x2/net13.t5 26.5955
R20836 x2/net13.n26 x2/net13.t7 26.5955
R20837 x2/net13.n26 x2/net13.t0 26.5955
R20838 x2/net13.n0 x2/net13.t6 24.9236
R20839 x2/net13.n0 x2/net13.t2 24.9236
R20840 x2/net13.n1 x2/net13.t4 24.9236
R20841 x2/net13.n1 x2/net13.t3 24.9236
R20842 x2/net13 x2/net13.n9 21.5045
R20843 x2/net13.n13 x2/net13 21.5045
R20844 x2/net13.n14 x2/net13 18.9445
R20845 x2/net13 x2/net13.n27 18.4569
R20846 x2/net13 x2/net13.n2 16.8965
R20847 x2/net13 x2/net13.n21 14.8485
R20848 x2/net13 x2/net13.n22 14.4935
R20849 x2/net13.n23 x2/net13 14.4935
R20850 x2/net13.n28 x2/net13 14.008
R20851 x2/net13.n28 x2/net13.n24 12.0894
R20852 x2/net13.n24 x2/net13.n23 11.8308
R20853 x2/net13.n21 x2/net13 8.7045
R20854 x2/net13.n14 x2/net13 4.6085
R20855 x2/net13.n22 x2/net13 4.3525
R20856 x2/net13 x2/net13.n13 2.5605
R20857 x2/net13 x2/net13.n28 2.41559
R20858 x2/net13.n22 x2/net13.n2 2.3045
R20859 x2/net13.n9 x2/net13 1.5365
R20860 a_4463_6717.n1 a_4463_6717.t4 530.01
R20861 a_4463_6717.t0 a_4463_6717.n5 421.021
R20862 a_4463_6717.n0 a_4463_6717.t2 337.171
R20863 a_4463_6717.n3 a_4463_6717.t1 280.223
R20864 a_4463_6717.n4 a_4463_6717.t6 263.173
R20865 a_4463_6717.n4 a_4463_6717.t7 227.826
R20866 a_4463_6717.n0 a_4463_6717.t5 199.762
R20867 a_4463_6717.n2 a_4463_6717.n1 170.81
R20868 a_4463_6717.n2 a_4463_6717.n0 167.321
R20869 a_4463_6717.n5 a_4463_6717.n4 152
R20870 a_4463_6717.n1 a_4463_6717.t3 141.923
R20871 a_4463_6717.n3 a_4463_6717.n2 10.8376
R20872 a_4463_6717.n5 a_4463_6717.n3 2.50485
R20873 a_4550_6941.n3 a_4550_6941.n2 647.119
R20874 a_4550_6941.n1 a_4550_6941.t5 350.253
R20875 a_4550_6941.n2 a_4550_6941.n0 260.339
R20876 a_4550_6941.n2 a_4550_6941.n1 246.119
R20877 a_4550_6941.n1 a_4550_6941.t4 189.588
R20878 a_4550_6941.n3 a_4550_6941.t3 89.1195
R20879 a_4550_6941.n0 a_4550_6941.t0 63.3338
R20880 a_4550_6941.t2 a_4550_6941.n3 41.0422
R20881 a_4550_6941.n0 a_4550_6941.t1 31.9797
R20882 a_9043_7125.n1 a_9043_7125.t4 530.01
R20883 a_9043_7125.t0 a_9043_7125.n5 421.021
R20884 a_9043_7125.n0 a_9043_7125.t7 337.142
R20885 a_9043_7125.n3 a_9043_7125.t1 280.223
R20886 a_9043_7125.n4 a_9043_7125.t3 263.173
R20887 a_9043_7125.n4 a_9043_7125.t6 227.826
R20888 a_9043_7125.n0 a_9043_7125.t2 199.762
R20889 a_9043_7125.n2 a_9043_7125.n1 170.81
R20890 a_9043_7125.n2 a_9043_7125.n0 167.321
R20891 a_9043_7125.n5 a_9043_7125.n4 152
R20892 a_9043_7125.n1 a_9043_7125.t5 141.923
R20893 a_9043_7125.n3 a_9043_7125.n2 10.8376
R20894 a_9043_7125.n5 a_9043_7125.n3 2.50485
R20895 a_10124_7497.n3 a_10124_7497.n2 636.953
R20896 a_10124_7497.n1 a_10124_7497.t4 366.856
R20897 a_10124_7497.n2 a_10124_7497.n0 300.2
R20898 a_10124_7497.n2 a_10124_7497.n1 225.036
R20899 a_10124_7497.n1 a_10124_7497.t5 174.056
R20900 a_10124_7497.n0 a_10124_7497.t0 70.0005
R20901 a_10124_7497.n3 a_10124_7497.t3 68.0124
R20902 a_10124_7497.t1 a_10124_7497.n3 63.3219
R20903 a_10124_7497.n0 a_10124_7497.t2 61.6672
R20904 a_10233_7497.n0 a_10233_7497.t1 68.3338
R20905 a_10233_7497.n0 a_10233_7497.t0 26.3935
R20906 a_10233_7497.n1 a_10233_7497.n0 14.4005
R20907 a_4330_7915.n3 a_4330_7915.n2 636.953
R20908 a_4330_7915.n1 a_4330_7915.t4 366.856
R20909 a_4330_7915.n2 a_4330_7915.n0 300.2
R20910 a_4330_7915.n2 a_4330_7915.n1 225.036
R20911 a_4330_7915.n1 a_4330_7915.t5 174.056
R20912 a_4330_7915.n0 a_4330_7915.t1 70.0005
R20913 a_4330_7915.t0 a_4330_7915.n3 68.0124
R20914 a_4330_7915.n3 a_4330_7915.t2 63.3219
R20915 a_4330_7915.n0 a_4330_7915.t3 61.6672
R20916 a_4365_7663.t0 a_4365_7663.t1 87.1434
R20917 a_10601_5321.n0 a_10601_5321.t0 68.3338
R20918 a_10601_5321.n0 a_10601_5321.t1 26.3935
R20919 a_10601_5321.n1 a_10601_5321.n0 14.4005
R20920 a_2019_6005.n5 a_2019_6005.n4 807.871
R20921 a_2019_6005.n0 a_2019_6005.t7 389.183
R20922 a_2019_6005.n1 a_2019_6005.n0 251.167
R20923 a_2019_6005.n1 a_2019_6005.t1 223.571
R20924 a_2019_6005.n3 a_2019_6005.t3 212.081
R20925 a_2019_6005.n2 a_2019_6005.t5 212.081
R20926 a_2019_6005.n4 a_2019_6005.n3 176.576
R20927 a_2019_6005.n0 a_2019_6005.t6 174.891
R20928 a_2019_6005.n3 a_2019_6005.t8 139.78
R20929 a_2019_6005.n2 a_2019_6005.t4 139.78
R20930 a_2019_6005.t0 a_2019_6005.n5 63.3219
R20931 a_2019_6005.n5 a_2019_6005.t2 63.3219
R20932 a_2019_6005.n3 a_2019_6005.n2 61.346
R20933 a_2019_6005.n4 a_2019_6005.n1 37.5061
R20934 a_2341_6397.t0 a_2341_6397.t1 87.1434
R20935 a_11030_3311.t0 a_11030_3311.t1 87.1434
R20936 a_7521_4399.t0 a_7521_4399.t1 60.0005
R20937 SWN[1].n2 SWN[1] 586.793
R20938 SWN[1].n3 SWN[1].n2 585
R20939 SWN[1].n1 SWN[1].n0 185
R20940 SWN[1] SWN[1].n1 49.0339
R20941 SWN[1].n2 SWN[1].t1 26.5955
R20942 SWN[1].n2 SWN[1].t0 26.5955
R20943 SWN[1].n0 SWN[1].t2 24.9236
R20944 SWN[1].n0 SWN[1].t3 24.9236
R20945 SWN[1].n3 SWN[1] 15.6165
R20946 SWN[1].n4 SWN[1] 13.0565
R20947 SWN[1].n1 SWN[1] 10.4965
R20948 SWN[1].n4 SWN[1] 9.66056
R20949 SWN[1] SWN[1].n4 4.3525
R20950 SWN[1] SWN[1].n3 1.7925
R20951 a_8178_4399.t0 a_8178_4399.t1 87.1434
R20952 a_10145_4917.n3 a_10145_4917.n2 647.119
R20953 a_10145_4917.n1 a_10145_4917.t4 350.253
R20954 a_10145_4917.n2 a_10145_4917.n0 260.339
R20955 a_10145_4917.n2 a_10145_4917.n1 246.119
R20956 a_10145_4917.n1 a_10145_4917.t5 189.588
R20957 a_10145_4917.n3 a_10145_4917.t0 89.1195
R20958 a_10145_4917.n0 a_10145_4917.t3 63.3338
R20959 a_10145_4917.t1 a_10145_4917.n3 41.0422
R20960 a_10145_4917.n0 a_10145_4917.t2 31.9797
R20961 a_10023_5321.t0 a_10023_5321.t1 198.571
R20962 a_10189_5309.t0 a_10189_5309.t1 60.0005
R20963 a_2905_5487.t1 a_2905_5487.t0 198.571
R20964 a_2595_5724.n3 a_2595_5724.n2 674.338
R20965 a_2595_5724.n1 a_2595_5724.t4 332.58
R20966 a_2595_5724.n2 a_2595_5724.n0 284.012
R20967 a_2595_5724.n2 a_2595_5724.n1 253.648
R20968 a_2595_5724.n1 a_2595_5724.t5 168.701
R20969 a_2595_5724.t0 a_2595_5724.n3 96.1553
R20970 a_2595_5724.n3 a_2595_5724.t3 65.6672
R20971 a_2595_5724.n0 a_2595_5724.t1 65.0005
R20972 a_2595_5724.n0 a_2595_5724.t2 45.0005
R20973 a_7185_6037.t0 a_7185_6037.n3 370.026
R20974 a_7185_6037.n0 a_7185_6037.t2 351.356
R20975 a_7185_6037.n1 a_7185_6037.t4 334.717
R20976 a_7185_6037.n3 a_7185_6037.t1 325.971
R20977 a_7185_6037.n1 a_7185_6037.t3 309.935
R20978 a_7185_6037.n0 a_7185_6037.t5 305.683
R20979 a_7185_6037.n2 a_7185_6037.n0 16.879
R20980 a_7185_6037.n3 a_7185_6037.n2 10.8867
R20981 a_7185_6037.n2 a_7185_6037.n1 9.3005
R20982 a_7753_6005.n3 a_7753_6005.n2 647.119
R20983 a_7753_6005.n1 a_7753_6005.t5 350.253
R20984 a_7753_6005.n2 a_7753_6005.n0 260.339
R20985 a_7753_6005.n2 a_7753_6005.n1 246.119
R20986 a_7753_6005.n1 a_7753_6005.t4 189.588
R20987 a_7753_6005.n3 a_7753_6005.t0 89.1195
R20988 a_7753_6005.n0 a_7753_6005.t1 63.3338
R20989 a_7753_6005.t2 a_7753_6005.n3 41.0422
R20990 a_7753_6005.n0 a_7753_6005.t3 31.9797
R20991 a_8100_6409.n3 a_8100_6409.n2 636.953
R20992 a_8100_6409.n1 a_8100_6409.t4 366.856
R20993 a_8100_6409.n2 a_8100_6409.n0 300.2
R20994 a_8100_6409.n2 a_8100_6409.n1 225.036
R20995 a_8100_6409.n1 a_8100_6409.t5 174.056
R20996 a_8100_6409.n0 a_8100_6409.t3 70.0005
R20997 a_8100_6409.t1 a_8100_6409.n3 68.0124
R20998 a_8100_6409.n3 a_8100_6409.t2 63.3219
R20999 a_8100_6409.n0 a_8100_6409.t0 61.6672
R21000 a_7156_6941.n0 a_7156_6941.t1 1327.82
R21001 a_7156_6941.n0 a_7156_6941.t2 194.655
R21002 a_7156_6941.t0 a_7156_6941.n0 63.3219
R21003 x2/TRIG1.n0 x2/TRIG1.t5 332.312
R21004 x2/TRIG1.n0 x2/TRIG1.t4 295.627
R21005 x2/TRIG1.n6 x2/TRIG1.n5 289.096
R21006 x2/TRIG1.n1 x2/TRIG1.n0 194.845
R21007 x2/TRIG1.n4 x2/TRIG1.n3 185
R21008 x2/TRIG1 x2/TRIG1.n4 49.0339
R21009 x2/TRIG1 x2/TRIG1.n1 31.4548
R21010 x2/TRIG1.n5 x2/TRIG1.t1 26.5955
R21011 x2/TRIG1.n5 x2/TRIG1.t0 26.5955
R21012 x2/TRIG1.n3 x2/TRIG1.t2 24.9236
R21013 x2/TRIG1.n3 x2/TRIG1.t3 24.9236
R21014 x2/TRIG1.n2 x2/TRIG1 15.4573
R21015 x2/TRIG1 x2/TRIG1.n6 9.48653
R21016 x2/TRIG1.n6 x2/TRIG1 7.7181
R21017 x2/TRIG1.n4 x2/TRIG1.n2 6.1445
R21018 x2/TRIG1.n2 x2/TRIG1 4.3525
R21019 x2/TRIG1.n1 x2/TRIG1 4.17441
R21020 a_9669_3861.t0 a_9669_3861.n3 370.026
R21021 a_9669_3861.n0 a_9669_3861.t3 351.356
R21022 a_9669_3861.n1 a_9669_3861.t4 334.717
R21023 a_9669_3861.n3 a_9669_3861.t1 325.971
R21024 a_9669_3861.n1 a_9669_3861.t5 309.935
R21025 a_9669_3861.n0 a_9669_3861.t2 305.683
R21026 a_9669_3861.n2 a_9669_3861.n0 16.879
R21027 a_9669_3861.n3 a_9669_3861.n2 10.8867
R21028 a_9669_3861.n2 a_9669_3861.n1 9.3005
R21029 a_10584_4233.n3 a_10584_4233.n2 636.953
R21030 a_10584_4233.n1 a_10584_4233.t5 366.856
R21031 a_10584_4233.n2 a_10584_4233.n0 300.2
R21032 a_10584_4233.n2 a_10584_4233.n1 225.036
R21033 a_10584_4233.n1 a_10584_4233.t4 174.056
R21034 a_10584_4233.n0 a_10584_4233.t2 70.0005
R21035 a_10584_4233.t0 a_10584_4233.n3 68.0124
R21036 a_10584_4233.n3 a_10584_4233.t3 63.3219
R21037 a_10584_4233.n0 a_10584_4233.t1 61.6672
R21038 a_10746_3855.t0 a_10746_3855.t1 126.644
R21039 a_7494_9117.n3 a_7494_9117.n2 647.119
R21040 a_7494_9117.n1 a_7494_9117.t4 350.253
R21041 a_7494_9117.n2 a_7494_9117.n0 260.339
R21042 a_7494_9117.n2 a_7494_9117.n1 246.119
R21043 a_7494_9117.n1 a_7494_9117.t5 189.588
R21044 a_7494_9117.n3 a_7494_9117.t0 89.1195
R21045 a_7494_9117.n0 a_7494_9117.t3 63.3338
R21046 a_7494_9117.t2 a_7494_9117.n3 41.0422
R21047 a_7494_9117.n0 a_7494_9117.t1 31.9797
R21048 a_7801_8751.t0 a_7801_8751.t1 60.0005
R21049 a_7873_8751.t1 a_7873_8751.t0 198.571
R21050 SWP[7].n0 SWP[7].t4 332.312
R21051 SWP[7].n0 SWP[7].t5 295.627
R21052 SWP[7].n2 SWP[7].n1 289.096
R21053 SWP[7] SWP[7].n0 196.004
R21054 SWP[7].n4 SWP[7].n3 185
R21055 SWP[7].n4 SWP[7] 49.0339
R21056 SWP[7].n6 SWP[7] 33.172
R21057 SWP[7].n1 SWP[7].t1 26.5955
R21058 SWP[7].n1 SWP[7].t0 26.5955
R21059 SWP[7].n3 SWP[7].t2 24.9236
R21060 SWP[7].n3 SWP[7].t3 24.9236
R21061 SWP[7] SWP[7].n6 21.5406
R21062 SWP[7] SWP[7].n5 11.0981
R21063 SWP[7] SWP[7].n2 9.48653
R21064 SWP[7].n2 SWP[7] 7.7181
R21065 SWP[7].n6 SWP[7] 6.61805
R21066 SWP[7].n5 SWP[7].n4 6.1445
R21067 SWP[7].n5 SWP[7] 4.3525
R21068 a_7365_8751.n0 a_7365_8751.t1 68.3338
R21069 a_7365_8751.n0 a_7365_8751.t0 26.3935
R21070 a_7365_8751.n1 a_7365_8751.n0 14.4005
R21071 a_8615_7457.n2 a_8615_7457.n1 672.948
R21072 a_8615_7457.n1 a_8615_7457.t1 314.563
R21073 a_8615_7457.n0 a_8615_7457.t3 236.18
R21074 a_8615_7457.n0 a_8615_7457.t4 163.881
R21075 a_8615_7457.n1 a_8615_7457.n0 152
R21076 a_8615_7457.t0 a_8615_7457.n2 63.3219
R21077 a_8615_7457.n2 a_8615_7457.t2 63.3219
R21078 a_7551_5853.t0 a_7551_5853.n0 1327.82
R21079 a_7551_5853.n0 a_7551_5853.t1 194.655
R21080 a_7551_5853.n0 a_7551_5853.t2 63.3219
R21081 a_7624_4221.n1 a_7624_4221.n0 926.024
R21082 a_7624_4221.n1 a_7624_4221.t2 82.0838
R21083 a_7624_4221.n0 a_7624_4221.t3 63.3338
R21084 a_7624_4221.t0 a_7624_4221.n1 63.3219
R21085 a_7624_4221.n0 a_7624_4221.t1 29.7268
R21086 a_2397_5487.n0 a_2397_5487.t1 68.3338
R21087 a_2397_5487.n0 a_2397_5487.t0 26.3935
R21088 a_2397_5487.n1 a_2397_5487.n0 14.4005
R21089 a_2122_5739.n3 a_2122_5739.n2 636.953
R21090 a_2122_5739.n1 a_2122_5739.t5 366.856
R21091 a_2122_5739.n2 a_2122_5739.n0 300.2
R21092 a_2122_5739.n2 a_2122_5739.n1 225.036
R21093 a_2122_5739.n1 a_2122_5739.t4 174.056
R21094 a_2122_5739.n0 a_2122_5739.t3 70.0005
R21095 a_2122_5739.t1 a_2122_5739.n3 68.0124
R21096 a_2122_5739.n3 a_2122_5739.t2 63.3219
R21097 a_2122_5739.n0 a_2122_5739.t0 61.6672
R21098 a_7019_6037.n1 a_7019_6037.t3 530.01
R21099 a_7019_6037.t0 a_7019_6037.n5 421.021
R21100 a_7019_6037.n0 a_7019_6037.t5 337.142
R21101 a_7019_6037.n3 a_7019_6037.t1 280.223
R21102 a_7019_6037.n4 a_7019_6037.t6 263.173
R21103 a_7019_6037.n4 a_7019_6037.t2 227.826
R21104 a_7019_6037.n0 a_7019_6037.t4 199.762
R21105 a_7019_6037.n2 a_7019_6037.n1 170.81
R21106 a_7019_6037.n2 a_7019_6037.n0 167.321
R21107 a_7019_6037.n5 a_7019_6037.n4 152
R21108 a_7019_6037.n1 a_7019_6037.t7 141.923
R21109 a_7019_6037.n3 a_7019_6037.n2 10.8376
R21110 a_7019_6037.n5 a_7019_6037.n3 2.50485
R21111 SWP[4].n3 SWP[4].n2 585
R21112 SWP[4].n2 SWP[4].n1 585
R21113 SWP[4].n0 SWP[4].t4 333.651
R21114 SWP[4].n0 SWP[4].t5 297.233
R21115 SWP[4].n7 SWP[4].n0 195.701
R21116 SWP[4].n5 SWP[4].n4 185
R21117 SWP[4].n7 SWP[4].n6 69.2636
R21118 SWP[4].n5 SWP[4] 57.7379
R21119 SWP[4].n2 SWP[4].t1 26.5955
R21120 SWP[4].n2 SWP[4].t0 26.5955
R21121 SWP[4].n4 SWP[4].t2 24.9236
R21122 SWP[4].n4 SWP[4].t3 24.9236
R21123 SWP[4].n6 SWP[4] 13.6525
R21124 SWP[4].n6 SWP[4] 11.0319
R21125 SWP[4] SWP[4].n3 10.4965
R21126 SWP[4].n1 SWP[4] 10.4965
R21127 SWP[4].n3 SWP[4] 6.9125
R21128 SWP[4].n1 SWP[4] 6.9125
R21129 SWP[4] SWP[4].n5 1.7925
R21130 SWP[4] SWP[4].n7 1.03669
R21131 a_9372_7663.n1 a_9372_7663.n0 926.024
R21132 a_9372_7663.t0 a_9372_7663.n1 82.0838
R21133 a_9372_7663.n0 a_9372_7663.t1 63.3338
R21134 a_9372_7663.n1 a_9372_7663.t2 63.3219
R21135 a_9372_7663.n0 a_9372_7663.t3 29.7268
R21136 a_5182_6941.n1 a_5182_6941.n0 926.024
R21137 a_5182_6941.t0 a_5182_6941.n1 82.0838
R21138 a_5182_6941.n0 a_5182_6941.t3 63.3338
R21139 a_5182_6941.n1 a_5182_6941.t1 63.3219
R21140 a_5182_6941.n0 a_5182_6941.t2 29.7268
R21141 a_2585_11477.t0 a_2585_11477.n3 370.026
R21142 a_2585_11477.n0 a_2585_11477.t3 351.356
R21143 a_2585_11477.n1 a_2585_11477.t2 334.717
R21144 a_2585_11477.n3 a_2585_11477.t1 325.971
R21145 a_2585_11477.n1 a_2585_11477.t4 309.935
R21146 a_2585_11477.n0 a_2585_11477.t5 305.683
R21147 a_2585_11477.n2 a_2585_11477.n0 16.879
R21148 a_2585_11477.n3 a_2585_11477.n2 10.8867
R21149 a_2585_11477.n2 a_2585_11477.n1 9.3005
R21150 a_2935_11849.n3 a_2935_11849.n2 674.338
R21151 a_2935_11849.n1 a_2935_11849.t4 332.58
R21152 a_2935_11849.n2 a_2935_11849.n0 284.012
R21153 a_2935_11849.n2 a_2935_11849.n1 253.648
R21154 a_2935_11849.n1 a_2935_11849.t5 168.701
R21155 a_2935_11849.t1 a_2935_11849.n3 96.1553
R21156 a_2935_11849.n3 a_2935_11849.t3 65.6672
R21157 a_2935_11849.n0 a_2935_11849.t0 65.0005
R21158 a_2935_11849.n0 a_2935_11849.t2 45.0005
R21159 a_3031_11849.t0 a_3031_11849.t1 198.571
R21160 DOUT[8].n4 DOUT[8].n3 585
R21161 DOUT[8].n3 DOUT[8].n2 585
R21162 DOUT[8].n1 DOUT[8].n0 185
R21163 DOUT[8].n2 DOUT[8] 49.758
R21164 DOUT[8] DOUT[8].n1 49.0339
R21165 DOUT[8].n3 DOUT[8].t1 26.5955
R21166 DOUT[8].n3 DOUT[8].t0 26.5955
R21167 DOUT[8].n0 DOUT[8].t3 24.9236
R21168 DOUT[8].n0 DOUT[8].t2 24.9236
R21169 DOUT[8].n4 DOUT[8] 15.6165
R21170 DOUT[8].n1 DOUT[8] 10.4965
R21171 DOUT[8].n2 DOUT[8] 1.7925
R21172 DOUT[8] DOUT[8].n4 1.7925
R21173 a_8701_7457.t0 a_8701_7457.t1 77.1434
R21174 a_5511_10927.n3 a_5511_10927.n2 674.338
R21175 a_5511_10927.n1 a_5511_10927.t5 332.58
R21176 a_5511_10927.n2 a_5511_10927.n0 284.012
R21177 a_5511_10927.n2 a_5511_10927.n1 253.648
R21178 a_5511_10927.n1 a_5511_10927.t4 168.701
R21179 a_5511_10927.n3 a_5511_10927.t2 96.1553
R21180 a_5511_10927.t0 a_5511_10927.n3 65.6672
R21181 a_5511_10927.n0 a_5511_10927.t3 65.0005
R21182 a_5511_10927.n0 a_5511_10927.t1 45.0005
R21183 a_5729_11169.n3 a_5729_11169.n2 647.119
R21184 a_5729_11169.n1 a_5729_11169.t4 350.253
R21185 a_5729_11169.n2 a_5729_11169.n0 260.339
R21186 a_5729_11169.n2 a_5729_11169.n1 246.119
R21187 a_5729_11169.n1 a_5729_11169.t5 189.588
R21188 a_5729_11169.n3 a_5729_11169.t1 89.1195
R21189 a_5729_11169.n0 a_5729_11169.t0 63.3338
R21190 a_5729_11169.t2 a_5729_11169.n3 41.0422
R21191 a_5729_11169.n0 a_5729_11169.t3 31.9797
R21192 a_4680_4221.n1 a_4680_4221.n0 926.024
R21193 a_4680_4221.n1 a_4680_4221.t3 82.0838
R21194 a_4680_4221.n0 a_4680_4221.t2 63.3338
R21195 a_4680_4221.t0 a_4680_4221.n1 63.3219
R21196 a_4680_4221.n0 a_4680_4221.t1 29.7268
R21197 a_4775_4233.n3 a_4775_4233.n2 674.338
R21198 a_4775_4233.n1 a_4775_4233.t5 332.58
R21199 a_4775_4233.n2 a_4775_4233.n0 284.012
R21200 a_4775_4233.n2 a_4775_4233.n1 253.648
R21201 a_4775_4233.n1 a_4775_4233.t4 168.701
R21202 a_4775_4233.t1 a_4775_4233.n3 96.1553
R21203 a_4775_4233.n3 a_4775_4233.t2 65.6672
R21204 a_4775_4233.n0 a_4775_4233.t0 65.0005
R21205 a_4775_4233.n0 a_4775_4233.t3 45.0005
R21206 a_10759_4159.n5 a_10759_4159.n4 807.871
R21207 a_10759_4159.n2 a_10759_4159.t6 389.183
R21208 a_10759_4159.n3 a_10759_4159.n2 251.167
R21209 a_10759_4159.n3 a_10759_4159.t1 223.571
R21210 a_10759_4159.n0 a_10759_4159.t3 212.081
R21211 a_10759_4159.n1 a_10759_4159.t4 212.081
R21212 a_10759_4159.n4 a_10759_4159.n1 176.576
R21213 a_10759_4159.n2 a_10759_4159.t5 174.891
R21214 a_10759_4159.n0 a_10759_4159.t7 139.78
R21215 a_10759_4159.n1 a_10759_4159.t8 139.78
R21216 a_10759_4159.n5 a_10759_4159.t2 63.3219
R21217 a_10759_4159.t0 a_10759_4159.n5 63.3219
R21218 a_10759_4159.n1 a_10759_4159.n0 61.346
R21219 a_10759_4159.n4 a_10759_4159.n3 37.7195
R21220 CF[5].n4 CF[5].n3 585
R21221 CF[5].n5 CF[5].n4 585
R21222 CF[5].n8 CF[5].t4 333.651
R21223 CF[5].n8 CF[5].t8 297.233
R21224 CF[5].n11 CF[5].t5 294.557
R21225 CF[5].n0 CF[5].t6 294.557
R21226 CF[5].n11 CF[5].t7 211.01
R21227 CF[5].n0 CF[5].t9 211.01
R21228 CF[5].n9 CF[5].n8 195.701
R21229 CF[5].n2 CF[5].n1 185
R21230 CF[5] CF[5].n11 156.207
R21231 CF[5] CF[5].n0 156.207
R21232 CF[5] CF[5].n2 57.7379
R21233 CF[5].n14 CF[5].n13 37.5972
R21234 CF[5].n13 CF[5].n10 29.6861
R21235 CF[5].n4 CF[5].t1 26.5955
R21236 CF[5].n4 CF[5].t0 26.5955
R21237 CF[5].n1 CF[5].t3 24.9236
R21238 CF[5].n1 CF[5].t2 24.9236
R21239 CF[5].n7 CF[5].n6 15.1865
R21240 CF[5] CF[5].n12 12.1248
R21241 CF[5].n10 CF[5].n7 10.5446
R21242 CF[5].n3 CF[5] 10.4965
R21243 CF[5].n5 CF[5] 10.4965
R21244 CF[5].n12 CF[5] 9.32621
R21245 CF[5].n14 CF[5] 9.32621
R21246 CF[5].n10 CF[5].n9 9.3005
R21247 CF[5].n3 CF[5] 6.9125
R21248 CF[5].n7 CF[5] 4.43761
R21249 CF[5].n6 CF[5] 4.3525
R21250 CF[5].n12 CF[5] 3.10907
R21251 CF[5] CF[5].n14 3.10907
R21252 CF[5].n13 CF[5] 2.80957
R21253 CF[5].n6 CF[5].n5 2.5605
R21254 CF[5].n2 CF[5] 1.7925
R21255 CF[5].n9 CF[5] 1.03669
R21256 a_4380_4765.t0 a_4380_4765.t1 126.644
R21257 a_5342_3563.n3 a_5342_3563.n2 636.953
R21258 a_5342_3563.n1 a_5342_3563.t4 366.856
R21259 a_5342_3563.n2 a_5342_3563.n0 300.2
R21260 a_5342_3563.n2 a_5342_3563.n1 225.036
R21261 a_5342_3563.n1 a_5342_3563.t5 174.056
R21262 a_5342_3563.n0 a_5342_3563.t3 70.0005
R21263 a_5342_3563.t1 a_5342_3563.n3 68.0124
R21264 a_5342_3563.n3 a_5342_3563.t2 63.3219
R21265 a_5342_3563.n0 a_5342_3563.t0 61.6672
R21266 a_5377_3311.t0 a_5377_3311.t1 87.1434
R21267 a_2419_11477.n1 a_2419_11477.t5 530.01
R21268 a_2419_11477.t0 a_2419_11477.n5 421.021
R21269 a_2419_11477.n0 a_2419_11477.t4 337.142
R21270 a_2419_11477.n3 a_2419_11477.t1 280.223
R21271 a_2419_11477.n4 a_2419_11477.t6 263.173
R21272 a_2419_11477.n4 a_2419_11477.t7 227.826
R21273 a_2419_11477.n0 a_2419_11477.t3 199.762
R21274 a_2419_11477.n2 a_2419_11477.n1 170.81
R21275 a_2419_11477.n2 a_2419_11477.n0 167.321
R21276 a_2419_11477.n5 a_2419_11477.n4 152
R21277 a_2419_11477.n1 a_2419_11477.t2 141.923
R21278 a_2419_11477.n3 a_2419_11477.n2 10.8376
R21279 a_2419_11477.n5 a_2419_11477.n3 2.50485
R21280 x2/net4.n0 x2/net4.t5 333.651
R21281 x2/net4.n0 x2/net4.t4 297.233
R21282 x2/net4.n6 x2/net4.n5 289.096
R21283 x2/net4.n1 x2/net4.n0 193.506
R21284 x2/net4.n4 x2/net4.n3 185
R21285 x2/net4 x2/net4.n4 49.0339
R21286 x2/net4 x2/net4.n1 26.979
R21287 x2/net4.n5 x2/net4.t0 26.5955
R21288 x2/net4.n5 x2/net4.t1 26.5955
R21289 x2/net4.n3 x2/net4.t2 24.9236
R21290 x2/net4.n3 x2/net4.t3 24.9236
R21291 x2/net4.n2 x2/net4 20.2272
R21292 x2/net4 x2/net4.n6 9.48653
R21293 x2/net4.n6 x2/net4 7.7181
R21294 x2/net4.n4 x2/net4.n2 6.1445
R21295 x2/net4.n2 x2/net4 4.3525
R21296 x2/net4.n1 x2/net4 4.17441
R21297 a_9287_10687.n4 a_9287_10687.n1 807.871
R21298 a_9287_10687.n0 a_9287_10687.t4 389.183
R21299 a_9287_10687.n5 a_9287_10687.n0 251.167
R21300 a_9287_10687.t0 a_9287_10687.n5 223.571
R21301 a_9287_10687.n2 a_9287_10687.t7 212.081
R21302 a_9287_10687.n3 a_9287_10687.t6 212.081
R21303 a_9287_10687.n4 a_9287_10687.n3 176.576
R21304 a_9287_10687.n0 a_9287_10687.t5 174.891
R21305 a_9287_10687.n2 a_9287_10687.t3 139.78
R21306 a_9287_10687.n3 a_9287_10687.t8 139.78
R21307 a_9287_10687.n1 a_9287_10687.t1 63.3219
R21308 a_9287_10687.n1 a_9287_10687.t2 63.3219
R21309 a_9287_10687.n3 a_9287_10687.n2 61.346
R21310 a_9287_10687.n5 a_9287_10687.n4 37.7195
R21311 a_9411_9839.n1 a_9411_9839.t5 530.01
R21312 a_9411_9839.t0 a_9411_9839.n5 421.021
R21313 a_9411_9839.n0 a_9411_9839.t4 337.142
R21314 a_9411_9839.n3 a_9411_9839.t1 280.223
R21315 a_9411_9839.n4 a_9411_9839.t2 263.173
R21316 a_9411_9839.n4 a_9411_9839.t6 227.826
R21317 a_9411_9839.n0 a_9411_9839.t7 199.762
R21318 a_9411_9839.n2 a_9411_9839.n1 170.81
R21319 a_9411_9839.n2 a_9411_9839.n0 167.321
R21320 a_9411_9839.n5 a_9411_9839.n4 152
R21321 a_9411_9839.n1 a_9411_9839.t3 141.923
R21322 a_9411_9839.n3 a_9411_9839.n2 10.8376
R21323 a_9411_9839.n5 a_9411_9839.n3 2.50485
R21324 a_9577_9839.t0 a_9577_9839.n3 370.026
R21325 a_9577_9839.n0 a_9577_9839.t4 351.356
R21326 a_9577_9839.n1 a_9577_9839.t2 334.717
R21327 a_9577_9839.n3 a_9577_9839.t1 325.971
R21328 a_9577_9839.n1 a_9577_9839.t3 309.935
R21329 a_9577_9839.n0 a_9577_9839.t5 305.683
R21330 a_9577_9839.n2 a_9577_9839.n0 16.879
R21331 a_9577_9839.n3 a_9577_9839.n2 10.8867
R21332 a_9577_9839.n2 a_9577_9839.n1 9.3005
R21333 a_7011_6812.n3 a_7011_6812.n2 674.338
R21334 a_7011_6812.n1 a_7011_6812.t4 332.58
R21335 a_7011_6812.n2 a_7011_6812.n0 284.012
R21336 a_7011_6812.n2 a_7011_6812.n1 253.648
R21337 a_7011_6812.n1 a_7011_6812.t5 168.701
R21338 a_7011_6812.n3 a_7011_6812.t3 96.1553
R21339 a_7011_6812.t0 a_7011_6812.n3 65.6672
R21340 a_7011_6812.n0 a_7011_6812.t2 65.0005
R21341 a_7011_6812.n0 a_7011_6812.t1 45.0005
R21342 a_2659_10761.n3 a_2659_10761.n2 674.338
R21343 a_2659_10761.n1 a_2659_10761.t4 332.58
R21344 a_2659_10761.n2 a_2659_10761.n0 284.012
R21345 a_2659_10761.n2 a_2659_10761.n1 253.648
R21346 a_2659_10761.n1 a_2659_10761.t5 168.701
R21347 a_2659_10761.t1 a_2659_10761.n3 96.1553
R21348 a_2659_10761.n3 a_2659_10761.t3 65.6672
R21349 a_2659_10761.n0 a_2659_10761.t0 65.0005
R21350 a_2659_10761.n0 a_2659_10761.t2 45.0005
R21351 a_8183_5461.n5 a_8183_5461.n4 807.871
R21352 a_8183_5461.n2 a_8183_5461.t3 389.183
R21353 a_8183_5461.n3 a_8183_5461.n2 251.167
R21354 a_8183_5461.n3 a_8183_5461.t2 223.571
R21355 a_8183_5461.n0 a_8183_5461.t4 212.081
R21356 a_8183_5461.n1 a_8183_5461.t8 212.081
R21357 a_8183_5461.n4 a_8183_5461.n1 176.576
R21358 a_8183_5461.n2 a_8183_5461.t6 174.891
R21359 a_8183_5461.n0 a_8183_5461.t7 139.78
R21360 a_8183_5461.n1 a_8183_5461.t5 139.78
R21361 a_8183_5461.n5 a_8183_5461.t1 63.3219
R21362 a_8183_5461.t0 a_8183_5461.n5 63.3219
R21363 a_8183_5461.n1 a_8183_5461.n0 61.346
R21364 a_8183_5461.n4 a_8183_5461.n3 37.7195
R21365 a_2291_10927.n3 a_2291_10927.n2 674.338
R21366 a_2291_10927.n1 a_2291_10927.t4 332.58
R21367 a_2291_10927.n2 a_2291_10927.n0 284.012
R21368 a_2291_10927.n2 a_2291_10927.n1 253.648
R21369 a_2291_10927.n1 a_2291_10927.t5 168.701
R21370 a_2291_10927.t1 a_2291_10927.n3 96.1553
R21371 a_2291_10927.n3 a_2291_10927.t2 65.6672
R21372 a_2291_10927.n0 a_2291_10927.t0 65.0005
R21373 a_2291_10927.n0 a_2291_10927.t3 45.0005
R21374 a_2399_11293.n0 a_2399_11293.t2 1327.82
R21375 a_2399_11293.t0 a_2399_11293.n0 194.655
R21376 a_2399_11293.n0 a_2399_11293.t1 63.3219
R21377 a_10759_3071.n4 a_10759_3071.n1 807.871
R21378 a_10759_3071.n0 a_10759_3071.t4 389.183
R21379 a_10759_3071.n5 a_10759_3071.n0 251.167
R21380 a_10759_3071.t0 a_10759_3071.n5 223.571
R21381 a_10759_3071.n2 a_10759_3071.t7 212.081
R21382 a_10759_3071.n3 a_10759_3071.t8 212.081
R21383 a_10759_3071.n4 a_10759_3071.n3 176.576
R21384 a_10759_3071.n0 a_10759_3071.t3 174.891
R21385 a_10759_3071.n2 a_10759_3071.t5 139.78
R21386 a_10759_3071.n3 a_10759_3071.t6 139.78
R21387 a_10759_3071.n1 a_10759_3071.t1 63.3219
R21388 a_10759_3071.n1 a_10759_3071.t2 63.3219
R21389 a_10759_3071.n3 a_10759_3071.n2 61.346
R21390 a_10759_3071.n5 a_10759_3071.n4 37.7195
R21391 a_2071_8893.n1 a_2071_8893.t7 530.01
R21392 a_2071_8893.t0 a_2071_8893.n5 421.021
R21393 a_2071_8893.n0 a_2071_8893.t3 337.171
R21394 a_2071_8893.n3 a_2071_8893.t1 280.223
R21395 a_2071_8893.n4 a_2071_8893.t2 263.173
R21396 a_2071_8893.n4 a_2071_8893.t5 227.826
R21397 a_2071_8893.n0 a_2071_8893.t4 199.762
R21398 a_2071_8893.n2 a_2071_8893.n1 170.81
R21399 a_2071_8893.n2 a_2071_8893.n0 167.321
R21400 a_2071_8893.n5 a_2071_8893.n4 152
R21401 a_2071_8893.n1 a_2071_8893.t6 141.923
R21402 a_2071_8893.n3 a_2071_8893.n2 10.8376
R21403 a_2071_8893.n5 a_2071_8893.n3 2.50485
R21404 a_4826_10383.n3 a_4826_10383.n2 647.119
R21405 a_4826_10383.n1 a_4826_10383.t4 350.253
R21406 a_4826_10383.n2 a_4826_10383.n0 260.339
R21407 a_4826_10383.n2 a_4826_10383.n1 246.119
R21408 a_4826_10383.n1 a_4826_10383.t5 189.588
R21409 a_4826_10383.n3 a_4826_10383.t0 89.1195
R21410 a_4826_10383.n0 a_4826_10383.t1 63.3338
R21411 a_4826_10383.t2 a_4826_10383.n3 41.0422
R21412 a_4826_10383.n0 a_4826_10383.t3 31.9797
R21413 a_9761_5487.t0 a_9761_5487.n3 370.026
R21414 a_9761_5487.n0 a_9761_5487.t3 351.356
R21415 a_9761_5487.n1 a_9761_5487.t4 334.717
R21416 a_9761_5487.n3 a_9761_5487.t1 325.971
R21417 a_9761_5487.n1 a_9761_5487.t2 309.935
R21418 a_9761_5487.n0 a_9761_5487.t5 305.683
R21419 a_9761_5487.n2 a_9761_5487.n0 16.879
R21420 a_9761_5487.n3 a_9761_5487.n2 10.8867
R21421 a_9761_5487.n2 a_9761_5487.n1 9.3005
R21422 a_3891_12015.n1 a_3891_12015.t7 530.01
R21423 a_3891_12015.t0 a_3891_12015.n5 421.021
R21424 a_3891_12015.n0 a_3891_12015.t2 337.142
R21425 a_3891_12015.n3 a_3891_12015.t1 280.223
R21426 a_3891_12015.n4 a_3891_12015.t4 263.173
R21427 a_3891_12015.n4 a_3891_12015.t5 227.826
R21428 a_3891_12015.n0 a_3891_12015.t6 199.762
R21429 a_3891_12015.n2 a_3891_12015.n1 170.81
R21430 a_3891_12015.n2 a_3891_12015.n0 167.321
R21431 a_3891_12015.n5 a_3891_12015.n4 152
R21432 a_3891_12015.n1 a_3891_12015.t3 141.923
R21433 a_3891_12015.n3 a_3891_12015.n2 10.8376
R21434 a_3891_12015.n5 a_3891_12015.n3 2.50485
R21435 a_6076_10927.n3 a_6076_10927.n2 636.953
R21436 a_6076_10927.n1 a_6076_10927.t4 366.856
R21437 a_6076_10927.n2 a_6076_10927.n0 300.2
R21438 a_6076_10927.n2 a_6076_10927.n1 225.036
R21439 a_6076_10927.n1 a_6076_10927.t5 174.056
R21440 a_6076_10927.n0 a_6076_10927.t1 70.0005
R21441 a_6076_10927.n3 a_6076_10927.t3 68.0124
R21442 a_6076_10927.t0 a_6076_10927.n3 63.3219
R21443 a_6076_10927.n0 a_6076_10927.t2 61.6672
R21444 a_6430_10927.t0 a_6430_10927.t1 87.1434
R21445 a_5383_5629.n1 a_5383_5629.t4 530.01
R21446 a_5383_5629.t0 a_5383_5629.n5 421.021
R21447 a_5383_5629.n0 a_5383_5629.t3 337.171
R21448 a_5383_5629.n3 a_5383_5629.t1 280.223
R21449 a_5383_5629.n4 a_5383_5629.t7 263.173
R21450 a_5383_5629.n4 a_5383_5629.t2 227.826
R21451 a_5383_5629.n0 a_5383_5629.t5 199.762
R21452 a_5383_5629.n2 a_5383_5629.n1 170.81
R21453 a_5383_5629.n2 a_5383_5629.n0 167.321
R21454 a_5383_5629.n5 a_5383_5629.n4 152
R21455 a_5383_5629.n1 a_5383_5629.t6 141.923
R21456 a_5383_5629.n3 a_5383_5629.n2 10.8376
R21457 a_5383_5629.n5 a_5383_5629.n3 2.50485
R21458 a_5344_5755.t0 a_5344_5755.n3 370.026
R21459 a_5344_5755.n0 a_5344_5755.t3 351.356
R21460 a_5344_5755.n1 a_5344_5755.t4 334.717
R21461 a_5344_5755.n3 a_5344_5755.t1 325.971
R21462 a_5344_5755.n1 a_5344_5755.t5 309.935
R21463 a_5344_5755.n0 a_5344_5755.t2 305.683
R21464 a_5344_5755.n2 a_5344_5755.n0 16.879
R21465 a_5344_5755.n3 a_5344_5755.n2 10.8867
R21466 a_5344_5755.n2 a_5344_5755.n1 9.3005
R21467 a_10851_5461.n5 a_10851_5461.n4 807.871
R21468 a_10851_5461.n2 a_10851_5461.t7 389.183
R21469 a_10851_5461.n3 a_10851_5461.n2 251.167
R21470 a_10851_5461.n3 a_10851_5461.t1 223.571
R21471 a_10851_5461.n0 a_10851_5461.t4 212.081
R21472 a_10851_5461.n1 a_10851_5461.t5 212.081
R21473 a_10851_5461.n4 a_10851_5461.n1 176.576
R21474 a_10851_5461.n2 a_10851_5461.t8 174.891
R21475 a_10851_5461.n0 a_10851_5461.t6 139.78
R21476 a_10851_5461.n1 a_10851_5461.t3 139.78
R21477 a_10851_5461.n5 a_10851_5461.t2 63.3219
R21478 a_10851_5461.t0 a_10851_5461.n5 63.3219
R21479 a_10851_5461.n1 a_10851_5461.n0 61.346
R21480 a_10851_5461.n4 a_10851_5461.n3 37.7195
R21481 CF[7].n0 CF[7] 586.793
R21482 CF[7].n1 CF[7].n0 585
R21483 CF[7].n11 CF[7].t9 333.651
R21484 CF[7].n11 CF[7].t7 297.233
R21485 CF[7].n5 CF[7].t6 294.557
R21486 CF[7].n8 CF[7].t4 294.557
R21487 CF[7].n5 CF[7].t8 211.01
R21488 CF[7].n8 CF[7].t5 211.01
R21489 CF[7].n12 CF[7].n11 195.701
R21490 CF[7].n3 CF[7].n2 185
R21491 CF[7].n6 CF[7].n5 152
R21492 CF[7].n9 CF[7].n8 152
R21493 CF[7].n3 CF[7] 49.0339
R21494 CF[7].n13 CF[7].n10 40.8439
R21495 CF[7].n0 CF[7].t1 26.5955
R21496 CF[7].n0 CF[7].t0 26.5955
R21497 CF[7].n2 CF[7].t2 24.9236
R21498 CF[7].n2 CF[7].t3 24.9236
R21499 CF[7].n10 CF[7] 20.107
R21500 CF[7].n1 CF[7] 15.6165
R21501 CF[7].n10 CF[7].n7 15.4806
R21502 CF[7] CF[7].n4 15.3283
R21503 CF[7].n14 CF[7].n13 11.7615
R21504 CF[7] CF[7].n9 10.4234
R21505 CF[7].n7 CF[7] 9.32621
R21506 CF[7].n13 CF[7].n12 9.3005
R21507 CF[7].n4 CF[7].n3 6.1445
R21508 CF[7] CF[7].n14 5.27626
R21509 CF[7].n4 CF[7] 4.3525
R21510 CF[7].n6 CF[7] 2.01193
R21511 CF[7].n9 CF[7] 2.01193
R21512 CF[7] CF[7].n1 1.7925
R21513 CF[7].n7 CF[7].n6 1.09764
R21514 CF[7].n12 CF[7] 1.03669
R21515 CF[7].n14 CF[7] 0.162245
R21516 a_4764_6941.t0 a_4764_6941.n0 1327.82
R21517 a_4764_6941.n0 a_4764_6941.t1 194.655
R21518 a_4764_6941.n0 a_4764_6941.t2 63.3219
R21519 a_4332_8323.t0 a_4332_8323.n3 370.026
R21520 a_4332_8323.n0 a_4332_8323.t2 351.356
R21521 a_4332_8323.n1 a_4332_8323.t3 334.717
R21522 a_4332_8323.n3 a_4332_8323.t1 325.971
R21523 a_4332_8323.n1 a_4332_8323.t4 309.935
R21524 a_4332_8323.n0 a_4332_8323.t5 305.683
R21525 a_4332_8323.n2 a_4332_8323.n0 16.879
R21526 a_4332_8323.n3 a_4332_8323.n2 10.8867
R21527 a_4332_8323.n2 a_4332_8323.n1 9.3005
R21528 a_4054_8339.n3 a_4054_8339.n2 636.953
R21529 a_4054_8339.n1 a_4054_8339.t4 366.856
R21530 a_4054_8339.n2 a_4054_8339.n0 300.2
R21531 a_4054_8339.n2 a_4054_8339.n1 225.036
R21532 a_4054_8339.n1 a_4054_8339.t5 174.056
R21533 a_4054_8339.n0 a_4054_8339.t2 70.0005
R21534 a_4054_8339.t0 a_4054_8339.n3 68.0124
R21535 a_4054_8339.n3 a_4054_8339.t3 63.3219
R21536 a_4054_8339.n0 a_4054_8339.t1 61.6672
R21537 a_4458_8207.n3 a_4458_8207.n2 647.119
R21538 a_4458_8207.n1 a_4458_8207.t4 350.253
R21539 a_4458_8207.n2 a_4458_8207.n0 260.339
R21540 a_4458_8207.n2 a_4458_8207.n1 246.119
R21541 a_4458_8207.n1 a_4458_8207.t5 189.588
R21542 a_4458_8207.n3 a_4458_8207.t2 89.1195
R21543 a_4458_8207.n0 a_4458_8207.t3 63.3338
R21544 a_4458_8207.t0 a_4458_8207.n3 41.0422
R21545 a_4458_8207.n0 a_4458_8207.t1 31.9797
R21546 a_7551_11293.n0 a_7551_11293.t1 1327.82
R21547 a_7551_11293.n0 a_7551_11293.t2 194.655
R21548 a_7551_11293.t0 a_7551_11293.n0 63.3219
R21549 a_2439_7805.n1 a_2439_7805.t2 530.01
R21550 a_2439_7805.t0 a_2439_7805.n5 421.021
R21551 a_2439_7805.n0 a_2439_7805.t6 337.171
R21552 a_2439_7805.n3 a_2439_7805.t1 280.223
R21553 a_2439_7805.n4 a_2439_7805.t4 263.173
R21554 a_2439_7805.n4 a_2439_7805.t7 227.826
R21555 a_2439_7805.n0 a_2439_7805.t5 199.762
R21556 a_2439_7805.n2 a_2439_7805.n1 170.81
R21557 a_2439_7805.n2 a_2439_7805.n0 167.321
R21558 a_2439_7805.n5 a_2439_7805.n4 152
R21559 a_2439_7805.n1 a_2439_7805.t3 141.923
R21560 a_2439_7805.n3 a_2439_7805.n2 10.8376
R21561 a_2439_7805.n5 a_2439_7805.n3 2.50485
R21562 a_2740_8029.n0 a_2740_8029.t2 1327.82
R21563 a_2740_8029.n0 a_2740_8029.t1 194.655
R21564 a_2740_8029.t0 a_2740_8029.n0 63.3219
R21565 a_2595_7900.n3 a_2595_7900.n2 674.338
R21566 a_2595_7900.n1 a_2595_7900.t4 332.58
R21567 a_2595_7900.n2 a_2595_7900.n0 284.012
R21568 a_2595_7900.n2 a_2595_7900.n1 253.648
R21569 a_2595_7900.n1 a_2595_7900.t5 168.701
R21570 a_2595_7900.n3 a_2595_7900.t1 96.1553
R21571 a_2595_7900.t0 a_2595_7900.n3 65.6672
R21572 a_2595_7900.n0 a_2595_7900.t2 65.0005
R21573 a_2595_7900.n0 a_2595_7900.t3 45.0005
R21574 a_2526_10205.n3 a_2526_10205.n2 647.119
R21575 a_2526_10205.n1 a_2526_10205.t4 350.253
R21576 a_2526_10205.n2 a_2526_10205.n0 260.339
R21577 a_2526_10205.n2 a_2526_10205.n1 246.119
R21578 a_2526_10205.n1 a_2526_10205.t5 189.588
R21579 a_2526_10205.n3 a_2526_10205.t3 89.1195
R21580 a_2526_10205.n0 a_2526_10205.t0 63.3338
R21581 a_2526_10205.t1 a_2526_10205.n3 41.0422
R21582 a_2526_10205.n0 a_2526_10205.t2 31.9797
R21583 a_2833_9839.t0 a_2833_9839.t1 60.0005
R21584 a_2905_9839.t1 a_2905_9839.t0 198.571
R21585 a_7171_7637.n3 a_7171_7637.n0 807.871
R21586 a_7171_7637.n4 a_7171_7637.t6 389.183
R21587 a_7171_7637.n5 a_7171_7637.n4 251.167
R21588 a_7171_7637.t0 a_7171_7637.n5 223.571
R21589 a_7171_7637.n1 a_7171_7637.t8 212.081
R21590 a_7171_7637.n2 a_7171_7637.t4 212.081
R21591 a_7171_7637.n3 a_7171_7637.n2 176.576
R21592 a_7171_7637.n4 a_7171_7637.t3 174.891
R21593 a_7171_7637.n1 a_7171_7637.t5 139.78
R21594 a_7171_7637.n2 a_7171_7637.t7 139.78
R21595 a_7171_7637.n0 a_7171_7637.t1 63.3219
R21596 a_7171_7637.n0 a_7171_7637.t2 63.3219
R21597 a_7171_7637.n2 a_7171_7637.n1 61.346
R21598 a_7171_7637.n5 a_7171_7637.n3 37.7195
R21599 a_7105_7663.t1 a_7105_7663.t0 94.7268
R21600 a_2397_9839.n0 a_2397_9839.t1 68.3338
R21601 a_2397_9839.n0 a_2397_9839.t0 26.3935
R21602 a_2397_9839.n1 a_2397_9839.n0 14.4005
R21603 a_1973_5309.t0 a_1973_5309.t1 87.1434
R21604 a_4733_3133.t0 a_4733_3133.t1 87.1434
R21605 DOUT[6].n3 DOUT[6].n2 585
R21606 DOUT[6].n4 DOUT[6].n3 585
R21607 DOUT[6].n1 DOUT[6].n0 185
R21608 DOUT[6] DOUT[6].n4 58.7606
R21609 DOUT[6] DOUT[6].n1 49.0339
R21610 DOUT[6].n3 DOUT[6].t0 26.5955
R21611 DOUT[6].n3 DOUT[6].t1 26.5955
R21612 DOUT[6].n0 DOUT[6].t3 24.9236
R21613 DOUT[6].n0 DOUT[6].t2 24.9236
R21614 DOUT[6].n2 DOUT[6] 15.6165
R21615 DOUT[6].n1 DOUT[6] 10.4965
R21616 DOUT[6].n4 DOUT[6] 1.7925
R21617 DOUT[6].n2 DOUT[6] 1.7925
R21618 a_4608_7931.t0 a_4608_7931.n3 370.026
R21619 a_4608_7931.n0 a_4608_7931.t4 351.356
R21620 a_4608_7931.n1 a_4608_7931.t5 334.717
R21621 a_4608_7931.n3 a_4608_7931.t1 325.971
R21622 a_4608_7931.n1 a_4608_7931.t3 309.935
R21623 a_4608_7931.n0 a_4608_7931.t2 305.683
R21624 a_4608_7931.n2 a_4608_7931.n0 16.879
R21625 a_4608_7931.n3 a_4608_7931.n2 10.8867
R21626 a_4608_7931.n2 a_4608_7931.n1 9.3005
R21627 a_4564_8029.t0 a_4564_8029.t1 126.644
R21628 a_4424_9019.t0 a_4424_9019.n3 370.026
R21629 a_4424_9019.n0 a_4424_9019.t4 351.356
R21630 a_4424_9019.n1 a_4424_9019.t2 334.717
R21631 a_4424_9019.n3 a_4424_9019.t1 325.971
R21632 a_4424_9019.n1 a_4424_9019.t5 309.935
R21633 a_4424_9019.n0 a_4424_9019.t3 305.683
R21634 a_4424_9019.n2 a_4424_9019.n0 16.879
R21635 a_4424_9019.n3 a_4424_9019.n2 10.8867
R21636 a_4424_9019.n2 a_4424_9019.n1 9.3005
R21637 a_3675_11775.n4 a_3675_11775.n1 807.871
R21638 a_3675_11775.n0 a_3675_11775.t4 389.183
R21639 a_3675_11775.n5 a_3675_11775.n0 251.167
R21640 a_3675_11775.t0 a_3675_11775.n5 223.571
R21641 a_3675_11775.n2 a_3675_11775.t7 212.081
R21642 a_3675_11775.n3 a_3675_11775.t6 212.081
R21643 a_3675_11775.n4 a_3675_11775.n3 176.576
R21644 a_3675_11775.n0 a_3675_11775.t5 174.891
R21645 a_3675_11775.n2 a_3675_11775.t3 139.78
R21646 a_3675_11775.n3 a_3675_11775.t8 139.78
R21647 a_3675_11775.n1 a_3675_11775.t1 63.3219
R21648 a_3675_11775.n1 a_3675_11775.t2 63.3219
R21649 a_3675_11775.n3 a_3675_11775.n2 61.346
R21650 a_3675_11775.n5 a_3675_11775.n4 37.7195
R21651 x2/net10.n4 x2/net10.n3 585
R21652 x2/net10.n5 x2/net10.n4 585
R21653 x2/net10.n0 x2/net10.t5 333.651
R21654 x2/net10.n0 x2/net10.t4 297.233
R21655 x2/net10 x2/net10.n0 194.062
R21656 x2/net10.n2 x2/net10.n1 185
R21657 x2/net10 x2/net10.n2 57.7379
R21658 x2/net10.n4 x2/net10.t0 26.5955
R21659 x2/net10.n4 x2/net10.t1 26.5955
R21660 x2/net10.n1 x2/net10.t3 24.9236
R21661 x2/net10.n1 x2/net10.t2 24.9236
R21662 x2/net10.n3 x2/net10 10.4965
R21663 x2/net10.n5 x2/net10 10.4965
R21664 x2/net10.n3 x2/net10 6.9125
R21665 x2/net10 x2/net10.n5 6.9125
R21666 x2/net10.n2 x2/net10 1.7925
R21667 a_2465_8573.t0 a_2465_8573.t1 60.0005
R21668 a_2537_8573.t0 a_2537_8573.t1 198.571
R21669 DOUT[3].n4 DOUT[3].n3 585
R21670 DOUT[3].n3 DOUT[3].n2 585
R21671 DOUT[3].n1 DOUT[3].n0 185
R21672 DOUT[3].n5 DOUT[3].n1 53.3859
R21673 DOUT[3] DOUT[3].n5 43.7315
R21674 DOUT[3].n3 DOUT[3].t1 26.5955
R21675 DOUT[3].n3 DOUT[3].t0 26.5955
R21676 DOUT[3].n0 DOUT[3].t2 24.9236
R21677 DOUT[3].n0 DOUT[3].t3 24.9236
R21678 DOUT[3] DOUT[3].n4 10.4965
R21679 DOUT[3].n2 DOUT[3] 10.4965
R21680 DOUT[3].n4 DOUT[3] 6.9125
R21681 DOUT[3].n2 DOUT[3] 6.9125
R21682 DOUT[3].n5 DOUT[3] 4.3525
R21683 DOUT[3].n1 DOUT[3] 1.7925
R21684 a_8425_6603.t0 a_8425_6603.t1 77.1434
R21685 a_2400_7931.t0 a_2400_7931.n3 370.026
R21686 a_2400_7931.n0 a_2400_7931.t3 351.356
R21687 a_2400_7931.n1 a_2400_7931.t4 334.717
R21688 a_2400_7931.n3 a_2400_7931.t1 325.971
R21689 a_2400_7931.n1 a_2400_7931.t2 309.935
R21690 a_2400_7931.n0 a_2400_7931.t5 305.683
R21691 a_2400_7931.n2 a_2400_7931.n0 16.879
R21692 a_2400_7931.n3 a_2400_7931.n2 10.8867
R21693 a_2400_7931.n2 a_2400_7931.n1 9.3005
R21694 a_3158_8029.n1 a_3158_8029.n0 926.024
R21695 a_3158_8029.t1 a_3158_8029.n1 82.0838
R21696 a_3158_8029.n0 a_3158_8029.t0 63.3338
R21697 a_3158_8029.n1 a_3158_8029.t3 63.3219
R21698 a_3158_8029.n0 a_3158_8029.t2 29.7268
R21699 a_7708_2767.n0 a_7708_2767.t1 1327.82
R21700 a_7708_2767.n0 a_7708_2767.t2 194.655
R21701 a_7708_2767.t0 a_7708_2767.n0 63.3219
R21702 a_10194_8029.t0 a_10194_8029.t1 126.644
R21703 a_4647_7805.n1 a_4647_7805.t6 530.01
R21704 a_4647_7805.t0 a_4647_7805.n5 421.021
R21705 a_4647_7805.n0 a_4647_7805.t3 337.171
R21706 a_4647_7805.n3 a_4647_7805.t1 280.223
R21707 a_4647_7805.n4 a_4647_7805.t2 263.173
R21708 a_4647_7805.n4 a_4647_7805.t5 227.826
R21709 a_4647_7805.n0 a_4647_7805.t4 199.762
R21710 a_4647_7805.n2 a_4647_7805.n1 170.81
R21711 a_4647_7805.n2 a_4647_7805.n0 167.321
R21712 a_4647_7805.n5 a_4647_7805.n4 152
R21713 a_4647_7805.n1 a_4647_7805.t7 141.923
R21714 a_4647_7805.n3 a_4647_7805.n2 10.8376
R21715 a_4647_7805.n5 a_4647_7805.n3 2.50485
R21716 a_4929_8751.t1 a_4929_8751.t0 198.571
R21717 a_4619_8988.n3 a_4619_8988.n2 674.338
R21718 a_4619_8988.n1 a_4619_8988.t4 332.58
R21719 a_4619_8988.n2 a_4619_8988.n0 284.012
R21720 a_4619_8988.n2 a_4619_8988.n1 253.648
R21721 a_4619_8988.n1 a_4619_8988.t5 168.701
R21722 a_4619_8988.n3 a_4619_8988.t2 96.1553
R21723 a_4619_8988.t1 a_4619_8988.n3 65.6672
R21724 a_4619_8988.n0 a_4619_8988.t3 65.0005
R21725 a_4619_8988.n0 a_4619_8988.t0 45.0005
R21726 a_5171_2741.n3 a_5171_2741.n2 674.338
R21727 a_5171_2741.n1 a_5171_2741.t4 332.58
R21728 a_5171_2741.n2 a_5171_2741.n0 284.012
R21729 a_5171_2741.n2 a_5171_2741.n1 253.648
R21730 a_5171_2741.n1 a_5171_2741.t5 168.701
R21731 a_5171_2741.t1 a_5171_2741.n3 96.1553
R21732 a_5171_2741.n3 a_5171_2741.t2 65.6672
R21733 a_5171_2741.n0 a_5171_2741.t0 65.0005
R21734 a_5171_2741.n0 a_5171_2741.t3 45.0005
R21735 a_10851_3285.n5 a_10851_3285.n4 807.871
R21736 a_10851_3285.n2 a_10851_3285.t3 389.183
R21737 a_10851_3285.n3 a_10851_3285.n2 251.167
R21738 a_10851_3285.n3 a_10851_3285.t1 223.571
R21739 a_10851_3285.n0 a_10851_3285.t8 212.081
R21740 a_10851_3285.n1 a_10851_3285.t5 212.081
R21741 a_10851_3285.n4 a_10851_3285.n1 176.576
R21742 a_10851_3285.n2 a_10851_3285.t6 174.891
R21743 a_10851_3285.n0 a_10851_3285.t4 139.78
R21744 a_10851_3285.n1 a_10851_3285.t7 139.78
R21745 a_10851_3285.n5 a_10851_3285.t2 63.3219
R21746 a_10851_3285.t0 a_10851_3285.n5 63.3219
R21747 a_10851_3285.n1 a_10851_3285.n0 61.346
R21748 a_10851_3285.n4 a_10851_3285.n3 37.7195
R21749 a_6927_5487.n1 a_6927_5487.t3 530.01
R21750 a_6927_5487.t0 a_6927_5487.n5 421.021
R21751 a_6927_5487.n0 a_6927_5487.t6 337.142
R21752 a_6927_5487.n3 a_6927_5487.t1 280.223
R21753 a_6927_5487.n4 a_6927_5487.t4 263.173
R21754 a_6927_5487.n4 a_6927_5487.t5 227.826
R21755 a_6927_5487.n0 a_6927_5487.t7 199.762
R21756 a_6927_5487.n2 a_6927_5487.n1 170.81
R21757 a_6927_5487.n2 a_6927_5487.n0 167.321
R21758 a_6927_5487.n5 a_6927_5487.n4 152
R21759 a_6927_5487.n1 a_6927_5487.t2 141.923
R21760 a_6927_5487.n3 a_6927_5487.n2 10.8376
R21761 a_6927_5487.n5 a_6927_5487.n3 2.50485
R21762 a_7443_5487.n3 a_7443_5487.n2 674.338
R21763 a_7443_5487.n1 a_7443_5487.t4 332.58
R21764 a_7443_5487.n2 a_7443_5487.n0 284.012
R21765 a_7443_5487.n2 a_7443_5487.n1 253.648
R21766 a_7443_5487.n1 a_7443_5487.t5 168.701
R21767 a_7443_5487.n3 a_7443_5487.t2 96.1553
R21768 a_7443_5487.t0 a_7443_5487.n3 65.6672
R21769 a_7443_5487.n0 a_7443_5487.t3 65.0005
R21770 a_7443_5487.n0 a_7443_5487.t1 45.0005
R21771 a_8170_5853.t0 a_8170_5853.t1 126.644
R21772 a_10019_6409.n3 a_10019_6409.n2 674.338
R21773 a_10019_6409.n1 a_10019_6409.t5 332.58
R21774 a_10019_6409.n2 a_10019_6409.n0 284.012
R21775 a_10019_6409.n2 a_10019_6409.n1 253.648
R21776 a_10019_6409.n1 a_10019_6409.t4 168.701
R21777 a_10019_6409.n3 a_10019_6409.t2 96.1553
R21778 a_10019_6409.t0 a_10019_6409.n3 65.6672
R21779 a_10019_6409.n0 a_10019_6409.t3 65.0005
R21780 a_10019_6409.n0 a_10019_6409.t1 45.0005
R21781 a_10115_6409.t1 a_10115_6409.t0 198.571
R21782 SWN[0].n4 SWN[0].n3 585
R21783 SWN[0].n3 SWN[0].n2 585
R21784 SWN[0].n1 SWN[0].n0 185
R21785 SWN[0] SWN[0].n1 49.0339
R21786 SWN[0].n3 SWN[0].t0 26.5955
R21787 SWN[0].n3 SWN[0].t1 26.5955
R21788 SWN[0].n0 SWN[0].t3 24.9236
R21789 SWN[0].n0 SWN[0].t2 24.9236
R21790 SWN[0].n2 SWN[0] 23.3526
R21791 SWN[0].n4 SWN[0] 15.6165
R21792 SWN[0].n1 SWN[0] 10.4965
R21793 SWN[0].n2 SWN[0] 1.7925
R21794 SWN[0] SWN[0].n4 1.7925
R21795 a_1835_7637.n3 a_1835_7637.n0 807.871
R21796 a_1835_7637.n4 a_1835_7637.t4 389.183
R21797 a_1835_7637.n5 a_1835_7637.n4 251.167
R21798 a_1835_7637.t0 a_1835_7637.n5 223.571
R21799 a_1835_7637.n2 a_1835_7637.t8 212.081
R21800 a_1835_7637.n1 a_1835_7637.t6 212.081
R21801 a_1835_7637.n3 a_1835_7637.n2 176.576
R21802 a_1835_7637.n4 a_1835_7637.t7 174.891
R21803 a_1835_7637.n2 a_1835_7637.t5 139.78
R21804 a_1835_7637.n1 a_1835_7637.t3 139.78
R21805 a_1835_7637.n0 a_1835_7637.t2 63.3219
R21806 a_1835_7637.n0 a_1835_7637.t1 63.3219
R21807 a_1835_7637.n2 a_1835_7637.n1 61.346
R21808 a_1835_7637.n5 a_1835_7637.n3 37.5061
R21809 DOUT[9].n4 DOUT[9].n3 585
R21810 DOUT[9].n3 DOUT[9].n2 585
R21811 DOUT[9].n1 DOUT[9].n0 185
R21812 DOUT[9].n2 DOUT[9] 51.9733
R21813 DOUT[9] DOUT[9].n1 49.0339
R21814 DOUT[9].n3 DOUT[9].t0 26.5955
R21815 DOUT[9].n3 DOUT[9].t1 26.5955
R21816 DOUT[9].n0 DOUT[9].t2 24.9236
R21817 DOUT[9].n0 DOUT[9].t3 24.9236
R21818 DOUT[9].n4 DOUT[9] 15.6165
R21819 DOUT[9].n1 DOUT[9] 10.4965
R21820 DOUT[9].n2 DOUT[9] 1.7925
R21821 DOUT[9] DOUT[9].n4 1.7925
R21822 a_2196_10927.n1 a_2196_10927.n0 926.024
R21823 a_2196_10927.n1 a_2196_10927.t3 82.0838
R21824 a_2196_10927.n0 a_2196_10927.t2 63.3338
R21825 a_2196_10927.t0 a_2196_10927.n1 63.3219
R21826 a_2196_10927.n0 a_2196_10927.t1 29.7268
R21827 a_8452_10749.n1 a_8452_10749.n0 926.024
R21828 a_8452_10749.t0 a_8452_10749.n1 82.0838
R21829 a_8452_10749.n0 a_8452_10749.t3 63.3338
R21830 a_8452_10749.n1 a_8452_10749.t1 63.3219
R21831 a_8452_10749.n0 a_8452_10749.t2 29.7268
R21832 a_9503_3861.n1 a_9503_3861.t2 530.01
R21833 a_9503_3861.t0 a_9503_3861.n5 421.021
R21834 a_9503_3861.n0 a_9503_3861.t3 337.142
R21835 a_9503_3861.n3 a_9503_3861.t1 280.223
R21836 a_9503_3861.n4 a_9503_3861.t5 263.173
R21837 a_9503_3861.n4 a_9503_3861.t6 227.826
R21838 a_9503_3861.n0 a_9503_3861.t4 199.762
R21839 a_9503_3861.n2 a_9503_3861.n1 170.81
R21840 a_9503_3861.n2 a_9503_3861.n0 167.321
R21841 a_9503_3861.n5 a_9503_3861.n4 152
R21842 a_9503_3861.n1 a_9503_3861.t7 141.923
R21843 a_9503_3861.n3 a_9503_3861.n2 10.8376
R21844 a_9503_3861.n5 a_9503_3861.n3 2.50485
R21845 a_10019_4233.n3 a_10019_4233.n2 674.338
R21846 a_10019_4233.n1 a_10019_4233.t5 332.58
R21847 a_10019_4233.n2 a_10019_4233.n0 284.012
R21848 a_10019_4233.n2 a_10019_4233.n1 253.648
R21849 a_10019_4233.n1 a_10019_4233.t4 168.701
R21850 a_10019_4233.t1 a_10019_4233.n3 96.1553
R21851 a_10019_4233.n3 a_10019_4233.t2 65.6672
R21852 a_10019_4233.n0 a_10019_4233.t0 65.0005
R21853 a_10019_4233.n0 a_10019_4233.t3 45.0005
R21854 a_10127_3855.n0 a_10127_3855.t2 1327.82
R21855 a_10127_3855.n0 a_10127_3855.t1 194.655
R21856 a_10127_3855.t0 a_10127_3855.n0 63.3219
R21857 a_4181_4399.t0 a_4181_4399.t1 87.1434
R21858 a_4421_8751.n0 a_4421_8751.t1 68.3338
R21859 a_4421_8751.n0 a_4421_8751.t0 26.3935
R21860 a_4421_8751.n1 a_4421_8751.n0 14.4005
R21861 a_4146_9003.n3 a_4146_9003.n2 636.953
R21862 a_4146_9003.n1 a_4146_9003.t4 366.856
R21863 a_4146_9003.n2 a_4146_9003.n0 300.2
R21864 a_4146_9003.n2 a_4146_9003.n1 225.036
R21865 a_4146_9003.n1 a_4146_9003.t5 174.056
R21866 a_4146_9003.n0 a_4146_9003.t0 70.0005
R21867 a_4146_9003.n3 a_4146_9003.t2 68.0124
R21868 a_4146_9003.t1 a_4146_9003.n3 63.3219
R21869 a_4146_9003.n0 a_4146_9003.t3 61.6672
R21870 a_8183_3285.n5 a_8183_3285.n4 807.871
R21871 a_8183_3285.n2 a_8183_3285.t5 389.183
R21872 a_8183_3285.n3 a_8183_3285.n2 251.167
R21873 a_8183_3285.n3 a_8183_3285.t1 223.571
R21874 a_8183_3285.n0 a_8183_3285.t8 212.081
R21875 a_8183_3285.n1 a_8183_3285.t6 212.081
R21876 a_8183_3285.n4 a_8183_3285.n1 176.576
R21877 a_8183_3285.n2 a_8183_3285.t3 174.891
R21878 a_8183_3285.n0 a_8183_3285.t4 139.78
R21879 a_8183_3285.n1 a_8183_3285.t7 139.78
R21880 a_8183_3285.n5 a_8183_3285.t2 63.3219
R21881 a_8183_3285.t0 a_8183_3285.n5 63.3219
R21882 a_8183_3285.n1 a_8183_3285.n0 61.346
R21883 a_8183_3285.n4 a_8183_3285.n3 37.7195
R21884 a_8117_3311.t1 a_8117_3311.t0 94.7268
R21885 a_5539_5724.n3 a_5539_5724.n2 674.338
R21886 a_5539_5724.n1 a_5539_5724.t4 332.58
R21887 a_5539_5724.n2 a_5539_5724.n0 284.012
R21888 a_5539_5724.n2 a_5539_5724.n1 253.648
R21889 a_5539_5724.n1 a_5539_5724.t5 168.701
R21890 a_5539_5724.t1 a_5539_5724.n3 96.1553
R21891 a_5539_5724.n3 a_5539_5724.t2 65.6672
R21892 a_5539_5724.n0 a_5539_5724.t0 65.0005
R21893 a_5539_5724.n0 a_5539_5724.t3 45.0005
R21894 a_5470_5853.n3 a_5470_5853.n2 647.119
R21895 a_5470_5853.n1 a_5470_5853.t4 350.253
R21896 a_5470_5853.n2 a_5470_5853.n0 260.339
R21897 a_5470_5853.n2 a_5470_5853.n1 246.119
R21898 a_5470_5853.n1 a_5470_5853.t5 189.588
R21899 a_5470_5853.n3 a_5470_5853.t0 89.1195
R21900 a_5470_5853.n0 a_5470_5853.t1 63.3338
R21901 a_5470_5853.t2 a_5470_5853.n3 41.0422
R21902 a_5470_5853.n0 a_5470_5853.t3 31.9797
R21903 a_7348_3311.n1 a_7348_3311.n0 926.024
R21904 a_7348_3311.t1 a_7348_3311.n1 82.0838
R21905 a_7348_3311.n0 a_7348_3311.t0 63.3338
R21906 a_7348_3311.n1 a_7348_3311.t2 63.3219
R21907 a_7348_3311.n0 a_7348_3311.t3 29.7268
R21908 a_6573_6575.t0 a_6573_6575.t1 87.1434
R21909 a_7443_3311.n3 a_7443_3311.n2 674.338
R21910 a_7443_3311.n1 a_7443_3311.t4 332.58
R21911 a_7443_3311.n2 a_7443_3311.n0 284.012
R21912 a_7443_3311.n2 a_7443_3311.n1 253.648
R21913 a_7443_3311.n1 a_7443_3311.t5 168.701
R21914 a_7443_3311.t1 a_7443_3311.n3 96.1553
R21915 a_7443_3311.n3 a_7443_3311.t3 65.6672
R21916 a_7443_3311.n0 a_7443_3311.t0 65.0005
R21917 a_7443_3311.n0 a_7443_3311.t2 45.0005
R21918 a_7661_3553.n3 a_7661_3553.n2 647.119
R21919 a_7661_3553.n1 a_7661_3553.t5 350.253
R21920 a_7661_3553.n2 a_7661_3553.n0 260.339
R21921 a_7661_3553.n2 a_7661_3553.n1 246.119
R21922 a_7661_3553.n1 a_7661_3553.t4 189.588
R21923 a_7661_3553.n3 a_7661_3553.t2 89.1195
R21924 a_7661_3553.n0 a_7661_3553.t3 63.3338
R21925 a_7661_3553.t0 a_7661_3553.n3 41.0422
R21926 a_7661_3553.n0 a_7661_3553.t1 31.9797
R21927 a_7981_4221.t0 a_7981_4221.t1 60.0005
R21928 a_7539_3311.t0 a_7539_3311.t1 198.571
R21929 a_9503_2773.n1 a_9503_2773.t6 530.01
R21930 a_9503_2773.t0 a_9503_2773.n5 421.021
R21931 a_9503_2773.n0 a_9503_2773.t7 337.142
R21932 a_9503_2773.n3 a_9503_2773.t1 280.223
R21933 a_9503_2773.n4 a_9503_2773.t3 263.173
R21934 a_9503_2773.n4 a_9503_2773.t4 227.826
R21935 a_9503_2773.n0 a_9503_2773.t2 199.762
R21936 a_9503_2773.n2 a_9503_2773.n1 170.81
R21937 a_9503_2773.n2 a_9503_2773.n0 167.321
R21938 a_9503_2773.n5 a_9503_2773.n4 152
R21939 a_9503_2773.n1 a_9503_2773.t5 141.923
R21940 a_9503_2773.n3 a_9503_2773.n2 10.8376
R21941 a_9503_2773.n5 a_9503_2773.n3 2.50485
R21942 a_7125_3133.t0 a_7125_3133.t1 87.1434
R21943 SWN[8].n2 SWN[8].n1 585
R21944 SWN[8].n1 SWN[8].n0 585
R21945 SWN[8].n4 SWN[8].n3 185
R21946 SWN[8].n4 SWN[8] 57.7379
R21947 SWN[8].n1 SWN[8].t1 26.5955
R21948 SWN[8].n1 SWN[8].t0 26.5955
R21949 SWN[8].n3 SWN[8].t2 24.9236
R21950 SWN[8].n3 SWN[8].t3 24.9236
R21951 SWN[8] SWN[8].n2 10.4965
R21952 SWN[8].n0 SWN[8] 10.4965
R21953 SWN[8].n2 SWN[8] 6.9125
R21954 SWN[8].n0 SWN[8] 6.9125
R21955 SWN[8] SWN[8].n4 1.7925
R21956 a_5015_6273.n1 a_5015_6273.t2 530.01
R21957 a_5015_6273.t0 a_5015_6273.n5 421.021
R21958 a_5015_6273.n0 a_5015_6273.t5 337.171
R21959 a_5015_6273.n3 a_5015_6273.t1 280.223
R21960 a_5015_6273.n4 a_5015_6273.t4 263.173
R21961 a_5015_6273.n4 a_5015_6273.t6 227.826
R21962 a_5015_6273.n0 a_5015_6273.t3 199.762
R21963 a_5015_6273.n2 a_5015_6273.n1 170.81
R21964 a_5015_6273.n2 a_5015_6273.n0 167.321
R21965 a_5015_6273.n5 a_5015_6273.n4 152
R21966 a_5015_6273.n1 a_5015_6273.t7 141.923
R21967 a_5015_6273.n3 a_5015_6273.n2 10.8376
R21968 a_5015_6273.n5 a_5015_6273.n3 2.50485
R21969 a_5316_6031.t0 a_5316_6031.n0 1327.82
R21970 a_5316_6031.n0 a_5316_6031.t2 194.655
R21971 a_5316_6031.n0 a_5316_6031.t1 63.3219
R21972 a_5171_6005.n3 a_5171_6005.n2 674.338
R21973 a_5171_6005.n1 a_5171_6005.t4 332.58
R21974 a_5171_6005.n2 a_5171_6005.n0 284.012
R21975 a_5171_6005.n2 a_5171_6005.n1 253.648
R21976 a_5171_6005.n1 a_5171_6005.t5 168.701
R21977 a_5171_6005.n3 a_5171_6005.t3 96.1553
R21978 a_5171_6005.t0 a_5171_6005.n3 65.6672
R21979 a_5171_6005.n0 a_5171_6005.t2 65.0005
R21980 a_5171_6005.n0 a_5171_6005.t1 45.0005
R21981 a_7407_8893.n1 a_7407_8893.t4 530.01
R21982 a_7407_8893.t0 a_7407_8893.n5 421.021
R21983 a_7407_8893.n0 a_7407_8893.t2 337.171
R21984 a_7407_8893.n3 a_7407_8893.t1 280.223
R21985 a_7407_8893.n4 a_7407_8893.t6 263.173
R21986 a_7407_8893.n4 a_7407_8893.t3 227.826
R21987 a_7407_8893.n0 a_7407_8893.t7 199.762
R21988 a_7407_8893.n2 a_7407_8893.n1 170.81
R21989 a_7407_8893.n2 a_7407_8893.n0 167.321
R21990 a_7407_8893.n5 a_7407_8893.n4 152
R21991 a_7407_8893.n1 a_7407_8893.t5 141.923
R21992 a_7407_8893.n3 a_7407_8893.n2 10.8376
R21993 a_7407_8893.n5 a_7407_8893.n3 2.50485
R21994 a_10492_5321.n3 a_10492_5321.n2 636.953
R21995 a_10492_5321.n1 a_10492_5321.t4 366.856
R21996 a_10492_5321.n2 a_10492_5321.n0 300.2
R21997 a_10492_5321.n2 a_10492_5321.n1 225.036
R21998 a_10492_5321.n1 a_10492_5321.t5 174.056
R21999 a_10492_5321.n0 a_10492_5321.t3 70.0005
R22000 a_10492_5321.t0 a_10492_5321.n3 68.0124
R22001 a_10492_5321.n3 a_10492_5321.t2 63.3219
R22002 a_10492_5321.n0 a_10492_5321.t1 61.6672
R22003 a_10846_5309.t0 a_10846_5309.t1 87.1434
R22004 a_2526_5853.n3 a_2526_5853.n2 647.119
R22005 a_2526_5853.n1 a_2526_5853.t5 350.253
R22006 a_2526_5853.n2 a_2526_5853.n0 260.339
R22007 a_2526_5853.n2 a_2526_5853.n1 246.119
R22008 a_2526_5853.n1 a_2526_5853.t4 189.588
R22009 a_2526_5853.n3 a_2526_5853.t2 89.1195
R22010 a_2526_5853.n0 a_2526_5853.t3 63.3338
R22011 a_2526_5853.t0 a_2526_5853.n3 41.0422
R22012 a_2526_5853.n0 a_2526_5853.t1 31.9797
R22013 a_2740_5853.t0 a_2740_5853.n0 1327.82
R22014 a_2740_5853.n0 a_2740_5853.t1 194.655
R22015 a_2740_5853.n0 a_2740_5853.t2 63.3219
R22016 a_3662_11471.t0 a_3662_11471.t1 126.644
R22017 a_10693_6409.n0 a_10693_6409.t0 68.3338
R22018 a_10693_6409.n0 a_10693_6409.t1 26.3935
R22019 a_10693_6409.n1 a_10693_6409.n0 14.4005
R22020 DOUT[7].n4 DOUT[7].n3 585
R22021 DOUT[7].n3 DOUT[7].n2 585
R22022 DOUT[7].n1 DOUT[7].n0 185
R22023 DOUT[7].n5 DOUT[7].n1 53.3859
R22024 DOUT[7].n3 DOUT[7].t1 26.5955
R22025 DOUT[7].n3 DOUT[7].t0 26.5955
R22026 DOUT[7].n0 DOUT[7].t3 24.9236
R22027 DOUT[7].n0 DOUT[7].t2 24.9236
R22028 DOUT[7] DOUT[7].n5 11.7141
R22029 DOUT[7] DOUT[7].n4 10.4965
R22030 DOUT[7].n2 DOUT[7] 10.4965
R22031 DOUT[7].n4 DOUT[7] 6.9125
R22032 DOUT[7].n2 DOUT[7] 6.9125
R22033 DOUT[7].n5 DOUT[7] 4.3525
R22034 DOUT[7].n1 DOUT[7] 1.7925
R22035 a_4883_3855.n0 a_4883_3855.t1 1327.82
R22036 a_4883_3855.t0 a_4883_3855.n0 194.655
R22037 a_4883_3855.n0 a_4883_3855.t2 63.3219
R22038 a_4089_8573.t0 a_4089_8573.t1 87.1434
R22039 a_10207_8725.n5 a_10207_8725.n4 807.871
R22040 a_10207_8725.n2 a_10207_8725.t7 389.183
R22041 a_10207_8725.n3 a_10207_8725.n2 251.167
R22042 a_10207_8725.n3 a_10207_8725.t1 223.571
R22043 a_10207_8725.n0 a_10207_8725.t3 212.081
R22044 a_10207_8725.n1 a_10207_8725.t8 212.081
R22045 a_10207_8725.n4 a_10207_8725.n1 176.576
R22046 a_10207_8725.n2 a_10207_8725.t4 174.891
R22047 a_10207_8725.n0 a_10207_8725.t6 139.78
R22048 a_10207_8725.n1 a_10207_8725.t5 139.78
R22049 a_10207_8725.n5 a_10207_8725.t2 63.3219
R22050 a_10207_8725.t0 a_10207_8725.n5 63.3219
R22051 a_10207_8725.n1 a_10207_8725.n0 61.346
R22052 a_10207_8725.n4 a_10207_8725.n3 37.7195
R22053 DOUT[2].n3 DOUT[2].n2 585
R22054 DOUT[2].n4 DOUT[2].n3 585
R22055 DOUT[2].n1 DOUT[2].n0 185
R22056 DOUT[2] DOUT[2].n1 49.0339
R22057 DOUT[2].n3 DOUT[2].t1 26.5955
R22058 DOUT[2].n3 DOUT[2].t0 26.5955
R22059 DOUT[2].n0 DOUT[2].t2 24.9236
R22060 DOUT[2].n0 DOUT[2].t3 24.9236
R22061 DOUT[2].n2 DOUT[2] 15.6165
R22062 DOUT[2] DOUT[2].n4 12.0152
R22063 DOUT[2].n1 DOUT[2] 10.4965
R22064 DOUT[2].n4 DOUT[2] 1.7925
R22065 DOUT[2].n2 DOUT[2] 1.7925
R22066 a_5340_4233.n3 a_5340_4233.n2 636.953
R22067 a_5340_4233.n1 a_5340_4233.t4 366.856
R22068 a_5340_4233.n2 a_5340_4233.n0 300.2
R22069 a_5340_4233.n2 a_5340_4233.n1 225.036
R22070 a_5340_4233.n1 a_5340_4233.t5 174.056
R22071 a_5340_4233.n0 a_5340_4233.t2 70.0005
R22072 a_5340_4233.t1 a_5340_4233.n3 68.0124
R22073 a_5340_4233.n3 a_5340_4233.t3 63.3219
R22074 a_5340_4233.n0 a_5340_4233.t0 61.6672
R22075 a_8008_3311.n3 a_8008_3311.n2 636.953
R22076 a_8008_3311.n1 a_8008_3311.t4 366.856
R22077 a_8008_3311.n2 a_8008_3311.n0 300.2
R22078 a_8008_3311.n2 a_8008_3311.n1 225.036
R22079 a_8008_3311.n1 a_8008_3311.t5 174.056
R22080 a_8008_3311.n0 a_8008_3311.t2 70.0005
R22081 a_8008_3311.t0 a_8008_3311.n3 68.0124
R22082 a_8008_3311.n3 a_8008_3311.t3 63.3219
R22083 a_8008_3311.n0 a_8008_3311.t1 61.6672
R22084 a_10838_3677.t0 a_10838_3677.t1 126.644
R22085 a_2032_9019.t0 a_2032_9019.n3 370.026
R22086 a_2032_9019.n0 a_2032_9019.t5 351.356
R22087 a_2032_9019.n1 a_2032_9019.t2 334.717
R22088 a_2032_9019.n3 a_2032_9019.t1 325.971
R22089 a_2032_9019.n1 a_2032_9019.t4 309.935
R22090 a_2032_9019.n0 a_2032_9019.t3 305.683
R22091 a_2032_9019.n2 a_2032_9019.n0 16.879
R22092 a_2032_9019.n3 a_2032_9019.n2 10.8867
R22093 a_2032_9019.n2 a_2032_9019.n1 9.3005
R22094 a_2537_8751.t1 a_2537_8751.t0 198.571
R22095 a_2227_8988.n3 a_2227_8988.n2 674.338
R22096 a_2227_8988.n1 a_2227_8988.t4 332.58
R22097 a_2227_8988.n2 a_2227_8988.n0 284.012
R22098 a_2227_8988.n2 a_2227_8988.n1 253.648
R22099 a_2227_8988.n1 a_2227_8988.t5 168.701
R22100 a_2227_8988.n3 a_2227_8988.t2 96.1553
R22101 a_2227_8988.t1 a_2227_8988.n3 65.6672
R22102 a_2227_8988.n0 a_2227_8988.t3 65.0005
R22103 a_2227_8988.n0 a_2227_8988.t0 45.0005
R22104 a_5081_12015.t1 a_5081_12015.t0 94.7268
R22105 a_7203_3861.n1 a_7203_3861.t7 530.01
R22106 a_7203_3861.t0 a_7203_3861.n5 421.021
R22107 a_7203_3861.n0 a_7203_3861.t2 337.142
R22108 a_7203_3861.n3 a_7203_3861.t1 280.223
R22109 a_7203_3861.n4 a_7203_3861.t3 263.173
R22110 a_7203_3861.n4 a_7203_3861.t5 227.826
R22111 a_7203_3861.n0 a_7203_3861.t4 199.762
R22112 a_7203_3861.n2 a_7203_3861.n1 170.81
R22113 a_7203_3861.n2 a_7203_3861.n0 167.321
R22114 a_7203_3861.n5 a_7203_3861.n4 152
R22115 a_7203_3861.n1 a_7203_3861.t6 141.923
R22116 a_7203_3861.n3 a_7203_3861.n2 10.8376
R22117 a_7203_3861.n5 a_7203_3861.n3 2.50485
R22118 a_10654_4943.t0 a_10654_4943.t1 126.644
R22119 a_4669_12015.t0 a_4669_12015.t1 60.0005
R22120 a_4976_6147.t0 a_4976_6147.n3 370.026
R22121 a_4976_6147.n0 a_4976_6147.t5 351.356
R22122 a_4976_6147.n1 a_4976_6147.t4 334.717
R22123 a_4976_6147.n3 a_4976_6147.t1 325.971
R22124 a_4976_6147.n1 a_4976_6147.t2 309.935
R22125 a_4976_6147.n0 a_4976_6147.t3 305.683
R22126 a_4976_6147.n2 a_4976_6147.n0 16.879
R22127 a_4976_6147.n3 a_4976_6147.n2 10.8867
R22128 a_4976_6147.n2 a_4976_6147.n1 9.3005
R22129 a_5734_6031.n1 a_5734_6031.n0 926.024
R22130 a_5734_6031.n1 a_5734_6031.t2 82.0838
R22131 a_5734_6031.n0 a_5734_6031.t3 63.3338
R22132 a_5734_6031.t0 a_5734_6031.n1 63.3219
R22133 a_5734_6031.n0 a_5734_6031.t1 29.7268
R22134 a_5734_11471.n1 a_5734_11471.n0 926.024
R22135 a_5734_11471.t0 a_5734_11471.n1 82.0838
R22136 a_5734_11471.n0 a_5734_11471.t1 63.3338
R22137 a_5734_11471.n1 a_5734_11471.t2 63.3219
R22138 a_5734_11471.n0 a_5734_11471.t3 29.7268
R22139 a_8209_6409.n0 a_8209_6409.t1 68.3338
R22140 a_8209_6409.n0 a_8209_6409.t0 26.3935
R22141 a_8209_6409.n1 a_8209_6409.n0 14.4005
R22142 a_5090_8207.n1 a_5090_8207.n0 926.024
R22143 a_5090_8207.t1 a_5090_8207.n1 82.0838
R22144 a_5090_8207.n0 a_5090_8207.t0 63.3338
R22145 a_5090_8207.n1 a_5090_8207.t2 63.3219
R22146 a_5090_8207.n0 a_5090_8207.t3 29.7268
R22147 a_8126_9117.n1 a_8126_9117.n0 926.024
R22148 a_8126_9117.n1 a_8126_9117.t3 82.0838
R22149 a_8126_9117.n0 a_8126_9117.t0 63.3338
R22150 a_8126_9117.t1 a_8126_9117.n1 63.3219
R22151 a_8126_9117.n0 a_8126_9117.t2 29.7268
R22152 a_10237_2741.n3 a_10237_2741.n2 647.119
R22153 a_10237_2741.n1 a_10237_2741.t5 350.253
R22154 a_10237_2741.n2 a_10237_2741.n0 260.339
R22155 a_10237_2741.n2 a_10237_2741.n1 246.119
R22156 a_10237_2741.n1 a_10237_2741.t4 189.588
R22157 a_10237_2741.n3 a_10237_2741.t1 89.1195
R22158 a_10237_2741.n0 a_10237_2741.t0 63.3338
R22159 a_10237_2741.t3 a_10237_2741.n3 41.0422
R22160 a_10237_2741.n0 a_10237_2741.t2 31.9797
R22161 a_10127_2767.t0 a_10127_2767.n0 1327.82
R22162 a_10127_2767.n0 a_10127_2767.t2 194.655
R22163 a_10127_2767.n0 a_10127_2767.t1 63.3219
R22164 a_7440_6397.n1 a_7440_6397.n0 926.024
R22165 a_7440_6397.n1 a_7440_6397.t3 82.0838
R22166 a_7440_6397.n0 a_7440_6397.t2 63.3338
R22167 a_7440_6397.t0 a_7440_6397.n1 63.3219
R22168 a_7440_6397.n0 a_7440_6397.t1 29.7268
R22169 a_7535_6409.n3 a_7535_6409.n2 674.338
R22170 a_7535_6409.n1 a_7535_6409.t5 332.58
R22171 a_7535_6409.n2 a_7535_6409.n0 284.012
R22172 a_7535_6409.n2 a_7535_6409.n1 253.648
R22173 a_7535_6409.n1 a_7535_6409.t4 168.701
R22174 a_7535_6409.t1 a_7535_6409.n3 96.1553
R22175 a_7535_6409.n3 a_7535_6409.t2 65.6672
R22176 a_7535_6409.n0 a_7535_6409.t0 65.0005
R22177 a_7535_6409.n0 a_7535_6409.t3 45.0005
R22178 SWP[5].n6 SWP[5].n5 585
R22179 SWP[5].n5 SWP[5].n4 585
R22180 SWP[5].n0 SWP[5].t5 333.651
R22181 SWP[5].n0 SWP[5].t4 297.233
R22182 SWP[5].n1 SWP[5].n0 193.506
R22183 SWP[5].n3 SWP[5].n2 185
R22184 SWP[5].n8 SWP[5].n1 58.0758
R22185 SWP[5].n7 SWP[5].n3 53.3859
R22186 SWP[5].n5 SWP[5].t1 26.5955
R22187 SWP[5].n5 SWP[5].t0 26.5955
R22188 SWP[5].n2 SWP[5].t2 24.9236
R22189 SWP[5].n2 SWP[5].t3 24.9236
R22190 SWP[5] SWP[5].n8 16.4812
R22191 SWP[5] SWP[5].n6 10.4965
R22192 SWP[5].n4 SWP[5] 10.4965
R22193 SWP[5].n8 SWP[5].n7 9.3005
R22194 SWP[5].n6 SWP[5] 6.9125
R22195 SWP[5].n4 SWP[5] 6.9125
R22196 SWP[5].n7 SWP[5] 4.3525
R22197 SWP[5].n1 SWP[5] 4.17441
R22198 SWP[5].n3 SWP[5] 1.7925
R22199 a_5409_6397.t0 a_5409_6397.t1 60.0005
R22200 a_8362_10927.t0 a_8362_10927.t1 87.1434
R22201 a_9467_7663.n3 a_9467_7663.n2 674.338
R22202 a_9467_7663.n1 a_9467_7663.t4 332.58
R22203 a_9467_7663.n2 a_9467_7663.n0 284.012
R22204 a_9467_7663.n2 a_9467_7663.n1 253.648
R22205 a_9467_7663.n1 a_9467_7663.t5 168.701
R22206 a_9467_7663.n3 a_9467_7663.t3 96.1553
R22207 a_9467_7663.t0 a_9467_7663.n3 65.6672
R22208 a_9467_7663.n0 a_9467_7663.t2 65.0005
R22209 a_9467_7663.n0 a_9467_7663.t1 45.0005
R22210 a_5458_10383.n1 a_5458_10383.n0 926.024
R22211 a_5458_10383.n1 a_5458_10383.t3 82.0838
R22212 a_5458_10383.n0 a_5458_10383.t2 63.3338
R22213 a_5458_10383.t0 a_5458_10383.n1 63.3219
R22214 a_5458_10383.n0 a_5458_10383.t1 29.7268
R22215 x2/TRIG2.n0 x2/TRIG2.t3 333.651
R22216 x2/TRIG2.n0 x2/TRIG2.t2 297.233
R22217 x2/TRIG2 x2/TRIG2.t0 230.518
R22218 x2/TRIG2.n1 x2/TRIG2.n0 193.506
R22219 x2/TRIG2.n2 x2/TRIG2.t1 130.594
R22220 x2/TRIG2.n2 x2/TRIG2 33.1945
R22221 x2/TRIG2 x2/TRIG2.n2 31.7575
R22222 x2/TRIG2 x2/TRIG2.n1 26.5122
R22223 x2/TRIG2.n3 x2/TRIG2 11.6875
R22224 x2/TRIG2.n3 x2/TRIG2 7.23528
R22225 x2/TRIG2 x2/TRIG2.n3 5.04292
R22226 x2/TRIG2.n1 x2/TRIG2 4.17441
R22227 a_9467_10927.n3 a_9467_10927.n2 674.338
R22228 a_9467_10927.n1 a_9467_10927.t5 332.58
R22229 a_9467_10927.n2 a_9467_10927.n0 284.012
R22230 a_9467_10927.n2 a_9467_10927.n1 253.648
R22231 a_9467_10927.n1 a_9467_10927.t4 168.701
R22232 a_9467_10927.n3 a_9467_10927.t2 96.1553
R22233 a_9467_10927.t0 a_9467_10927.n3 65.6672
R22234 a_9467_10927.n0 a_9467_10927.t1 65.0005
R22235 a_9467_10927.n0 a_9467_10927.t3 45.0005
R22236 a_9685_11169.n3 a_9685_11169.n2 647.119
R22237 a_9685_11169.n1 a_9685_11169.t5 350.253
R22238 a_9685_11169.n2 a_9685_11169.n0 260.339
R22239 a_9685_11169.n2 a_9685_11169.n1 246.119
R22240 a_9685_11169.n1 a_9685_11169.t4 189.588
R22241 a_9685_11169.n3 a_9685_11169.t0 89.1195
R22242 a_9685_11169.n0 a_9685_11169.t3 63.3338
R22243 a_9685_11169.t1 a_9685_11169.n3 41.0422
R22244 a_9685_11169.n0 a_9685_11169.t2 31.9797
R22245 a_6467_11477.n1 a_6467_11477.t7 530.01
R22246 a_6467_11477.t0 a_6467_11477.n5 421.021
R22247 a_6467_11477.n0 a_6467_11477.t6 337.142
R22248 a_6467_11477.n3 a_6467_11477.t1 280.223
R22249 a_6467_11477.n4 a_6467_11477.t3 263.173
R22250 a_6467_11477.n4 a_6467_11477.t5 227.826
R22251 a_6467_11477.n0 a_6467_11477.t2 199.762
R22252 a_6467_11477.n2 a_6467_11477.n1 170.81
R22253 a_6467_11477.n2 a_6467_11477.n0 167.321
R22254 a_6467_11477.n5 a_6467_11477.n4 152
R22255 a_6467_11477.n1 a_6467_11477.t4 141.923
R22256 a_6467_11477.n3 a_6467_11477.n2 10.8376
R22257 a_6467_11477.n5 a_6467_11477.n3 2.50485
R22258 a_7548_11849.n3 a_7548_11849.n2 636.953
R22259 a_7548_11849.n1 a_7548_11849.t4 366.856
R22260 a_7548_11849.n2 a_7548_11849.n0 300.2
R22261 a_7548_11849.n2 a_7548_11849.n1 225.036
R22262 a_7548_11849.n1 a_7548_11849.t5 174.056
R22263 a_7548_11849.n0 a_7548_11849.t2 70.0005
R22264 a_7548_11849.t1 a_7548_11849.n3 68.0124
R22265 a_7548_11849.n3 a_7548_11849.t3 63.3219
R22266 a_7548_11849.n0 a_7548_11849.t0 61.6672
R22267 a_7657_11849.n0 a_7657_11849.t1 68.3338
R22268 a_7657_11849.n0 a_7657_11849.t0 26.3935
R22269 a_7657_11849.n1 a_7657_11849.n0 14.4005
R22270 a_6927_10927.n1 a_6927_10927.t2 530.01
R22271 a_6927_10927.t0 a_6927_10927.n5 421.021
R22272 a_6927_10927.n0 a_6927_10927.t7 337.142
R22273 a_6927_10927.n3 a_6927_10927.t1 280.223
R22274 a_6927_10927.n4 a_6927_10927.t5 263.173
R22275 a_6927_10927.n4 a_6927_10927.t4 227.826
R22276 a_6927_10927.n0 a_6927_10927.t6 199.762
R22277 a_6927_10927.n2 a_6927_10927.n1 170.81
R22278 a_6927_10927.n2 a_6927_10927.n0 167.321
R22279 a_6927_10927.n5 a_6927_10927.n4 152
R22280 a_6927_10927.n1 a_6927_10927.t3 141.923
R22281 a_6927_10927.n3 a_6927_10927.n2 10.8376
R22282 a_6927_10927.n5 a_6927_10927.n3 2.50485
R22283 a_7443_10927.n3 a_7443_10927.n2 674.338
R22284 a_7443_10927.n1 a_7443_10927.t4 332.58
R22285 a_7443_10927.n2 a_7443_10927.n0 284.012
R22286 a_7443_10927.n2 a_7443_10927.n1 253.648
R22287 a_7443_10927.n1 a_7443_10927.t5 168.701
R22288 a_7443_10927.t1 a_7443_10927.n3 96.1553
R22289 a_7443_10927.n3 a_7443_10927.t2 65.6672
R22290 a_7443_10927.n0 a_7443_10927.t0 65.0005
R22291 a_7443_10927.n0 a_7443_10927.t3 45.0005
R22292 a_7643_6031.t0 a_7643_6031.n0 1327.82
R22293 a_7643_6031.n0 a_7643_6031.t2 194.655
R22294 a_7643_6031.n0 a_7643_6031.t1 63.3219
R22295 a_9927_9839.n3 a_9927_9839.n2 674.338
R22296 a_9927_9839.n1 a_9927_9839.t5 332.58
R22297 a_9927_9839.n2 a_9927_9839.n0 284.012
R22298 a_9927_9839.n2 a_9927_9839.n1 253.648
R22299 a_9927_9839.n1 a_9927_9839.t4 168.701
R22300 a_9927_9839.t1 a_9927_9839.n3 96.1553
R22301 a_9927_9839.n3 a_9927_9839.t2 65.6672
R22302 a_9927_9839.n0 a_9927_9839.t0 65.0005
R22303 a_9927_9839.n0 a_9927_9839.t3 45.0005
R22304 a_10023_9839.t0 a_10023_9839.t1 198.571
R22305 a_9924_4221.n1 a_9924_4221.n0 926.024
R22306 a_9924_4221.n1 a_9924_4221.t3 82.0838
R22307 a_9924_4221.n0 a_9924_4221.t0 63.3338
R22308 a_9924_4221.t1 a_9924_4221.n1 63.3219
R22309 a_9924_4221.n0 a_9924_4221.t2 29.7268
R22310 SWP[9].n4 SWP[9].t4 332.312
R22311 SWP[9].n4 SWP[9].t5 295.627
R22312 SWP[9].n1 SWP[9].n0 289.096
R22313 SWP[9] SWP[9].n4 195.401
R22314 SWP[9].n3 SWP[9].n2 185
R22315 SWP[9].n5 SWP[9] 54.8293
R22316 SWP[9].n3 SWP[9] 49.0339
R22317 SWP[9].n5 SWP[9] 28.3116
R22318 SWP[9].n0 SWP[9].t1 26.5955
R22319 SWP[9].n0 SWP[9].t0 26.5955
R22320 SWP[9].n2 SWP[9].t2 24.9236
R22321 SWP[9].n2 SWP[9].t3 24.9236
R22322 SWP[9].n6 SWP[9].n5 12.8803
R22323 SWP[9] SWP[9].n1 9.48653
R22324 SWP[9].n1 SWP[9] 7.7181
R22325 SWP[9].n6 SWP[9].n3 6.1445
R22326 SWP[9] SWP[9].n6 4.3525
R22327 a_6816_6843.t0 a_6816_6843.n3 370.026
R22328 a_6816_6843.n0 a_6816_6843.t5 351.356
R22329 a_6816_6843.n1 a_6816_6843.t3 334.717
R22330 a_6816_6843.n3 a_6816_6843.t1 325.971
R22331 a_6816_6843.n1 a_6816_6843.t2 309.935
R22332 a_6816_6843.n0 a_6816_6843.t4 305.683
R22333 a_6816_6843.n2 a_6816_6843.n0 16.879
R22334 a_6816_6843.n3 a_6816_6843.n2 10.8867
R22335 a_6816_6843.n2 a_6816_6843.n1 9.3005
R22336 a_7574_6941.n1 a_7574_6941.n0 926.024
R22337 a_7574_6941.n1 a_7574_6941.t2 82.0838
R22338 a_7574_6941.n0 a_7574_6941.t3 63.3338
R22339 a_7574_6941.t0 a_7574_6941.n1 63.3219
R22340 a_7574_6941.n0 a_7574_6941.t1 29.7268
R22341 a_6996_7663.n3 a_6996_7663.n2 636.953
R22342 a_6996_7663.n1 a_6996_7663.t4 366.856
R22343 a_6996_7663.n2 a_6996_7663.n0 300.2
R22344 a_6996_7663.n2 a_6996_7663.n1 225.036
R22345 a_6996_7663.n1 a_6996_7663.t5 174.056
R22346 a_6996_7663.n0 a_6996_7663.t3 70.0005
R22347 a_6996_7663.t1 a_6996_7663.n3 68.0124
R22348 a_6996_7663.n3 a_6996_7663.t2 63.3219
R22349 a_6996_7663.n0 a_6996_7663.t0 61.6672
R22350 a_7350_7663.t0 a_7350_7663.t1 87.1434
R22351 a_4995_10927.n1 a_4995_10927.t4 530.01
R22352 a_4995_10927.t0 a_4995_10927.n5 421.021
R22353 a_4995_10927.n0 a_4995_10927.t3 337.142
R22354 a_4995_10927.n3 a_4995_10927.t1 280.223
R22355 a_4995_10927.n4 a_4995_10927.t7 263.173
R22356 a_4995_10927.n4 a_4995_10927.t6 227.826
R22357 a_4995_10927.n0 a_4995_10927.t2 199.762
R22358 a_4995_10927.n2 a_4995_10927.n1 170.81
R22359 a_4995_10927.n2 a_4995_10927.n0 167.321
R22360 a_4995_10927.n5 a_4995_10927.n4 152
R22361 a_4995_10927.n1 a_4995_10927.t5 141.923
R22362 a_4995_10927.n3 a_4995_10927.n2 10.8376
R22363 a_4995_10927.n5 a_4995_10927.n3 2.50485
R22364 a_6185_10927.t0 a_6185_10927.t1 94.7268
R22365 x2/net12.n2 x2/net12.t9 212.081
R22366 x2/net12.n10 x2/net12.t5 212.081
R22367 x2/net12.n3 x2/net12.t7 212.081
R22368 x2/net12.n5 x2/net12.t8 212.081
R22369 x2/net12.n15 x2/net12.n14 208.965
R22370 x2/net12.n5 x2/net12.n4 188.516
R22371 x2/net12.n7 x2/net12.n6 152
R22372 x2/net12.n9 x2/net12.n8 152
R22373 x2/net12.n12 x2/net12.n11 152
R22374 x2/net12.n2 x2/net12.t4 139.78
R22375 x2/net12.n10 x2/net12.t11 139.78
R22376 x2/net12.n3 x2/net12.t6 139.78
R22377 x2/net12.n5 x2/net12.t10 139.78
R22378 x2/net12 x2/net12.n0 96.8352
R22379 x2/net12.n11 x2/net12.n2 30.6732
R22380 x2/net12.n11 x2/net12.n10 30.6732
R22381 x2/net12.n10 x2/net12.n9 30.6732
R22382 x2/net12.n9 x2/net12.n3 30.6732
R22383 x2/net12.n6 x2/net12.n3 30.6732
R22384 x2/net12.n6 x2/net12.n5 30.6732
R22385 x2/net12.n14 x2/net12.t1 26.5955
R22386 x2/net12.n14 x2/net12.t0 26.5955
R22387 x2/net12.n0 x2/net12.t3 24.9236
R22388 x2/net12.n0 x2/net12.t2 24.9236
R22389 x2/net12.n8 x2/net12 19.2005
R22390 x2/net12 x2/net12.n7 17.1525
R22391 x2/net12.n4 x2/net12 17.1525
R22392 x2/net12 x2/net12.n13 13.0565
R22393 x2/net12 x2/net12.n12 11.9139
R22394 x2/net12 x2/net12.n1 11.2645
R22395 x2/net12.n13 x2/net12 9.86591
R22396 x2/net12.n7 x2/net12 6.4005
R22397 x2/net12.n4 x2/net12 6.4005
R22398 x2/net12.n1 x2/net12 6.1445
R22399 x2/net12.n1 x2/net12 4.65505
R22400 x2/net12.n8 x2/net12 4.3525
R22401 x2/net12.n13 x2/net12 4.3525
R22402 x2/net12.n12 x2/net12 2.3045
R22403 x2/net12.n15 x2/net12 2.0485
R22404 x2/net12 x2/net12.n15 1.55202
R22405 a_7369_3861.t0 a_7369_3861.n3 370.026
R22406 a_7369_3861.n0 a_7369_3861.t5 351.356
R22407 a_7369_3861.n1 a_7369_3861.t3 334.717
R22408 a_7369_3861.n3 a_7369_3861.t1 325.971
R22409 a_7369_3861.n1 a_7369_3861.t4 309.935
R22410 a_7369_3861.n0 a_7369_3861.t2 305.683
R22411 a_7369_3861.n2 a_7369_3861.n0 16.879
R22412 a_7369_3861.n3 a_7369_3861.n2 10.8867
R22413 a_7369_3861.n2 a_7369_3861.n1 9.3005
R22414 a_8446_3855.t0 a_8446_3855.t1 126.644
R22415 a_10035_4943.n0 a_10035_4943.t1 1327.82
R22416 a_10035_4943.t0 a_10035_4943.n0 194.655
R22417 a_10035_4943.n0 a_10035_4943.t2 63.3219
R22418 a_2439_9981.n1 a_2439_9981.t6 530.01
R22419 a_2439_9981.t0 a_2439_9981.n5 421.021
R22420 a_2439_9981.n0 a_2439_9981.t5 337.171
R22421 a_2439_9981.n3 a_2439_9981.t1 280.223
R22422 a_2439_9981.n4 a_2439_9981.t3 263.173
R22423 a_2439_9981.n4 a_2439_9981.t2 227.826
R22424 a_2439_9981.n0 a_2439_9981.t7 199.762
R22425 a_2439_9981.n2 a_2439_9981.n1 170.81
R22426 a_2439_9981.n2 a_2439_9981.n0 167.321
R22427 a_2439_9981.n5 a_2439_9981.n4 152
R22428 a_2439_9981.n1 a_2439_9981.t4 141.923
R22429 a_2439_9981.n3 a_2439_9981.n2 10.8376
R22430 a_2439_9981.n5 a_2439_9981.n3 2.50485
R22431 DOUT[1].n3 DOUT[1].n2 585
R22432 DOUT[1].n4 DOUT[1].n3 585
R22433 DOUT[1].n1 DOUT[1].n0 185
R22434 DOUT[1] DOUT[1].n1 49.0339
R22435 DOUT[1].n3 DOUT[1].t1 26.5955
R22436 DOUT[1].n3 DOUT[1].t0 26.5955
R22437 DOUT[1].n0 DOUT[1].t3 24.9236
R22438 DOUT[1].n0 DOUT[1].t2 24.9236
R22439 DOUT[1].n2 DOUT[1] 15.6165
R22440 DOUT[1] DOUT[1].n4 12.0152
R22441 DOUT[1].n1 DOUT[1] 10.4965
R22442 DOUT[1].n4 DOUT[1] 1.7925
R22443 DOUT[1].n2 DOUT[1] 1.7925
R22444 a_9575_11293.n0 a_9575_11293.t1 1327.82
R22445 a_9575_11293.t0 a_9575_11293.n0 194.655
R22446 a_9575_11293.n0 a_9575_11293.t2 63.3219
R22447 a_7367_4765.n0 a_7367_4765.t1 1327.82
R22448 a_7367_4765.n0 a_7367_4765.t2 194.655
R22449 a_7367_4765.t0 a_7367_4765.n0 63.3219
R22450 a_3017_6397.t0 a_3017_6397.t1 60.0005
R22451 a_7539_10927.t0 a_7539_10927.t1 198.571
R22452 a_7705_10927.t0 a_7705_10927.t1 60.0005
R22453 a_4857_4399.t0 a_4857_4399.t1 60.0005
R22454 COMP_P.n1 COMP_P.t5 235.763
R22455 COMP_P.n5 COMP_P.t3 221.72
R22456 COMP_P.n2 COMP_P.t4 221.72
R22457 COMP_P.n1 COMP_P.t2 163.464
R22458 COMP_P.n1 COMP_P.n0 152
R22459 COMP_P.n7 COMP_P.n6 152
R22460 COMP_P.n4 COMP_P.n3 152
R22461 COMP_P.n5 COMP_P.t0 149.421
R22462 COMP_P.n2 COMP_P.t1 149.421
R22463 COMP_P.n4 COMP_P.n2 58.019
R22464 COMP_P.n6 COMP_P.n5 43.7375
R22465 COMP_P.n0 COMP_P 22.2533
R22466 COMP_P COMP_P.n7 20.8005
R22467 COMP_P.n6 COMP_P.n1 17.8524
R22468 COMP_P.n5 COMP_P.n4 16.9598
R22469 COMP_P.n3 COMP_P 16.3205
R22470 COMP_P.n3 COMP_P 13.1205
R22471 COMP_P.n7 COMP_P 8.6405
R22472 COMP_P COMP_P.n0 0.9605
R22473 a_2071_8449.n1 a_2071_8449.t7 530.01
R22474 a_2071_8449.t0 a_2071_8449.n5 421.021
R22475 a_2071_8449.n0 a_2071_8449.t3 337.171
R22476 a_2071_8449.n3 a_2071_8449.t1 280.223
R22477 a_2071_8449.n4 a_2071_8449.t6 263.173
R22478 a_2071_8449.n4 a_2071_8449.t2 227.826
R22479 a_2071_8449.n0 a_2071_8449.t4 199.762
R22480 a_2071_8449.n2 a_2071_8449.n1 170.81
R22481 a_2071_8449.n2 a_2071_8449.n0 167.321
R22482 a_2071_8449.n5 a_2071_8449.n4 152
R22483 a_2071_8449.n1 a_2071_8449.t5 141.923
R22484 a_2071_8449.n3 a_2071_8449.n2 10.8376
R22485 a_2071_8449.n5 a_2071_8449.n3 2.50485
R22486 a_10219_3677.t0 a_10219_3677.n0 1327.82
R22487 a_10219_3677.n0 a_10219_3677.t2 194.655
R22488 a_10219_3677.n0 a_10219_3677.t1 63.3219
R22489 a_9209_7125.t0 a_9209_7125.n3 370.026
R22490 a_9209_7125.n0 a_9209_7125.t4 351.356
R22491 a_9209_7125.n1 a_9209_7125.t2 334.717
R22492 a_9209_7125.n3 a_9209_7125.t1 325.971
R22493 a_9209_7125.n1 a_9209_7125.t3 309.935
R22494 a_9209_7125.n0 a_9209_7125.t5 305.683
R22495 a_9209_7125.n2 a_9209_7125.n0 16.879
R22496 a_9209_7125.n3 a_9209_7125.n2 10.8867
R22497 a_9209_7125.n2 a_9209_7125.n1 9.3005
R22498 a_4312_12015.n1 a_4312_12015.n0 926.024
R22499 a_4312_12015.t1 a_4312_12015.n1 82.0838
R22500 a_4312_12015.n0 a_4312_12015.t0 63.3338
R22501 a_4312_12015.n1 a_4312_12015.t2 63.3219
R22502 a_4312_12015.n0 a_4312_12015.t3 29.7268
R22503 a_4135_10357.n5 a_4135_10357.n4 807.871
R22504 a_4135_10357.n0 a_4135_10357.t7 389.183
R22505 a_4135_10357.n1 a_4135_10357.n0 251.167
R22506 a_4135_10357.n1 a_4135_10357.t1 223.571
R22507 a_4135_10357.n3 a_4135_10357.t4 212.081
R22508 a_4135_10357.n2 a_4135_10357.t3 212.081
R22509 a_4135_10357.n4 a_4135_10357.n3 176.576
R22510 a_4135_10357.n0 a_4135_10357.t6 174.891
R22511 a_4135_10357.n3 a_4135_10357.t8 139.78
R22512 a_4135_10357.n2 a_4135_10357.t5 139.78
R22513 a_4135_10357.n5 a_4135_10357.t2 63.3219
R22514 a_4135_10357.t0 a_4135_10357.n5 63.3219
R22515 a_4135_10357.n3 a_4135_10357.n2 61.346
R22516 a_4135_10357.n4 a_4135_10357.n1 37.5061
R22517 x2/net7.n3 x2/net7.n2 585
R22518 x2/net7.n4 x2/net7.n3 585
R22519 x2/net7.n5 x2/net7.t5 332.312
R22520 x2/net7.n5 x2/net7.t4 295.627
R22521 x2/net7 x2/net7.n5 196.004
R22522 x2/net7.n1 x2/net7.n0 185
R22523 x2/net7 x2/net7.n1 57.7379
R22524 x2/net7.n3 x2/net7.t0 26.5955
R22525 x2/net7.n3 x2/net7.t1 26.5955
R22526 x2/net7.n0 x2/net7.t2 24.9236
R22527 x2/net7.n0 x2/net7.t3 24.9236
R22528 x2/net7.n6 x2/net7 22.6647
R22529 x2/net7.n2 x2/net7 10.4965
R22530 x2/net7.n4 x2/net7 10.4965
R22531 x2/net7.n2 x2/net7 6.9125
R22532 x2/net7 x2/net7.n6 4.3525
R22533 x2/net7.n6 x2/net7.n4 2.5605
R22534 x2/net7.n1 x2/net7 1.7925
R22535 a_4734_8029.n3 a_4734_8029.n2 647.119
R22536 a_4734_8029.n1 a_4734_8029.t5 350.253
R22537 a_4734_8029.n2 a_4734_8029.n0 260.339
R22538 a_4734_8029.n2 a_4734_8029.n1 246.119
R22539 a_4734_8029.n1 a_4734_8029.t4 189.588
R22540 a_4734_8029.n3 a_4734_8029.t1 89.1195
R22541 a_4734_8029.n0 a_4734_8029.t3 63.3338
R22542 a_4734_8029.t0 a_4734_8029.n3 41.0422
R22543 a_4734_8029.n0 a_4734_8029.t2 31.9797
R22544 a_10492_9839.n3 a_10492_9839.n2 636.953
R22545 a_10492_9839.n1 a_10492_9839.t5 366.856
R22546 a_10492_9839.n2 a_10492_9839.n0 300.2
R22547 a_10492_9839.n2 a_10492_9839.n1 225.036
R22548 a_10492_9839.n1 a_10492_9839.t4 174.056
R22549 a_10492_9839.n0 a_10492_9839.t2 70.0005
R22550 a_10492_9839.t1 a_10492_9839.n3 68.0124
R22551 a_10492_9839.n3 a_10492_9839.t3 63.3219
R22552 a_10492_9839.n0 a_10492_9839.t0 61.6672
R22553 a_2216_5059.t0 a_2216_5059.n3 370.026
R22554 a_2216_5059.n0 a_2216_5059.t5 351.356
R22555 a_2216_5059.n1 a_2216_5059.t4 334.717
R22556 a_2216_5059.n3 a_2216_5059.t1 325.971
R22557 a_2216_5059.n1 a_2216_5059.t3 309.935
R22558 a_2216_5059.n0 a_2216_5059.t2 305.683
R22559 a_2216_5059.n2 a_2216_5059.n0 16.879
R22560 a_2216_5059.n3 a_2216_5059.n2 10.8867
R22561 a_2216_5059.n2 a_2216_5059.n1 9.3005
R22562 a_2172_4943.t0 a_2172_4943.t1 126.644
R22563 a_1938_5075.n3 a_1938_5075.n2 636.953
R22564 a_1938_5075.n1 a_1938_5075.t5 366.856
R22565 a_1938_5075.n2 a_1938_5075.n0 300.2
R22566 a_1938_5075.n2 a_1938_5075.n1 225.036
R22567 a_1938_5075.n1 a_1938_5075.t4 174.056
R22568 a_1938_5075.n0 a_1938_5075.t2 70.0005
R22569 a_1938_5075.t0 a_1938_5075.n3 68.0124
R22570 a_1938_5075.n3 a_1938_5075.t3 63.3219
R22571 a_1938_5075.n0 a_1938_5075.t1 61.6672
R22572 a_2924_6031.n0 a_2924_6031.t1 1327.82
R22573 a_2924_6031.n0 a_2924_6031.t2 194.655
R22574 a_2924_6031.t0 a_2924_6031.n0 63.3219
R22575 a_10237_3829.n3 a_10237_3829.n2 647.119
R22576 a_10237_3829.n1 a_10237_3829.t5 350.253
R22577 a_10237_3829.n2 a_10237_3829.n0 260.339
R22578 a_10237_3829.n2 a_10237_3829.n1 246.119
R22579 a_10237_3829.n1 a_10237_3829.t4 189.588
R22580 a_10237_3829.n3 a_10237_3829.t0 89.1195
R22581 a_10237_3829.n0 a_10237_3829.t3 63.3338
R22582 a_10237_3829.t1 a_10237_3829.n3 41.0422
R22583 a_10237_3829.n0 a_10237_3829.t2 31.9797
R22584 a_4605_7663.n0 a_4605_7663.t1 68.3338
R22585 a_4605_7663.n0 a_4605_7663.t0 26.3935
R22586 a_4605_7663.n1 a_4605_7663.n0 14.4005
R22587 a_3386_10383.t0 a_3386_10383.t1 126.644
R22588 a_9503_6037.n1 a_9503_6037.t4 530.01
R22589 a_9503_6037.t0 a_9503_6037.n5 421.021
R22590 a_9503_6037.n0 a_9503_6037.t6 337.142
R22591 a_9503_6037.n3 a_9503_6037.t1 280.223
R22592 a_9503_6037.n4 a_9503_6037.t7 263.173
R22593 a_9503_6037.n4 a_9503_6037.t3 227.826
R22594 a_9503_6037.n0 a_9503_6037.t5 199.762
R22595 a_9503_6037.n2 a_9503_6037.n1 170.81
R22596 a_9503_6037.n2 a_9503_6037.n0 167.321
R22597 a_9503_6037.n5 a_9503_6037.n4 152
R22598 a_9503_6037.n1 a_9503_6037.t2 141.923
R22599 a_9503_6037.n3 a_9503_6037.n2 10.8376
R22600 a_9503_6037.n5 a_9503_6037.n3 2.50485
R22601 a_9924_6397.n1 a_9924_6397.n0 926.024
R22602 a_9924_6397.n1 a_9924_6397.t2 82.0838
R22603 a_9924_6397.n0 a_9924_6397.t3 63.3338
R22604 a_9924_6397.t0 a_9924_6397.n1 63.3219
R22605 a_9924_6397.n0 a_9924_6397.t1 29.7268
R22606 a_9411_9301.n1 a_9411_9301.t6 530.01
R22607 a_9411_9301.t0 a_9411_9301.n5 421.021
R22608 a_9411_9301.n0 a_9411_9301.t7 337.142
R22609 a_9411_9301.n3 a_9411_9301.t1 280.223
R22610 a_9411_9301.n4 a_9411_9301.t2 263.173
R22611 a_9411_9301.n4 a_9411_9301.t4 227.826
R22612 a_9411_9301.n0 a_9411_9301.t3 199.762
R22613 a_9411_9301.n2 a_9411_9301.n1 170.81
R22614 a_9411_9301.n2 a_9411_9301.n0 167.321
R22615 a_9411_9301.n5 a_9411_9301.n4 152
R22616 a_9411_9301.n1 a_9411_9301.t5 141.923
R22617 a_9411_9301.n3 a_9411_9301.n2 10.8376
R22618 a_9411_9301.n5 a_9411_9301.n3 2.50485
R22619 a_9577_9301.t0 a_9577_9301.n3 370.026
R22620 a_9577_9301.n0 a_9577_9301.t4 351.356
R22621 a_9577_9301.n1 a_9577_9301.t2 334.717
R22622 a_9577_9301.n3 a_9577_9301.t1 325.971
R22623 a_9577_9301.n1 a_9577_9301.t3 309.935
R22624 a_9577_9301.n0 a_9577_9301.t5 305.683
R22625 a_9577_9301.n2 a_9577_9301.n0 16.879
R22626 a_9577_9301.n3 a_9577_9301.n2 10.8867
R22627 a_9577_9301.n2 a_9577_9301.n1 9.3005
R22628 a_6813_6575.n0 a_6813_6575.t1 68.3338
R22629 a_6813_6575.n0 a_6813_6575.t0 26.3935
R22630 a_6813_6575.n1 a_6813_6575.n0 14.4005
R22631 a_8362_3311.t0 a_8362_3311.t1 87.1434
R22632 a_3018_11293.t0 a_3018_11293.t1 126.644
R22633 a_2227_8181.n3 a_2227_8181.n2 674.338
R22634 a_2227_8181.n1 a_2227_8181.t5 332.58
R22635 a_2227_8181.n2 a_2227_8181.n0 284.012
R22636 a_2227_8181.n2 a_2227_8181.n1 253.648
R22637 a_2227_8181.n1 a_2227_8181.t4 168.701
R22638 a_2227_8181.n3 a_2227_8181.t3 96.1553
R22639 a_2227_8181.t0 a_2227_8181.n3 65.6672
R22640 a_2227_8181.n0 a_2227_8181.t2 65.0005
R22641 a_2227_8181.n0 a_2227_8181.t1 45.0005
R22642 a_2526_8029.n3 a_2526_8029.n2 647.119
R22643 a_2526_8029.n1 a_2526_8029.t5 350.253
R22644 a_2526_8029.n2 a_2526_8029.n0 260.339
R22645 a_2526_8029.n2 a_2526_8029.n1 246.119
R22646 a_2526_8029.n1 a_2526_8029.t4 189.588
R22647 a_2526_8029.n3 a_2526_8029.t0 89.1195
R22648 a_2526_8029.n0 a_2526_8029.t3 63.3338
R22649 a_2526_8029.t1 a_2526_8029.n3 41.0422
R22650 a_2526_8029.n0 a_2526_8029.t2 31.9797
R22651 a_7456_8585.n3 a_7456_8585.n2 636.953
R22652 a_7456_8585.n1 a_7456_8585.t5 366.856
R22653 a_7456_8585.n2 a_7456_8585.n0 300.2
R22654 a_7456_8585.n2 a_7456_8585.n1 225.036
R22655 a_7456_8585.n1 a_7456_8585.t4 174.056
R22656 a_7456_8585.n0 a_7456_8585.t3 70.0005
R22657 a_7456_8585.t1 a_7456_8585.n3 68.0124
R22658 a_7456_8585.n3 a_7456_8585.t2 63.3219
R22659 a_7456_8585.n0 a_7456_8585.t0 61.6672
R22660 a_7937_3829.n3 a_7937_3829.n2 647.119
R22661 a_7937_3829.n1 a_7937_3829.t5 350.253
R22662 a_7937_3829.n2 a_7937_3829.n0 260.339
R22663 a_7937_3829.n2 a_7937_3829.n1 246.119
R22664 a_7937_3829.n1 a_7937_3829.t4 189.588
R22665 a_7937_3829.n3 a_7937_3829.t1 89.1195
R22666 a_7937_3829.n0 a_7937_3829.t0 63.3338
R22667 a_7937_3829.t3 a_7937_3829.n3 41.0422
R22668 a_7937_3829.n0 a_7937_3829.t2 31.9797
R22669 a_10032_10927.n3 a_10032_10927.n2 636.953
R22670 a_10032_10927.n1 a_10032_10927.t5 366.856
R22671 a_10032_10927.n2 a_10032_10927.n0 300.2
R22672 a_10032_10927.n2 a_10032_10927.n1 225.036
R22673 a_10032_10927.n1 a_10032_10927.t4 174.056
R22674 a_10032_10927.n0 a_10032_10927.t2 70.0005
R22675 a_10032_10927.t1 a_10032_10927.n3 68.0124
R22676 a_10032_10927.n3 a_10032_10927.t3 63.3219
R22677 a_10032_10927.n0 a_10032_10927.t0 61.6672
R22678 a_2387_10927.t1 a_2387_10927.t0 198.571
R22679 a_2553_10927.t0 a_2553_10927.t1 60.0005
R22680 a_6633_11477.t0 a_6633_11477.n3 370.026
R22681 a_6633_11477.n0 a_6633_11477.t2 351.356
R22682 a_6633_11477.n1 a_6633_11477.t4 334.717
R22683 a_6633_11477.n3 a_6633_11477.t1 325.971
R22684 a_6633_11477.n1 a_6633_11477.t5 309.935
R22685 a_6633_11477.n0 a_6633_11477.t3 305.683
R22686 a_6633_11477.n2 a_6633_11477.n0 16.879
R22687 a_6633_11477.n3 a_6633_11477.n2 10.8867
R22688 a_6633_11477.n2 a_6633_11477.n1 9.3005
R22689 a_7201_11445.n3 a_7201_11445.n2 647.119
R22690 a_7201_11445.n1 a_7201_11445.t5 350.253
R22691 a_7201_11445.n2 a_7201_11445.n0 260.339
R22692 a_7201_11445.n2 a_7201_11445.n1 246.119
R22693 a_7201_11445.n1 a_7201_11445.t4 189.588
R22694 a_7201_11445.n3 a_7201_11445.t3 89.1195
R22695 a_7201_11445.n0 a_7201_11445.t2 63.3338
R22696 a_7201_11445.t0 a_7201_11445.n3 41.0422
R22697 a_7201_11445.n0 a_7201_11445.t1 31.9797
R22698 a_4288_8207.t0 a_4288_8207.t1 126.644
R22699 a_4837_8573.t0 a_4837_8573.t1 198.571
R22700 a_5620_3579.t0 a_5620_3579.n3 370.026
R22701 a_5620_3579.n0 a_5620_3579.t5 351.356
R22702 a_5620_3579.n1 a_5620_3579.t2 334.717
R22703 a_5620_3579.n3 a_5620_3579.t1 325.971
R22704 a_5620_3579.n1 a_5620_3579.t4 309.935
R22705 a_5620_3579.n0 a_5620_3579.t3 305.683
R22706 a_5620_3579.n2 a_5620_3579.n0 16.879
R22707 a_5620_3579.n3 a_5620_3579.n2 10.8867
R22708 a_5620_3579.n2 a_5620_3579.n1 9.3005
R22709 a_6125_3311.t0 a_6125_3311.t1 198.571
R22710 a_5815_3548.n3 a_5815_3548.n2 674.338
R22711 a_5815_3548.n1 a_5815_3548.t4 332.58
R22712 a_5815_3548.n2 a_5815_3548.n0 284.012
R22713 a_5815_3548.n2 a_5815_3548.n1 253.648
R22714 a_5815_3548.n1 a_5815_3548.t5 168.701
R22715 a_5815_3548.t0 a_5815_3548.n3 96.1553
R22716 a_5815_3548.n3 a_5815_3548.t3 65.6672
R22717 a_5815_3548.n0 a_5815_3548.t1 65.0005
R22718 a_5815_3548.n0 a_5815_3548.t2 45.0005
R22719 a_5366_8029.n1 a_5366_8029.n0 926.024
R22720 a_5366_8029.t1 a_5366_8029.n1 82.0838
R22721 a_5366_8029.n0 a_5366_8029.t0 63.3338
R22722 a_5366_8029.n1 a_5366_8029.t2 63.3219
R22723 a_5366_8029.n0 a_5366_8029.t3 29.7268
R22724 a_7723_11775.n5 a_7723_11775.n4 807.871
R22725 a_7723_11775.n2 a_7723_11775.t5 389.183
R22726 a_7723_11775.n3 a_7723_11775.n2 251.167
R22727 a_7723_11775.n3 a_7723_11775.t1 223.571
R22728 a_7723_11775.n0 a_7723_11775.t7 212.081
R22729 a_7723_11775.n1 a_7723_11775.t6 212.081
R22730 a_7723_11775.n4 a_7723_11775.n1 176.576
R22731 a_7723_11775.n2 a_7723_11775.t8 174.891
R22732 a_7723_11775.n0 a_7723_11775.t4 139.78
R22733 a_7723_11775.n1 a_7723_11775.t3 139.78
R22734 a_7723_11775.n5 a_7723_11775.t2 63.3219
R22735 a_7723_11775.t0 a_7723_11775.n5 63.3219
R22736 a_7723_11775.n1 a_7723_11775.n0 61.346
R22737 a_7723_11775.n4 a_7723_11775.n3 37.7195
R22738 a_5161_10927.t0 a_5161_10927.n3 370.026
R22739 a_5161_10927.n0 a_5161_10927.t2 351.356
R22740 a_5161_10927.n1 a_5161_10927.t3 334.717
R22741 a_5161_10927.n3 a_5161_10927.t1 325.971
R22742 a_5161_10927.n1 a_5161_10927.t5 309.935
R22743 a_5161_10927.n0 a_5161_10927.t4 305.683
R22744 a_5161_10927.n2 a_5161_10927.n0 16.879
R22745 a_5161_10927.n3 a_5161_10927.n2 10.8867
R22746 a_5161_10927.n2 a_5161_10927.n1 9.3005
R22747 a_5617_3311.n0 a_5617_3311.t0 68.3338
R22748 a_5617_3311.n0 a_5617_3311.t1 26.3935
R22749 a_5617_3311.n1 a_5617_3311.n0 14.4005
R22750 a_2540_6031.t0 a_2540_6031.t1 126.644
R22751 a_8454_6397.t0 a_8454_6397.t1 87.1434
R22752 a_6431_7663.n3 a_6431_7663.n2 674.338
R22753 a_6431_7663.n1 a_6431_7663.t5 332.58
R22754 a_6431_7663.n2 a_6431_7663.n0 284.012
R22755 a_6431_7663.n2 a_6431_7663.n1 253.648
R22756 a_6431_7663.n1 a_6431_7663.t4 168.701
R22757 a_6431_7663.t1 a_6431_7663.n3 96.1553
R22758 a_6431_7663.n3 a_6431_7663.t3 65.6672
R22759 a_6431_7663.n0 a_6431_7663.t0 65.0005
R22760 a_6431_7663.n0 a_6431_7663.t2 45.0005
R22761 a_6539_8029.n0 a_6539_8029.t2 1327.82
R22762 a_6539_8029.t0 a_6539_8029.n0 194.655
R22763 a_6539_8029.n0 a_6539_8029.t1 63.3219
R22764 a_10145_10081.n3 a_10145_10081.n2 647.119
R22765 a_10145_10081.n1 a_10145_10081.t5 350.253
R22766 a_10145_10081.n2 a_10145_10081.n0 260.339
R22767 a_10145_10081.n2 a_10145_10081.n1 246.119
R22768 a_10145_10081.n1 a_10145_10081.t4 189.588
R22769 a_10145_10081.n3 a_10145_10081.t0 89.1195
R22770 a_10145_10081.n0 a_10145_10081.t1 63.3338
R22771 a_10145_10081.t2 a_10145_10081.n3 41.0422
R22772 a_10145_10081.n0 a_10145_10081.t3 31.9797
R22773 a_4422_10515.n3 a_4422_10515.n2 636.953
R22774 a_4422_10515.n1 a_4422_10515.t5 366.856
R22775 a_4422_10515.n2 a_4422_10515.n0 300.2
R22776 a_4422_10515.n2 a_4422_10515.n1 225.036
R22777 a_4422_10515.n1 a_4422_10515.t4 174.056
R22778 a_4422_10515.n0 a_4422_10515.t2 70.0005
R22779 a_4422_10515.t0 a_4422_10515.n3 68.0124
R22780 a_4422_10515.n3 a_4422_10515.t3 63.3219
R22781 a_4422_10515.n0 a_4422_10515.t1 61.6672
R22782 a_3870_5075.n3 a_3870_5075.n2 636.953
R22783 a_3870_5075.n1 a_3870_5075.t4 366.856
R22784 a_3870_5075.n2 a_3870_5075.n0 300.2
R22785 a_3870_5075.n2 a_3870_5075.n1 225.036
R22786 a_3870_5075.n1 a_3870_5075.t5 174.056
R22787 a_3870_5075.n0 a_3870_5075.t3 70.0005
R22788 a_3870_5075.t1 a_3870_5075.n3 68.0124
R22789 a_3870_5075.n3 a_3870_5075.t2 63.3219
R22790 a_3870_5075.n0 a_3870_5075.t0 61.6672
R22791 a_4973_6397.t0 a_4973_6397.t1 94.7268
R22792 a_2356_4765.t0 a_2356_4765.t1 126.644
R22793 a_2122_4651.n3 a_2122_4651.n2 636.953
R22794 a_2122_4651.n1 a_2122_4651.t5 366.856
R22795 a_2122_4651.n2 a_2122_4651.n0 300.2
R22796 a_2122_4651.n2 a_2122_4651.n1 225.036
R22797 a_2122_4651.n1 a_2122_4651.t4 174.056
R22798 a_2122_4651.n0 a_2122_4651.t0 70.0005
R22799 a_2122_4651.n3 a_2122_4651.t2 68.0124
R22800 a_2122_4651.t1 a_2122_4651.n3 63.3219
R22801 a_2122_4651.n0 a_2122_4651.t3 61.6672
R22802 a_10785_5487.t1 a_10785_5487.t0 94.7268
R22803 a_9832_9839.n1 a_9832_9839.n0 926.024
R22804 a_9832_9839.n0 a_9832_9839.t3 82.0838
R22805 a_9832_9839.n1 a_9832_9839.t2 63.3338
R22806 a_9832_9839.n0 a_9832_9839.t1 63.3219
R22807 a_9832_9839.n2 a_9832_9839.t0 26.3935
R22808 a_9832_9839.n3 a_9832_9839.n2 14.4005
R22809 a_9832_9839.n2 a_9832_9839.n1 3.33383
R22810 a_10584_3145.n3 a_10584_3145.n2 636.953
R22811 a_10584_3145.n1 a_10584_3145.t4 366.856
R22812 a_10584_3145.n2 a_10584_3145.n0 300.2
R22813 a_10584_3145.n2 a_10584_3145.n1 225.036
R22814 a_10584_3145.n1 a_10584_3145.t5 174.056
R22815 a_10584_3145.n0 a_10584_3145.t0 70.0005
R22816 a_10584_3145.n3 a_10584_3145.t3 68.0124
R22817 a_10584_3145.t1 a_10584_3145.n3 63.3219
R22818 a_10584_3145.n0 a_10584_3145.t2 61.6672
R22819 a_10693_3145.n0 a_10693_3145.t1 68.3338
R22820 a_10693_3145.n0 a_10693_3145.t0 26.3935
R22821 a_10693_3145.n1 a_10693_3145.n0 14.4005
R22822 a_8170_3677.t0 a_8170_3677.t1 126.644
R22823 a_3224_10761.n3 a_3224_10761.n2 636.953
R22824 a_3224_10761.n1 a_3224_10761.t5 366.856
R22825 a_3224_10761.n2 a_3224_10761.n0 300.2
R22826 a_3224_10761.n2 a_3224_10761.n1 225.036
R22827 a_3224_10761.n1 a_3224_10761.t4 174.056
R22828 a_3224_10761.n0 a_3224_10761.t2 70.0005
R22829 a_3224_10761.t0 a_3224_10761.n3 68.0124
R22830 a_3224_10761.n3 a_3224_10761.t3 63.3219
R22831 a_3224_10761.n0 a_3224_10761.t1 61.6672
R22832 a_3333_10761.n0 a_3333_10761.t0 68.3338
R22833 a_3333_10761.n0 a_3333_10761.t1 26.3935
R22834 a_3333_10761.n1 a_3333_10761.n0 14.4005
R22835 CLKSB.n0 CLKSB.t0 235.56
R22836 CLKSB.n2 CLKSB.t1 130.594
R22837 CLKSB CLKSB.n2 22.2966
R22838 CLKSB.n2 CLKSB.n1 13.7066
R22839 CLKSB.n1 CLKSB 4.55579
R22840 CLKSB CLKSB.n0 2.22659
R22841 CLKSB.n0 CLKSB 1.55202
R22842 a_9117_10927.t0 a_9117_10927.n3 370.026
R22843 a_9117_10927.n0 a_9117_10927.t3 351.356
R22844 a_9117_10927.n1 a_9117_10927.t5 334.717
R22845 a_9117_10927.n3 a_9117_10927.t1 325.971
R22846 a_9117_10927.n1 a_9117_10927.t2 309.935
R22847 a_9117_10927.n0 a_9117_10927.t4 305.683
R22848 a_9117_10927.n2 a_9117_10927.n0 16.879
R22849 a_9117_10927.n3 a_9117_10927.n2 10.8867
R22850 a_9117_10927.n2 a_9117_10927.n1 9.3005
R22851 x2/net2.n5 x2/net2.n4 585
R22852 x2/net2.n6 x2/net2.n5 585
R22853 x2/net2.n2 x2/net2.t5 333.651
R22854 x2/net2.n2 x2/net2.t4 297.233
R22855 x2/net2.n3 x2/net2.n2 195.701
R22856 x2/net2.n1 x2/net2.n0 185
R22857 x2/net2 x2/net2.n1 49.0339
R22858 x2/net2.n5 x2/net2.t1 26.5955
R22859 x2/net2.n5 x2/net2.t0 26.5955
R22860 x2/net2.n0 x2/net2.t3 24.9236
R22861 x2/net2.n0 x2/net2.t2 24.9236
R22862 x2/net2.n4 x2/net2 17.0535
R22863 x2/net2.n6 x2/net2 15.6165
R22864 x2/net2 x2/net2.n3 14.4935
R22865 x2/net2.n1 x2/net2 10.4965
R22866 x2/net2.n4 x2/net2 1.7925
R22867 x2/net2 x2/net2.n6 1.7925
R22868 x2/net2.n3 x2/net2 1.03669
R22869 a_10219_5853.n0 a_10219_5853.t1 1327.82
R22870 a_10219_5853.n0 a_10219_5853.t2 194.655
R22871 a_10219_5853.t0 a_10219_5853.n0 63.3219
R22872 a_4976_11587.t0 a_4976_11587.n3 370.026
R22873 a_4976_11587.n0 a_4976_11587.t4 351.356
R22874 a_4976_11587.n1 a_4976_11587.t3 334.717
R22875 a_4976_11587.n3 a_4976_11587.t1 325.971
R22876 a_4976_11587.n1 a_4976_11587.t5 309.935
R22877 a_4976_11587.n0 a_4976_11587.t2 305.683
R22878 a_4976_11587.n2 a_4976_11587.n0 16.879
R22879 a_4976_11587.n3 a_4976_11587.n2 10.8867
R22880 a_4976_11587.n2 a_4976_11587.n1 9.3005
R22881 a_4932_11471.t0 a_4932_11471.t1 126.644
R22882 a_4698_11603.n3 a_4698_11603.n2 636.953
R22883 a_4698_11603.n1 a_4698_11603.t4 366.856
R22884 a_4698_11603.n2 a_4698_11603.n0 300.2
R22885 a_4698_11603.n2 a_4698_11603.n1 225.036
R22886 a_4698_11603.n1 a_4698_11603.t5 174.056
R22887 a_4698_11603.n0 a_4698_11603.t0 70.0005
R22888 a_4698_11603.n3 a_4698_11603.t2 68.0124
R22889 a_4698_11603.t1 a_4698_11603.n3 63.3219
R22890 a_4698_11603.n0 a_4698_11603.t3 61.6672
R22891 SWP[1].n0 SWP[1].t4 333.651
R22892 SWP[1].n0 SWP[1].t5 297.233
R22893 SWP[1].n2 SWP[1].n1 289.096
R22894 SWP[1] SWP[1].n0 194.062
R22895 SWP[1].n4 SWP[1].n3 185
R22896 SWP[1] SWP[1].n6 60.323
R22897 SWP[1].n4 SWP[1] 49.0339
R22898 SWP[1].n1 SWP[1].t1 26.5955
R22899 SWP[1].n1 SWP[1].t0 26.5955
R22900 SWP[1].n3 SWP[1].t2 24.9236
R22901 SWP[1].n3 SWP[1].t3 24.9236
R22902 SWP[1].n6 SWP[1] 15.9249
R22903 SWP[1] SWP[1].n2 9.48653
R22904 SWP[1].n6 SWP[1].n5 9.3005
R22905 SWP[1].n2 SWP[1] 7.7181
R22906 SWP[1].n5 SWP[1].n4 6.1445
R22907 SWP[1].n5 SWP[1] 4.3525
R22908 a_7710_11471.t0 a_7710_11471.t1 126.644
R22909 a_5316_2767.n0 a_5316_2767.t1 1327.82
R22910 a_5316_2767.n0 a_5316_2767.t2 194.655
R22911 a_5316_2767.t0 a_5316_2767.n0 63.3219
R22912 a_2356_8029.t0 a_2356_8029.t1 126.644
R22913 a_3609_11849.n0 a_3609_11849.t0 68.3338
R22914 a_3609_11849.n0 a_3609_11849.t1 26.3935
R22915 a_3609_11849.n1 a_3609_11849.n0 14.4005
R22916 a_7093_5487.t0 a_7093_5487.n3 370.026
R22917 a_7093_5487.n0 a_7093_5487.t5 351.356
R22918 a_7093_5487.n1 a_7093_5487.t3 334.717
R22919 a_7093_5487.n3 a_7093_5487.t1 325.971
R22920 a_7093_5487.n1 a_7093_5487.t2 309.935
R22921 a_7093_5487.n0 a_7093_5487.t4 305.683
R22922 a_7093_5487.n2 a_7093_5487.n0 16.879
R22923 a_7093_5487.n3 a_7093_5487.n2 10.8867
R22924 a_7093_5487.n2 a_7093_5487.n1 9.3005
R22925 a_4698_6163.n3 a_4698_6163.n2 636.953
R22926 a_4698_6163.n1 a_4698_6163.t4 366.856
R22927 a_4698_6163.n2 a_4698_6163.n0 300.2
R22928 a_4698_6163.n2 a_4698_6163.n1 225.036
R22929 a_4698_6163.n1 a_4698_6163.t5 174.056
R22930 a_4698_6163.n0 a_4698_6163.t1 70.0005
R22931 a_4698_6163.n3 a_4698_6163.t2 68.0124
R22932 a_4698_6163.t0 a_4698_6163.n3 63.3219
R22933 a_4698_6163.n0 a_4698_6163.t3 61.6672
R22934 a_7091_11471.n0 a_7091_11471.t2 1327.82
R22935 a_7091_11471.n0 a_7091_11471.t1 194.655
R22936 a_7091_11471.t0 a_7091_11471.n0 63.3219
R22937 a_9729_10927.t0 a_9729_10927.t1 60.0005
R22938 a_10141_8751.t0 a_10141_8751.t1 94.7268
R22939 a_7551_3677.n0 a_7551_3677.t1 1327.82
R22940 a_7551_3677.n0 a_7551_3677.t2 194.655
R22941 a_7551_3677.t0 a_7551_3677.n0 63.3219
R22942 a_4976_2883.t0 a_4976_2883.n3 370.026
R22943 a_4976_2883.n0 a_4976_2883.t4 351.356
R22944 a_4976_2883.n1 a_4976_2883.t3 334.717
R22945 a_4976_2883.n3 a_4976_2883.t1 325.971
R22946 a_4976_2883.n1 a_4976_2883.t2 309.935
R22947 a_4976_2883.n0 a_4976_2883.t5 305.683
R22948 a_4976_2883.n2 a_4976_2883.n0 16.879
R22949 a_4976_2883.n3 a_4976_2883.n2 10.8867
R22950 a_4976_2883.n2 a_4976_2883.n1 9.3005
R22951 a_7801_3133.t0 a_7801_3133.t1 60.0005
R22952 a_7708_9117.t0 a_7708_9117.n0 1327.82
R22953 a_7708_9117.n0 a_7708_9117.t1 194.655
R22954 a_7708_9117.n0 a_7708_9117.t2 63.3219
R22955 a_7563_8988.n3 a_7563_8988.n2 674.338
R22956 a_7563_8988.n1 a_7563_8988.t5 332.58
R22957 a_7563_8988.n2 a_7563_8988.n0 284.012
R22958 a_7563_8988.n2 a_7563_8988.n1 253.648
R22959 a_7563_8988.n1 a_7563_8988.t4 168.701
R22960 a_7563_8988.t1 a_7563_8988.n3 96.1553
R22961 a_7563_8988.n3 a_7563_8988.t3 65.6672
R22962 a_7563_8988.n0 a_7563_8988.t0 65.0005
R22963 a_7563_8988.n0 a_7563_8988.t2 45.0005
R22964 a_5300_5853.t0 a_5300_5853.t1 126.644
R22965 a_5066_5739.n3 a_5066_5739.n2 636.953
R22966 a_5066_5739.n1 a_5066_5739.t5 366.856
R22967 a_5066_5739.n2 a_5066_5739.n0 300.2
R22968 a_5066_5739.n2 a_5066_5739.n1 225.036
R22969 a_5066_5739.n1 a_5066_5739.t4 174.056
R22970 a_5066_5739.n0 a_5066_5739.t2 70.0005
R22971 a_5066_5739.t0 a_5066_5739.n3 68.0124
R22972 a_5066_5739.n3 a_5066_5739.t3 63.3219
R22973 a_5066_5739.n0 a_5066_5739.t1 61.6672
R22974 a_10035_10205.n0 a_10035_10205.t2 1327.82
R22975 a_10035_10205.t0 a_10035_10205.n0 194.655
R22976 a_10035_10205.n0 a_10035_10205.t1 63.3219
R22977 a_3089_6397.t0 a_3089_6397.t1 198.571
R22978 a_4619_6812.n3 a_4619_6812.n2 674.338
R22979 a_4619_6812.n1 a_4619_6812.t5 332.58
R22980 a_4619_6812.n2 a_4619_6812.n0 284.012
R22981 a_4619_6812.n2 a_4619_6812.n1 253.648
R22982 a_4619_6812.n1 a_4619_6812.t4 168.701
R22983 a_4619_6812.n3 a_4619_6812.t3 96.1553
R22984 a_4619_6812.t0 a_4619_6812.n3 65.6672
R22985 a_4619_6812.n0 a_4619_6812.t2 65.0005
R22986 a_4619_6812.n0 a_4619_6812.t1 45.0005
R22987 a_6649_7905.n3 a_6649_7905.n2 647.119
R22988 a_6649_7905.n1 a_6649_7905.t4 350.253
R22989 a_6649_7905.n2 a_6649_7905.n0 260.339
R22990 a_6649_7905.n2 a_6649_7905.n1 246.119
R22991 a_6649_7905.n1 a_6649_7905.t5 189.588
R22992 a_6649_7905.n3 a_6649_7905.t0 89.1195
R22993 a_6649_7905.n0 a_6649_7905.t1 63.3338
R22994 a_6649_7905.t2 a_6649_7905.n3 41.0422
R22995 a_6649_7905.n0 a_6649_7905.t3 31.9797
R22996 a_4932_6031.t0 a_4932_6031.t1 126.644
R22997 a_9559_7497.n3 a_9559_7497.n2 674.338
R22998 a_9559_7497.n1 a_9559_7497.t4 332.58
R22999 a_9559_7497.n2 a_9559_7497.n0 284.012
R23000 a_9559_7497.n2 a_9559_7497.n1 253.648
R23001 a_9559_7497.n1 a_9559_7497.t5 168.701
R23002 a_9559_7497.t1 a_9559_7497.n3 96.1553
R23003 a_9559_7497.n3 a_9559_7497.t2 65.6672
R23004 a_9559_7497.n0 a_9559_7497.t0 65.0005
R23005 a_9559_7497.n0 a_9559_7497.t3 45.0005
R23006 a_9655_7497.t1 a_9655_7497.t0 198.571
R23007 a_5102_6031.n3 a_5102_6031.n2 647.119
R23008 a_5102_6031.n1 a_5102_6031.t4 350.253
R23009 a_5102_6031.n2 a_5102_6031.n0 260.339
R23010 a_5102_6031.n2 a_5102_6031.n1 246.119
R23011 a_5102_6031.n1 a_5102_6031.t5 189.588
R23012 a_5102_6031.n3 a_5102_6031.t1 89.1195
R23013 a_5102_6031.n0 a_5102_6031.t0 63.3338
R23014 a_5102_6031.t2 a_5102_6031.n3 41.0422
R23015 a_5102_6031.n0 a_5102_6031.t3 31.9797
R23016 a_2581_6397.t0 a_2581_6397.t1 94.7268
R23017 SWP[2].n0 SWP[2].t4 333.651
R23018 SWP[2].n0 SWP[2].t5 297.233
R23019 SWP[2].n2 SWP[2].n1 289.096
R23020 SWP[2] SWP[2].n0 194.062
R23021 SWP[2].n4 SWP[2].n3 185
R23022 SWP[2].n6 SWP[2] 59.0725
R23023 SWP[2].n4 SWP[2] 49.0339
R23024 SWP[2].n1 SWP[2].t0 26.5955
R23025 SWP[2].n1 SWP[2].t1 26.5955
R23026 SWP[2].n3 SWP[2].t3 24.9236
R23027 SWP[2].n3 SWP[2].t2 24.9236
R23028 SWP[2] SWP[2].n2 9.48653
R23029 SWP[2].n6 SWP[2].n5 9.3005
R23030 SWP[2].n2 SWP[2] 7.7181
R23031 SWP[2].n5 SWP[2].n4 6.1445
R23032 SWP[2] SWP[2].n6 5.1176
R23033 SWP[2].n5 SWP[2] 4.3525
R23034 a_6909_4399.t0 a_6909_4399.n3 370.026
R23035 a_6909_4399.n0 a_6909_4399.t3 351.356
R23036 a_6909_4399.n1 a_6909_4399.t2 334.717
R23037 a_6909_4399.n3 a_6909_4399.t1 325.971
R23038 a_6909_4399.n1 a_6909_4399.t4 309.935
R23039 a_6909_4399.n0 a_6909_4399.t5 305.683
R23040 a_6909_4399.n2 a_6909_4399.n0 16.879
R23041 a_6909_4399.n3 a_6909_4399.n2 10.8867
R23042 a_6909_4399.n2 a_6909_4399.n1 9.3005
R23043 a_7259_4399.n3 a_7259_4399.n2 674.338
R23044 a_7259_4399.n1 a_7259_4399.t4 332.58
R23045 a_7259_4399.n2 a_7259_4399.n0 284.012
R23046 a_7259_4399.n2 a_7259_4399.n1 253.648
R23047 a_7259_4399.n1 a_7259_4399.t5 168.701
R23048 a_7259_4399.t0 a_7259_4399.n3 96.1553
R23049 a_7259_4399.n3 a_7259_4399.t3 65.6672
R23050 a_7259_4399.n0 a_7259_4399.t1 65.0005
R23051 a_7259_4399.n0 a_7259_4399.t2 45.0005
R23052 a_7355_4399.t0 a_7355_4399.t1 198.571
R23053 a_2833_5487.t0 a_2833_5487.t1 60.0005
R23054 a_4411_11445.n4 a_4411_11445.n1 807.871
R23055 a_4411_11445.n0 a_4411_11445.t5 389.183
R23056 a_4411_11445.n5 a_4411_11445.n0 251.167
R23057 a_4411_11445.t0 a_4411_11445.n5 223.571
R23058 a_4411_11445.n3 a_4411_11445.t7 212.081
R23059 a_4411_11445.n2 a_4411_11445.t8 212.081
R23060 a_4411_11445.n4 a_4411_11445.n3 176.576
R23061 a_4411_11445.n0 a_4411_11445.t3 174.891
R23062 a_4411_11445.n3 a_4411_11445.t4 139.78
R23063 a_4411_11445.n2 a_4411_11445.t6 139.78
R23064 a_4411_11445.n1 a_4411_11445.t2 63.3219
R23065 a_4411_11445.n1 a_4411_11445.t1 63.3219
R23066 a_4411_11445.n3 a_4411_11445.n2 61.346
R23067 a_4411_11445.n5 a_4411_11445.n4 37.5061
R23068 a_4973_11837.t0 a_4973_11837.t1 94.7268
R23069 a_10654_9295.t0 a_10654_9295.t1 126.644
R23070 a_2974_4943.n1 a_2974_4943.n0 926.024
R23071 a_2974_4943.n1 a_2974_4943.t3 82.0838
R23072 a_2974_4943.n0 a_2974_4943.t2 63.3338
R23073 a_2974_4943.t0 a_2974_4943.n1 63.3219
R23074 a_2974_4943.n0 a_2974_4943.t1 29.7268
R23075 a_10386_7663.t0 a_10386_7663.t1 87.1434
R23076 a_9669_2773.t0 a_9669_2773.n3 370.026
R23077 a_9669_2773.n0 a_9669_2773.t2 351.356
R23078 a_9669_2773.n1 a_9669_2773.t3 334.717
R23079 a_9669_2773.n3 a_9669_2773.t1 325.971
R23080 a_9669_2773.n1 a_9669_2773.t4 309.935
R23081 a_9669_2773.n0 a_9669_2773.t5 305.683
R23082 a_9669_2773.n2 a_9669_2773.n0 16.879
R23083 a_9669_2773.n3 a_9669_2773.n2 10.8867
R23084 a_9669_2773.n2 a_9669_2773.n1 9.3005
R23085 a_10746_6031.t0 a_10746_6031.t1 126.644
R23086 a_7368_2883.t0 a_7368_2883.n3 370.026
R23087 a_7368_2883.n0 a_7368_2883.t2 351.356
R23088 a_7368_2883.n1 a_7368_2883.t3 334.717
R23089 a_7368_2883.n3 a_7368_2883.t1 325.971
R23090 a_7368_2883.n1 a_7368_2883.t4 309.935
R23091 a_7368_2883.n0 a_7368_2883.t5 305.683
R23092 a_7368_2883.n2 a_7368_2883.n0 16.879
R23093 a_7368_2883.n3 a_7368_2883.n2 10.8867
R23094 a_7368_2883.n2 a_7368_2883.n1 9.3005
R23095 a_6772_6941.t0 a_6772_6941.t1 126.644
R23096 a_10286_7119.t0 a_10286_7119.t1 126.644
R23097 a_2465_8751.t0 a_2465_8751.t1 60.0005
R23098 a_7719_4233.n3 a_7719_4233.n2 674.338
R23099 a_7719_4233.n1 a_7719_4233.t5 332.58
R23100 a_7719_4233.n2 a_7719_4233.n0 284.012
R23101 a_7719_4233.n2 a_7719_4233.n1 253.648
R23102 a_7719_4233.n1 a_7719_4233.t4 168.701
R23103 a_7719_4233.n3 a_7719_4233.t3 96.1553
R23104 a_7719_4233.t1 a_7719_4233.n3 65.6672
R23105 a_7719_4233.n0 a_7719_4233.t2 65.0005
R23106 a_7719_4233.n0 a_7719_4233.t0 45.0005
R23107 a_5694_4221.t0 a_5694_4221.t1 87.1434
R23108 a_10421_6817.n3 a_10421_6817.n2 647.119
R23109 a_10421_6817.n1 a_10421_6817.t5 350.253
R23110 a_10421_6817.n2 a_10421_6817.n0 260.339
R23111 a_10421_6817.n2 a_10421_6817.n1 246.119
R23112 a_10421_6817.n1 a_10421_6817.t4 189.588
R23113 a_10421_6817.n3 a_10421_6817.t0 89.1195
R23114 a_10421_6817.n0 a_10421_6817.t1 63.3338
R23115 a_10421_6817.t2 a_10421_6817.n3 41.0422
R23116 a_10421_6817.n0 a_10421_6817.t3 31.9797
R23117 a_5746_3677.n3 a_5746_3677.n2 647.119
R23118 a_5746_3677.n1 a_5746_3677.t5 350.253
R23119 a_5746_3677.n2 a_5746_3677.n0 260.339
R23120 a_5746_3677.n2 a_5746_3677.n1 246.119
R23121 a_5746_3677.n1 a_5746_3677.t4 189.588
R23122 a_5746_3677.n3 a_5746_3677.t0 89.1195
R23123 a_5746_3677.n0 a_5746_3677.t3 63.3338
R23124 a_5746_3677.t1 a_5746_3677.n3 41.0422
R23125 a_5746_3677.n0 a_5746_3677.t2 31.9797
R23126 a_7661_5729.n3 a_7661_5729.n2 647.119
R23127 a_7661_5729.n1 a_7661_5729.t4 350.253
R23128 a_7661_5729.n2 a_7661_5729.n0 260.339
R23129 a_7661_5729.n2 a_7661_5729.n1 246.119
R23130 a_7661_5729.n1 a_7661_5729.t5 189.588
R23131 a_7661_5729.n3 a_7661_5729.t3 89.1195
R23132 a_7661_5729.n0 a_7661_5729.t0 63.3338
R23133 a_7661_5729.t1 a_7661_5729.n3 41.0422
R23134 a_7661_5729.n0 a_7661_5729.t2 31.9797
R23135 a_7539_5487.t1 a_7539_5487.t0 198.571
R23136 a_7705_5487.t0 a_7705_5487.t1 60.0005
R23137 a_10145_9269.n3 a_10145_9269.n2 647.119
R23138 a_10145_9269.n1 a_10145_9269.t5 350.253
R23139 a_10145_9269.n2 a_10145_9269.n0 260.339
R23140 a_10145_9269.n2 a_10145_9269.n1 246.119
R23141 a_10145_9269.n1 a_10145_9269.t4 189.588
R23142 a_10145_9269.n3 a_10145_9269.t0 89.1195
R23143 a_10145_9269.n0 a_10145_9269.t1 63.3338
R23144 a_10145_9269.t3 a_10145_9269.n3 41.0422
R23145 a_10145_9269.n0 a_10145_9269.t2 31.9797
R23146 a_10035_9295.n0 a_10035_9295.t2 1327.82
R23147 a_10035_9295.t0 a_10035_9295.n0 194.655
R23148 a_10035_9295.n0 a_10035_9295.t1 63.3219
R23149 a_7618_8207.t0 a_7618_8207.t1 126.644
R23150 a_5134_12381.t0 a_5134_12381.t1 126.644
R23151 a_8339_6603.n2 a_8339_6603.n1 672.948
R23152 a_8339_6603.n1 a_8339_6603.t1 314.563
R23153 a_8339_6603.n0 a_8339_6603.t3 236.18
R23154 a_8339_6603.n0 a_8339_6603.t4 163.881
R23155 a_8339_6603.n1 a_8339_6603.n0 152
R23156 a_8339_6603.t0 a_8339_6603.n2 63.3219
R23157 a_8339_6603.n2 a_8339_6603.t2 63.3219
R23158 a_4380_9117.t0 a_4380_9117.t1 126.644
R23159 a_2556_4943.n0 a_2556_4943.t2 1327.82
R23160 a_2556_4943.n0 a_2556_4943.t1 194.655
R23161 a_2556_4943.t0 a_2556_4943.n0 63.3219
R23162 a_9464_7485.n1 a_9464_7485.n0 926.024
R23163 a_9464_7485.t1 a_9464_7485.n1 82.0838
R23164 a_9464_7485.n0 a_9464_7485.t0 63.3338
R23165 a_9464_7485.n1 a_9464_7485.t2 63.3219
R23166 a_9464_7485.n0 a_9464_7485.t3 29.7268
R23167 a_2595_4636.n3 a_2595_4636.n2 674.338
R23168 a_2595_4636.n1 a_2595_4636.t5 332.58
R23169 a_2595_4636.n2 a_2595_4636.n0 284.012
R23170 a_2595_4636.n2 a_2595_4636.n1 253.648
R23171 a_2595_4636.n1 a_2595_4636.t4 168.701
R23172 a_2595_4636.n3 a_2595_4636.t2 96.1553
R23173 a_2595_4636.t1 a_2595_4636.n3 65.6672
R23174 a_2595_4636.n0 a_2595_4636.t3 65.0005
R23175 a_2595_4636.n0 a_2595_4636.t0 45.0005
R23176 a_3158_4765.n1 a_3158_4765.n0 926.024
R23177 a_3158_4765.t0 a_3158_4765.n1 82.0838
R23178 a_3158_4765.n0 a_3158_4765.t3 63.3338
R23179 a_3158_4765.n1 a_3158_4765.t1 63.3219
R23180 a_3158_4765.n0 a_3158_4765.t2 29.7268
R23181 a_2158_9117.n3 a_2158_9117.n2 647.119
R23182 a_2158_9117.n1 a_2158_9117.t5 350.253
R23183 a_2158_9117.n2 a_2158_9117.n0 260.339
R23184 a_2158_9117.n2 a_2158_9117.n1 246.119
R23185 a_2158_9117.n1 a_2158_9117.t4 189.588
R23186 a_2158_9117.n3 a_2158_9117.t1 89.1195
R23187 a_2158_9117.n0 a_2158_9117.t0 63.3338
R23188 a_2158_9117.t2 a_2158_9117.n3 41.0422
R23189 a_2158_9117.n0 a_2158_9117.t3 31.9797
R23190 a_2372_9117.n0 a_2372_9117.t2 1327.82
R23191 a_2372_9117.t0 a_2372_9117.n0 194.655
R23192 a_2372_9117.n0 a_2372_9117.t1 63.3219
R23193 a_7873_3133.t0 a_7873_3133.t1 198.571
R23194 a_3153_11445.n3 a_3153_11445.n2 647.119
R23195 a_3153_11445.n1 a_3153_11445.t4 350.253
R23196 a_3153_11445.n2 a_3153_11445.n0 260.339
R23197 a_3153_11445.n2 a_3153_11445.n1 246.119
R23198 a_3153_11445.n1 a_3153_11445.t5 189.588
R23199 a_3153_11445.n3 a_3153_11445.t0 89.1195
R23200 a_3153_11445.n0 a_3153_11445.t1 63.3338
R23201 a_3153_11445.t2 a_3153_11445.n3 41.0422
R23202 a_3153_11445.n0 a_3153_11445.t3 31.9797
R23203 a_3500_11849.n3 a_3500_11849.n2 636.953
R23204 a_3500_11849.n1 a_3500_11849.t4 366.856
R23205 a_3500_11849.n2 a_3500_11849.n0 300.2
R23206 a_3500_11849.n2 a_3500_11849.n1 225.036
R23207 a_3500_11849.n1 a_3500_11849.t5 174.056
R23208 a_3500_11849.n0 a_3500_11849.t2 70.0005
R23209 a_3500_11849.t0 a_3500_11849.n3 68.0124
R23210 a_3500_11849.n3 a_3500_11849.t3 63.3219
R23211 a_3500_11849.n0 a_3500_11849.t1 61.6672
R23212 a_6888_11837.n1 a_6888_11837.n0 926.024
R23213 a_6888_11837.t0 a_6888_11837.n1 82.0838
R23214 a_6888_11837.n0 a_6888_11837.t1 63.3338
R23215 a_6888_11837.n1 a_6888_11837.t2 63.3219
R23216 a_6888_11837.n0 a_6888_11837.t3 29.7268
R23217 a_4550_9117.n3 a_4550_9117.n2 647.119
R23218 a_4550_9117.n1 a_4550_9117.t4 350.253
R23219 a_4550_9117.n2 a_4550_9117.n0 260.339
R23220 a_4550_9117.n2 a_4550_9117.n1 246.119
R23221 a_4550_9117.n1 a_4550_9117.t5 189.588
R23222 a_4550_9117.n3 a_4550_9117.t3 89.1195
R23223 a_4550_9117.n0 a_4550_9117.t0 63.3338
R23224 a_4550_9117.t1 a_4550_9117.n3 41.0422
R23225 a_4550_9117.n0 a_4550_9117.t2 31.9797
R23226 a_4857_8751.t0 a_4857_8751.t1 60.0005
R23227 a_8170_11293.t0 a_8170_11293.t1 126.644
R23228 a_10492_9673.n3 a_10492_9673.n2 636.953
R23229 a_10492_9673.n1 a_10492_9673.t4 366.856
R23230 a_10492_9673.n2 a_10492_9673.n0 300.2
R23231 a_10492_9673.n2 a_10492_9673.n1 225.036
R23232 a_10492_9673.n1 a_10492_9673.t5 174.056
R23233 a_10492_9673.n0 a_10492_9673.t2 70.0005
R23234 a_10492_9673.t0 a_10492_9673.n3 68.0124
R23235 a_10492_9673.n3 a_10492_9673.t3 63.3219
R23236 a_10492_9673.n0 a_10492_9673.t1 61.6672
R23237 a_10601_9673.n0 a_10601_9673.t0 68.3338
R23238 a_10601_9673.n0 a_10601_9673.t1 26.3935
R23239 a_10601_9673.n1 a_10601_9673.n0 14.4005
R23240 a_2157_7663.t0 a_2157_7663.t1 87.1434
R23241 a_10016_3311.n1 a_10016_3311.n0 926.024
R23242 a_10016_3311.t0 a_10016_3311.n1 82.0838
R23243 a_10016_3311.n0 a_10016_3311.t3 63.3338
R23244 a_10016_3311.n1 a_10016_3311.t1 63.3219
R23245 a_10016_3311.n0 a_10016_3311.t2 29.7268
R23246 a_5041_7663.t0 a_5041_7663.t1 60.0005
R23247 a_2564_10749.n1 a_2564_10749.n0 926.024
R23248 a_2564_10749.t1 a_2564_10749.n1 82.0838
R23249 a_2564_10749.n0 a_2564_10749.t0 63.3338
R23250 a_2564_10749.n1 a_2564_10749.t2 63.3219
R23251 a_2564_10749.n0 a_2564_10749.t3 29.7268
R23252 a_9575_8029.n0 a_9575_8029.t2 1327.82
R23253 a_9575_8029.n0 a_9575_8029.t1 194.655
R23254 a_9575_8029.t0 a_9575_8029.n0 63.3219
R23255 x2/net8.n4 x2/net8.n3 585
R23256 x2/net8.n5 x2/net8.n4 585
R23257 x2/net8.n2 x2/net8.t5 333.651
R23258 x2/net8.n2 x2/net8.t4 297.233
R23259 x2/net8 x2/net8.n2 194.062
R23260 x2/net8.n1 x2/net8.n0 185
R23261 x2/net8 x2/net8.n1 49.0339
R23262 x2/net8.n4 x2/net8.t0 26.5955
R23263 x2/net8.n4 x2/net8.t1 26.5955
R23264 x2/net8.n0 x2/net8.t2 24.9236
R23265 x2/net8.n0 x2/net8.t3 24.9236
R23266 x2/net8.n5 x2/net8 15.6165
R23267 x2/net8.n3 x2/net8 12.2206
R23268 x2/net8.n1 x2/net8 10.4965
R23269 x2/net8.n3 x2/net8 1.7925
R23270 x2/net8 x2/net8.n5 1.7925
R23271 a_3197_11837.t0 a_3197_11837.t1 60.0005
R23272 a_5481_3133.t0 a_5481_3133.t1 198.571
R23273 a_4948_8029.n0 a_4948_8029.t1 1327.82
R23274 a_4948_8029.n0 a_4948_8029.t2 194.655
R23275 a_4948_8029.t0 a_4948_8029.n0 63.3219
R23276 x2/net1.n3 x2/net1.n2 585
R23277 x2/net1.n4 x2/net1.n3 585
R23278 x2/net1.n5 x2/net1.t5 333.651
R23279 x2/net1.n5 x2/net1.t4 297.233
R23280 x2/net1 x2/net1.n5 196.493
R23281 x2/net1.n1 x2/net1.n0 185
R23282 x2/net1 x2/net1.n1 57.7379
R23283 x2/net1.n3 x2/net1.t1 26.5955
R23284 x2/net1.n3 x2/net1.t0 26.5955
R23285 x2/net1.n0 x2/net1.t3 24.9236
R23286 x2/net1.n0 x2/net1.t2 24.9236
R23287 x2/net1.n6 x2/net1 21.7272
R23288 x2/net1.n2 x2/net1 10.4965
R23289 x2/net1.n4 x2/net1 10.4965
R23290 x2/net1.n2 x2/net1 6.9125
R23291 x2/net1 x2/net1.n6 4.3525
R23292 x2/net1.n6 x2/net1.n4 2.5605
R23293 x2/net1.n1 x2/net1 1.7925
R23294 a_9221_10761.n0 a_9221_10761.t0 68.3338
R23295 a_9221_10761.n0 a_9221_10761.t1 26.3935
R23296 a_9221_10761.n1 a_9221_10761.n0 14.4005
R23297 a_8809_10749.t0 a_8809_10749.t1 60.0005
R23298 a_7158_8029.t0 a_7158_8029.t1 126.644
R23299 a_2372_8207.n0 a_2372_8207.t2 1327.82
R23300 a_2372_8207.n0 a_2372_8207.t1 194.655
R23301 a_2372_8207.t0 a_2372_8207.n0 63.3219
R23302 a_9667_7119.n0 a_9667_7119.t1 1327.82
R23303 a_9667_7119.t0 a_9667_7119.n0 194.655
R23304 a_9667_7119.n0 a_9667_7119.t2 63.3219
R23305 a_2029_8751.n0 a_2029_8751.t0 68.3338
R23306 a_2029_8751.n0 a_2029_8751.t1 26.3935
R23307 a_2029_8751.n1 a_2029_8751.n0 14.4005
R23308 a_6053_3311.t0 a_6053_3311.t1 60.0005
R23309 a_9563_8751.t1 a_9563_8751.t0 198.571
R23310 a_9729_8751.t0 a_9729_8751.t1 60.0005
R23311 a_6102_5853.n1 a_6102_5853.n0 926.024
R23312 a_6102_5853.n1 a_6102_5853.t3 82.0838
R23313 a_6102_5853.n0 a_6102_5853.t2 63.3338
R23314 a_6102_5853.t0 a_6102_5853.n1 63.3219
R23315 a_6102_5853.n0 a_6102_5853.t1 29.7268
R23316 a_4857_6575.t0 a_4857_6575.t1 60.0005
R23317 a_4503_12015.t0 a_4503_12015.t1 198.571
R23318 a_5619_11293.n0 a_5619_11293.t1 1327.82
R23319 a_5619_11293.n0 a_5619_11293.t2 194.655
R23320 a_5619_11293.t0 a_5619_11293.n0 63.3219
R23321 a_2790_8207.n1 a_2790_8207.n0 926.024
R23322 a_2790_8207.t0 a_2790_8207.n1 82.0838
R23323 a_2790_8207.n0 a_2790_8207.t1 63.3338
R23324 a_2790_8207.n1 a_2790_8207.t2 63.3219
R23325 a_2790_8207.n0 a_2790_8207.t3 29.7268
R23326 a_5409_3133.t0 a_5409_3133.t1 60.0005
R23327 a_2122_7915.n3 a_2122_7915.n2 636.953
R23328 a_2122_7915.n1 a_2122_7915.t4 366.856
R23329 a_2122_7915.n2 a_2122_7915.n0 300.2
R23330 a_2122_7915.n2 a_2122_7915.n1 225.036
R23331 a_2122_7915.n1 a_2122_7915.t5 174.056
R23332 a_2122_7915.n0 a_2122_7915.t3 70.0005
R23333 a_2122_7915.t0 a_2122_7915.n3 68.0124
R23334 a_2122_7915.n3 a_2122_7915.t2 63.3219
R23335 a_2122_7915.n0 a_2122_7915.t1 61.6672
R23336 a_6527_7663.t0 a_6527_7663.t1 198.571
R23337 SWN[3].n4 SWN[3].n3 585
R23338 SWN[3].n3 SWN[3].n2 585
R23339 SWN[3].n1 SWN[3].n0 185
R23340 SWN[3] SWN[3].n1 49.0339
R23341 SWN[3].n2 SWN[3] 28.327
R23342 SWN[3].n3 SWN[3].t1 26.5955
R23343 SWN[3].n3 SWN[3].t0 26.5955
R23344 SWN[3].n0 SWN[3].t2 24.9236
R23345 SWN[3].n0 SWN[3].t3 24.9236
R23346 SWN[3].n4 SWN[3] 15.6165
R23347 SWN[3].n1 SWN[3] 10.4965
R23348 SWN[3].n2 SWN[3] 1.7925
R23349 SWN[3] SWN[3].n4 1.7925
R23350 a_4932_2767.t0 a_4932_2767.t1 126.644
R23351 a_5133_10749.t0 a_5133_10749.t1 60.0005
R23352 a_5205_10749.t0 a_5205_10749.t1 198.571
R23353 a_5102_2767.n3 a_5102_2767.n2 647.119
R23354 a_5102_2767.n1 a_5102_2767.t4 350.253
R23355 a_5102_2767.n2 a_5102_2767.n0 260.339
R23356 a_5102_2767.n2 a_5102_2767.n1 246.119
R23357 a_5102_2767.n1 a_5102_2767.t5 189.588
R23358 a_5102_2767.n3 a_5102_2767.t0 89.1195
R23359 a_5102_2767.n0 a_5102_2767.t3 63.3338
R23360 a_5102_2767.t1 a_5102_2767.n3 41.0422
R23361 a_5102_2767.n0 a_5102_2767.t2 31.9797
R23362 a_5684_5853.n0 a_5684_5853.t1 1327.82
R23363 a_5684_5853.n0 a_5684_5853.t2 194.655
R23364 a_5684_5853.t0 a_5684_5853.n0 63.3219
R23365 a_7810_8573.t0 a_7810_8573.t1 87.1434
R23366 a_4697_10749.t0 a_4697_10749.t1 94.7268
R23367 a_6983_11849.n3 a_6983_11849.n2 674.338
R23368 a_6983_11849.n1 a_6983_11849.t4 332.58
R23369 a_6983_11849.n2 a_6983_11849.n0 284.012
R23370 a_6983_11849.n2 a_6983_11849.n1 253.648
R23371 a_6983_11849.n1 a_6983_11849.t5 168.701
R23372 a_6983_11849.n3 a_6983_11849.t3 96.1553
R23373 a_6983_11849.t1 a_6983_11849.n3 65.6672
R23374 a_6983_11849.n0 a_6983_11849.t2 65.0005
R23375 a_6983_11849.n0 a_6983_11849.t0 45.0005
R23376 a_10746_2767.t0 a_10746_2767.t1 126.644
R23377 a_2356_10205.t0 a_2356_10205.t1 126.644
R23378 a_5416_10927.n1 a_5416_10927.n0 926.024
R23379 a_5416_10927.n1 a_5416_10927.t3 82.0838
R23380 a_5416_10927.n0 a_5416_10927.t2 63.3338
R23381 a_5416_10927.t0 a_5416_10927.n1 63.3219
R23382 a_5416_10927.n0 a_5416_10927.t1 29.7268
R23383 a_4057_12015.t0 a_4057_12015.n3 370.026
R23384 a_4057_12015.n0 a_4057_12015.t5 351.356
R23385 a_4057_12015.n1 a_4057_12015.t2 334.717
R23386 a_4057_12015.n3 a_4057_12015.t1 325.971
R23387 a_4057_12015.n1 a_4057_12015.t4 309.935
R23388 a_4057_12015.n0 a_4057_12015.t3 305.683
R23389 a_4057_12015.n2 a_4057_12015.n0 16.879
R23390 a_4057_12015.n3 a_4057_12015.n2 10.8867
R23391 a_4057_12015.n2 a_4057_12015.n1 9.3005
R23392 a_10299_6575.t1 a_10299_6575.t0 198.571
R23393 a_10281_6397.t0 a_10281_6397.t1 60.0005
R23394 a_7365_3133.t1 a_7365_3133.t0 94.7268
R23395 a_5182_9117.n1 a_5182_9117.n0 926.024
R23396 a_5182_9117.t0 a_5182_9117.n1 82.0838
R23397 a_5182_9117.n0 a_5182_9117.t3 63.3338
R23398 a_5182_9117.n1 a_5182_9117.t1 63.3219
R23399 a_5182_9117.n0 a_5182_9117.t2 29.7268
R23400 a_10194_9117.t0 a_10194_9117.t1 126.644
R23401 a_10938_6397.t0 a_10938_6397.t1 87.1434
R23402 a_6999_8207.n0 a_6999_8207.t1 1327.82
R23403 a_6999_8207.t0 a_6999_8207.n0 194.655
R23404 a_6999_8207.n0 a_6999_8207.t2 63.3219
R23405 a_3043_11471.n0 a_3043_11471.t2 1327.82
R23406 a_3043_11471.t0 a_3043_11471.n0 194.655
R23407 a_3043_11471.n0 a_3043_11471.t1 63.3219
R23408 a_4764_9117.t0 a_4764_9117.n0 1327.82
R23409 a_4764_9117.n0 a_4764_9117.t2 194.655
R23410 a_4764_9117.n0 a_4764_9117.t1 63.3219
R23411 a_3905_5309.t0 a_3905_5309.t1 87.1434
R23412 a_3854_11837.t0 a_3854_11837.t1 87.1434
R23413 a_4733_11837.t0 a_4733_11837.t1 87.1434
R23414 a_8008_5487.n3 a_8008_5487.n2 636.953
R23415 a_8008_5487.n1 a_8008_5487.t5 366.856
R23416 a_8008_5487.n2 a_8008_5487.n0 300.2
R23417 a_8008_5487.n2 a_8008_5487.n1 225.036
R23418 a_8008_5487.n1 a_8008_5487.t4 174.056
R23419 a_8008_5487.n0 a_8008_5487.t0 70.0005
R23420 a_8008_5487.n3 a_8008_5487.t3 68.0124
R23421 a_8008_5487.t1 a_8008_5487.n3 63.3219
R23422 a_8008_5487.n0 a_8008_5487.t2 61.6672
R23423 a_5015_11713.n1 a_5015_11713.t6 530.01
R23424 a_5015_11713.t0 a_5015_11713.n5 421.021
R23425 a_5015_11713.n0 a_5015_11713.t3 337.171
R23426 a_5015_11713.n3 a_5015_11713.t1 280.223
R23427 a_5015_11713.n4 a_5015_11713.t2 263.173
R23428 a_5015_11713.n4 a_5015_11713.t4 227.826
R23429 a_5015_11713.n0 a_5015_11713.t7 199.762
R23430 a_5015_11713.n2 a_5015_11713.n1 170.81
R23431 a_5015_11713.n2 a_5015_11713.n0 167.321
R23432 a_5015_11713.n5 a_5015_11713.n4 152
R23433 a_5015_11713.n1 a_5015_11713.t5 141.923
R23434 a_5015_11713.n3 a_5015_11713.n2 10.8376
R23435 a_5015_11713.n5 a_5015_11713.n3 2.50485
R23436 a_4973_3133.t1 a_4973_3133.t0 94.7268
R23437 a_2790_9117.n1 a_2790_9117.n0 926.024
R23438 a_2790_9117.t0 a_2790_9117.n1 82.0838
R23439 a_2790_9117.n0 a_2790_9117.t1 63.3338
R23440 a_2790_9117.n1 a_2790_9117.t2 63.3219
R23441 a_2790_9117.n0 a_2790_9117.t3 29.7268
R23442 a_9927_5321.n3 a_9927_5321.n2 674.338
R23443 a_9927_5321.n1 a_9927_5321.t4 332.58
R23444 a_9927_5321.n2 a_9927_5321.n0 284.012
R23445 a_9927_5321.n2 a_9927_5321.n1 253.648
R23446 a_9927_5321.n1 a_9927_5321.t5 168.701
R23447 a_9927_5321.t0 a_9927_5321.n3 96.1553
R23448 a_9927_5321.n3 a_9927_5321.t3 65.6672
R23449 a_9927_5321.n0 a_9927_5321.t1 65.0005
R23450 a_9927_5321.n0 a_9927_5321.t2 45.0005
R23451 a_2833_7663.t0 a_2833_7663.t1 60.0005
R23452 a_10023_9673.t1 a_10023_9673.t0 198.571
R23453 a_10189_9661.t0 a_10189_9661.t1 60.0005
R23454 a_10141_10927.t1 a_10141_10927.t0 94.7268
R23455 a_5316_11471.n0 a_5316_11471.t1 1327.82
R23456 a_5316_11471.n0 a_5316_11471.t2 194.655
R23457 a_5316_11471.t0 a_5316_11471.n0 63.3219
R23458 a_9832_5309.n1 a_9832_5309.n0 926.024
R23459 a_9832_5309.n1 a_9832_5309.t3 82.0838
R23460 a_9832_5309.n0 a_9832_5309.t0 63.3338
R23461 a_9832_5309.t1 a_9832_5309.n1 63.3219
R23462 a_9832_5309.n0 a_9832_5309.t2 29.7268
R23463 a_5171_11445.n3 a_5171_11445.n2 674.338
R23464 a_5171_11445.n1 a_5171_11445.t4 332.58
R23465 a_5171_11445.n2 a_5171_11445.n0 284.012
R23466 a_5171_11445.n2 a_5171_11445.n1 253.648
R23467 a_5171_11445.n1 a_5171_11445.t5 168.701
R23468 a_5171_11445.n3 a_5171_11445.t2 96.1553
R23469 a_5171_11445.t0 a_5171_11445.n3 65.6672
R23470 a_5171_11445.n0 a_5171_11445.t3 65.0005
R23471 a_5171_11445.n0 a_5171_11445.t1 45.0005
R23472 a_9563_10927.t1 a_9563_10927.t0 198.571
R23473 a_4329_8573.t1 a_4329_8573.t0 94.7268
R23474 a_11122_6575.t0 a_11122_6575.t1 87.1434
R23475 a_6238_11293.t0 a_6238_11293.t1 126.644
R23476 a_6336_7663.n1 a_6336_7663.n0 926.024
R23477 a_6336_7663.t1 a_6336_7663.n1 82.0838
R23478 a_6336_7663.n0 a_6336_7663.t0 63.3338
R23479 a_6336_7663.n1 a_6336_7663.t2 63.3219
R23480 a_6336_7663.n0 a_6336_7663.t3 29.7268
R23481 a_10601_9839.t1 a_10601_9839.t0 94.7268
R23482 a_9924_3133.n1 a_9924_3133.n0 926.024
R23483 a_9924_3133.n1 a_9924_3133.t3 82.0838
R23484 a_9924_3133.n0 a_9924_3133.t2 63.3338
R23485 a_9924_3133.t0 a_9924_3133.n1 63.3219
R23486 a_9924_3133.n0 a_9924_3133.t1 29.7268
R23487 a_5607_10927.t0 a_5607_10927.t1 198.571
R23488 a_5773_10927.t0 a_5773_10927.t1 60.0005
R23489 a_10785_3311.t1 a_10785_3311.t0 94.7268
R23490 a_10189_9839.t0 a_10189_9839.t1 60.0005
R23491 a_10373_3311.t0 a_10373_3311.t1 60.0005
R23492 a_10141_7663.t0 a_10141_7663.t1 94.7268
R23493 a_2157_4399.t0 a_2157_4399.t1 87.1434
R23494 a_5849_5487.t0 a_5849_5487.t1 198.571
R23495 a_8547_10761.n3 a_8547_10761.n2 674.338
R23496 a_8547_10761.n1 a_8547_10761.t4 332.58
R23497 a_8547_10761.n2 a_8547_10761.n0 284.012
R23498 a_8547_10761.n2 a_8547_10761.n1 253.648
R23499 a_8547_10761.n1 a_8547_10761.t5 168.701
R23500 a_8547_10761.t0 a_8547_10761.n3 96.1553
R23501 a_8547_10761.n3 a_8547_10761.t2 65.6672
R23502 a_8547_10761.n0 a_8547_10761.t3 65.0005
R23503 a_8547_10761.n0 a_8547_10761.t1 45.0005
R23504 a_8765_10357.n3 a_8765_10357.n2 647.119
R23505 a_8765_10357.n1 a_8765_10357.t4 350.253
R23506 a_8765_10357.n2 a_8765_10357.n0 260.339
R23507 a_8765_10357.n2 a_8765_10357.n1 246.119
R23508 a_8765_10357.n1 a_8765_10357.t5 189.588
R23509 a_8765_10357.n3 a_8765_10357.t0 89.1195
R23510 a_8765_10357.n0 a_8765_10357.t1 63.3338
R23511 a_8765_10357.t2 a_8765_10357.n3 41.0422
R23512 a_8765_10357.n0 a_8765_10357.t3 31.9797
R23513 a_4803_7900.n3 a_4803_7900.n2 674.338
R23514 a_4803_7900.n1 a_4803_7900.t4 332.58
R23515 a_4803_7900.n2 a_4803_7900.n0 284.012
R23516 a_4803_7900.n2 a_4803_7900.n1 253.648
R23517 a_4803_7900.n1 a_4803_7900.t5 168.701
R23518 a_4803_7900.t0 a_4803_7900.n3 96.1553
R23519 a_4803_7900.n3 a_4803_7900.t2 65.6672
R23520 a_4803_7900.n0 a_4803_7900.t1 65.0005
R23521 a_4803_7900.n0 a_4803_7900.t3 45.0005
R23522 a_8031_10389.n1 a_8031_10389.t6 530.01
R23523 a_8031_10389.t0 a_8031_10389.n5 421.021
R23524 a_8031_10389.n0 a_8031_10389.t4 337.142
R23525 a_8031_10389.n3 a_8031_10389.t1 280.223
R23526 a_8031_10389.n4 a_8031_10389.t5 263.173
R23527 a_8031_10389.n4 a_8031_10389.t7 227.826
R23528 a_8031_10389.n0 a_8031_10389.t3 199.762
R23529 a_8031_10389.n2 a_8031_10389.n1 170.81
R23530 a_8031_10389.n2 a_8031_10389.n0 167.321
R23531 a_8031_10389.n5 a_8031_10389.n4 152
R23532 a_8031_10389.n1 a_8031_10389.t2 141.923
R23533 a_8031_10389.n3 a_8031_10389.n2 10.8376
R23534 a_8031_10389.n5 a_8031_10389.n3 2.50485
R23535 a_4181_6575.t0 a_4181_6575.t1 87.1434
R23536 a_2721_5309.t0 a_2721_5309.t1 198.571
R23537 a_2740_4765.n0 a_2740_4765.t1 1327.82
R23538 a_2740_4765.n0 a_2740_4765.t2 194.655
R23539 a_2740_4765.t0 a_2740_4765.n0 63.3219
R23540 a_10478_7485.t0 a_10478_7485.t1 87.1434
R23541 a_2755_10761.t0 a_2755_10761.t1 198.571
R23542 a_2921_10749.t0 a_2921_10749.t1 60.0005
R23543 a_2356_5853.t0 a_2356_5853.t1 126.644
R23544 a_10693_4233.n0 a_10693_4233.t0 68.3338
R23545 a_10693_4233.n0 a_10693_4233.t1 26.3935
R23546 a_10693_4233.n1 a_10693_4233.n0 14.4005
R23547 a_10846_9661.t0 a_10846_9661.t1 87.1434
R23548 a_4104_4943.t0 a_4104_4943.t1 126.644
R23549 a_5182_4765.n1 a_5182_4765.n0 926.024
R23550 a_5182_4765.n1 a_5182_4765.t3 82.0838
R23551 a_5182_4765.n0 a_5182_4765.t2 63.3338
R23552 a_5182_4765.t0 a_5182_4765.n1 63.3219
R23553 a_5182_4765.n0 a_5182_4765.t1 29.7268
R23554 a_9927_9673.n3 a_9927_9673.n2 674.338
R23555 a_9927_9673.n1 a_9927_9673.t5 332.58
R23556 a_9927_9673.n2 a_9927_9673.n0 284.012
R23557 a_9927_9673.n2 a_9927_9673.n1 253.648
R23558 a_9927_9673.n1 a_9927_9673.t4 168.701
R23559 a_9927_9673.t0 a_9927_9673.n3 96.1553
R23560 a_9927_9673.n3 a_9927_9673.t3 65.6672
R23561 a_9927_9673.n0 a_9927_9673.t1 65.0005
R23562 a_9927_9673.n0 a_9927_9673.t2 45.0005
R23563 a_9466_10749.t0 a_9466_10749.t1 87.1434
R23564 a_10846_9839.t0 a_10846_9839.t1 87.1434
R23565 a_10930_6941.t0 a_10930_6941.t1 126.644
R23566 a_7631_6409.t0 a_7631_6409.t1 198.571
R23567 a_9777_7093.n3 a_9777_7093.n2 647.119
R23568 a_9777_7093.n1 a_9777_7093.t4 350.253
R23569 a_9777_7093.n2 a_9777_7093.n0 260.339
R23570 a_9777_7093.n2 a_9777_7093.n1 246.119
R23571 a_9777_7093.n1 a_9777_7093.t5 189.588
R23572 a_9777_7093.n3 a_9777_7093.t2 89.1195
R23573 a_9777_7093.n0 a_9777_7093.t3 63.3338
R23574 a_9777_7093.t0 a_9777_7093.n3 41.0422
R23575 a_9777_7093.n0 a_9777_7093.t1 31.9797
R23576 a_9821_7485.t0 a_9821_7485.t1 60.0005
R23577 a_4929_6575.t1 a_4929_6575.t0 198.571
R23578 a_8643_10761.t1 a_8643_10761.t0 198.571
R23579 a_5481_6397.t0 a_5481_6397.t1 198.571
R23580 a_10386_8751.t0 a_10386_8751.t1 87.1434
R23581 a_10019_3145.n3 a_10019_3145.n2 674.338
R23582 a_10019_3145.n1 a_10019_3145.t5 332.58
R23583 a_10019_3145.n2 a_10019_3145.n0 284.012
R23584 a_10019_3145.n2 a_10019_3145.n1 253.648
R23585 a_10019_3145.n1 a_10019_3145.t4 168.701
R23586 a_10019_3145.t0 a_10019_3145.n3 96.1553
R23587 a_10019_3145.n3 a_10019_3145.t3 65.6672
R23588 a_10019_3145.n0 a_10019_3145.t1 65.0005
R23589 a_10019_3145.n0 a_10019_3145.t2 45.0005
R23590 a_10115_3145.t0 a_10115_3145.t1 198.571
R23591 a_2740_10205.n0 a_2740_10205.t1 1327.82
R23592 a_2740_10205.t0 a_2740_10205.n0 194.655
R23593 a_2740_10205.n0 a_2740_10205.t2 63.3219
R23594 a_11030_5487.t0 a_11030_5487.t1 87.1434
R23595 a_4457_10749.t0 a_4457_10749.t1 87.1434
R23596 a_7324_2767.t0 a_7324_2767.t1 126.644
R23597 a_2157_9839.t0 a_2157_9839.t1 87.1434
R23598 a_3158_5853.n1 a_3158_5853.n0 926.024
R23599 a_3158_5853.t1 a_3158_5853.n1 82.0838
R23600 a_3158_5853.n0 a_3158_5853.t0 63.3338
R23601 a_3158_5853.n1 a_3158_5853.t2 63.3219
R23602 a_3158_5853.n0 a_3158_5853.t3 29.7268
R23603 a_10281_3133.t0 a_10281_3133.t1 60.0005
R23604 a_8393_4233.n0 a_8393_4233.t1 68.3338
R23605 a_8393_4233.n0 a_8393_4233.t0 26.3935
R23606 a_8393_4233.n1 a_8393_4233.n0 14.4005
R23607 a_10938_3133.t0 a_10938_3133.t1 87.1434
R23608 a_7815_4233.t0 a_7815_4233.t1 198.571
R23609 a_2649_5309.t0 a_2649_5309.t1 60.0005
R23610 a_10386_10927.t0 a_10386_10927.t1 87.1434
R23611 a_2213_5309.t1 a_2213_5309.t0 94.7268
R23612 a_5777_5487.t0 a_5777_5487.t1 60.0005
R23613 a_7079_11849.t1 a_7079_11849.t0 198.571
R23614 a_4656_10383.t0 a_4656_10383.t1 126.644
R23615 a_8655_10383.n0 a_8655_10383.t2 1327.82
R23616 a_8655_10383.n0 a_8655_10383.t1 194.655
R23617 a_8655_10383.t0 a_8655_10383.n0 63.3219
R23618 a_8117_5487.t1 a_8117_5487.t0 94.7268
R23619 a_2905_7663.t0 a_2905_7663.t1 198.571
R23620 a_2397_7663.n0 a_2397_7663.t1 68.3338
R23621 a_2397_7663.n0 a_2397_7663.t0 26.3935
R23622 a_2397_7663.n1 a_2397_7663.n0 14.4005
R23623 a_7933_4399.t0 a_7933_4399.t1 94.7268
R23624 a_7245_11837.t0 a_7245_11837.t1 60.0005
R23625 a_1988_9117.t0 a_1988_9117.t1 126.644
R23626 a_6378_3677.n1 a_6378_3677.n0 926.024
R23627 a_6378_3677.n1 a_6378_3677.t3 82.0838
R23628 a_6378_3677.n0 a_6378_3677.t2 63.3338
R23629 a_6378_3677.t0 a_6378_3677.n1 63.3219
R23630 a_6378_3677.n0 a_6378_3677.t1 29.7268
R23631 a_8362_5487.t0 a_8362_5487.t1 87.1434
R23632 a_1988_8207.t0 a_1988_8207.t1 126.644
R23633 a_10838_5853.t0 a_10838_5853.t1 126.644
R23634 a_1789_8573.t0 a_1789_8573.t1 87.1434
R23635 a_7902_11837.t0 a_7902_11837.t1 87.1434
R23636 a_5113_7663.t0 a_5113_7663.t1 198.571
R23637 a_3578_10749.t0 a_3578_10749.t1 87.1434
R23638 a_7986_4765.t0 a_7986_4765.t1 126.644
R23639 a_2157_5487.t0 a_2157_5487.t1 87.1434
R23640 a_5101_5487.t0 a_5101_5487.t1 87.1434
R23641 a_6693_7663.t0 a_6693_7663.t1 60.0005
R23642 a_7705_3311.t0 a_7705_3311.t1 60.0005
R23643 a_10465_6575.t0 a_10465_6575.t1 60.0005
R23644 a_7797_6397.t0 a_7797_6397.t1 60.0005
R23645 a_10115_4233.t0 a_10115_4233.t1 198.571
R23646 a_8117_10927.t1 a_8117_10927.t0 94.7268
R23647 a_10938_4221.t0 a_10938_4221.t1 87.1434
R23648 a_4733_6397.t0 a_4733_6397.t1 87.1434
C0 x2/net6 x2/net13 0.02875f
C1 clknet_1_1__leaf_CLK x2/net2 0.180971f
C2 DOUT[5] DOUT[6] 0.623568f
C3 x2/net6 SWN[1] 0.036799f
C4 CF[6] CF[9] 0.024426f
C5 CKO CF[5] 0.10093f
C6 CKO SWP[2] 0.044087f
C7 CF[7] SWN[9] 0.239031f
C8 SWP[8] SWP[3] 0.042477f
C9 EN SWN[3] 0.144684f
C10 x3/COMP_BUF_P CF[2] 0.075709f
C11 x3/COMP_BUF_P DOUT[5] 0.050276f
C12 clknet_1_1__leaf_CLK x2/net8 0.052035f
C13 x2/net13 CLKS 0.864784f
C14 x3/COMP_BUF_N CF[5] 1.37051f
C15 EN DOUT[2] 0.090076f
C16 CLKS SWN[1] 0.026046f
C17 CF[6] CF[2] 0.087219f
C18 SWP[9] SWN[6] 0.037011f
C19 EN SWN[7] 0.124426f
C20 EN SWP[4] 0.221612f
C21 VDDD SWP[8] 2.08571f
C22 DOUT[9] SWN[1] 0.041174f
C23 CLK DOUT[3] 0.094231f
C24 COMP_P DOUT[3] 0.040582f
C25 x3/COMP_BUF_N SWN[9] 0.048631f
C26 clknet_1_0__leaf_CLK EN 0.016254f
C27 x2/net9 DOUT[7] 0.019131f
C28 clknet_0_CLK EN 0.315642f
C29 SWP[1] SWP[7] 0.068141f
C30 CLKS SWP[7] 0.679825f
C31 SWP[0] CF[5] 0.03218f
C32 SWP[0] SWP[2] 0.144313f
C33 SWP[8] CF[7] 0.012276f
C34 x3/COMP_BUF_P SWP[3] 0.058328f
C35 SWP[8] SWP[5] 0.041708f
C36 SWN[0] DOUT[7] 0.035391f
C37 clknet_1_1__leaf_CLK EN 1.87671f
C38 VDDD SWN[4] 1.27778f
C39 clknet_1_1__leaf_CLK x2/net1 0.110885f
C40 SWP[7] DOUT[9] 0.020614f
C41 SWP[2] SWP[9] 0.037287f
C42 CF[3] DOUT[6] 0.110708f
C43 CF[5] SWP[9] 0.966443f
C44 x2/net11 DOUT[4] 0.034125f
C45 VDDD SWN[2] 1.69527f
C46 VDDD DOUT[6] 2.02121f
C47 SWP[3] CF[6] 0.026255f
C48 SWP[0] SWN[9] 0.385956f
C49 CF[4] SWP[4] 0.023577f
C50 x3/COMP_BUF_P CF[3] 0.050691f
C51 x3/COMP_BUF_P VDDD 6.55023f
C52 clknet_0_CLK SWN[3] 0.074764f
C53 FINAL CF[4] 0.046696f
C54 x2/net5 EN 0.28253f
C55 x3/COMP_BUF_N SWP[8] 0.014671f
C56 clknet_1_0__leaf_CLK CF[4] 0.531711f
C57 EN DOUT[8] 1.33334f
C58 clknet_1_1__leaf_CLK SWN[3] 0.174339f
C59 CKO SWN[4] 0.080062f
C60 CF[0] CF[1] 0.589781f
C61 CF[3] CF[6] 0.025599f
C62 FINAL SWP[4] 0.178144f
C63 EN COMP_N 0.099628f
C64 x2/net4 x2/net11 0.016612f
C65 VDDD CF[6] 2.50788f
C66 clknet_1_0__leaf_CLK SWP[4] 0.049091f
C67 x2/TRIG2 x2/net6 0.037127f
C68 x3/COMP_BUF_P CF[7] 0.196288f
C69 x3/COMP_BUF_P SWP[5] 0.077101f
C70 CKO SWN[2] 0.022137f
C71 CLKS DOUT[3] 0.21641f
C72 CKO DOUT[6] 0.107337f
C73 clknet_0_CLK SWP[4] 0.025435f
C74 SWP[7] SWN[6] 0.047952f
C75 EN DOUT[5] 0.295931f
C76 clknet_0_CLK FINAL 0.385606f
C77 CF[6] CF[7] 0.394906f
C78 x3/COMP_BUF_P CKO 0.351403f
C79 SWP[0] SWP[8] 0.047648f
C80 SWP[1] CF[0] 0.065524f
C81 CLKS CF[0] 1.08162f
C82 SWP[5] CF[6] 0.023941f
C83 CF[0] CF[8] 0.020372f
C84 x3/COMP_BUF_N SWN[2] 0.179377f
C85 x2/net2 VDDD 0.580562f
C86 x3/COMP_BUF_N DOUT[6] 0.039329f
C87 DOUT[8] SWN[3] 0.041585f
C88 CF[4] CF[9] 0.020836f
C89 DOUT[7] SWN[1] 0.034767f
C90 clknet_1_1__leaf_CLK clknet_0_CLK 0.043152f
C91 SWN[0] SWN[4] 0.170789f
C92 VDDD DOUT[1] 0.861961f
C93 x2/net9 SWN[2] 0.014245f
C94 x3/COMP_BUF_N x3/COMP_BUF_P 0.140088f
C95 x2/net8 VDDD 0.77249f
C96 x2/TRIG2 DOUT[9] 0.022592f
C97 COMP_N DOUT[2] 0.038407f
C98 x2/net7 SWN[2] 0.030093f
C99 SWN[0] SWN[2] 0.109431f
C100 DOUT[0] COMP_P 0.221929f
C101 SWP[2] SWP[7] 0.059564f
C102 VDDD SWN[5] 0.335767f
C103 CLKS CLK 0.403272f
C104 x3/COMP_BUF_N CF[6] 0.026492f
C105 SWP[1] SWP[6] 0.04429f
C106 SWP[1] CLK 0.017543f
C107 CLKS SWP[6] 0.285389f
C108 clkload0.X SWP[4] 0.171861f
C109 clknet_1_0__leaf_CLK CF[9] 0.084131f
C110 CF[4] CF[2] 0.09812f
C111 SWP[6] CF[8] 0.093958f
C112 SWP[1] COMP_P 0.020601f
C113 SWP[9] SWN[4] 0.019962f
C114 SWP[7] DOUT[7] 0.069816f
C115 clknet_0_CLK CF[9] 0.015542f
C116 x3/COMP_BUF_P SWP[0] 0.063136f
C117 SWP[9] SWN[2] 0.022143f
C118 SWP[7] SWN[9] 0.034143f
C119 x2/net10 VDDD 0.440941f
C120 clknet_1_1__leaf_CLK DOUT[8] 0.04865f
C121 x2/net12 SWN[2] 0.032589f
C122 clknet_1_0__leaf_CLK CF[2] 0.040498f
C123 DOUT[6] DOUT[4] 0.022948f
C124 x3/COMP_BUF_P SWP[9] 0.029201f
C125 SWP[0] CF[6] 0.033274f
C126 clknet_0_CLK CF[2] 0.023188f
C127 VDDD EN 8.16485f
C128 CKO SWN[5] 0.142195f
C129 x2/net1 VDDD 1.1286f
C130 x2/net11 DOUT[3] 0.02765f
C131 clknet_1_1__leaf_CLK DOUT[5] 0.27076f
C132 SWP[1] CF[1] 0.032338f
C133 CLKS CF[1] 0.690374f
C134 CF[1] CF[8] 0.077979f
C135 SWP[9] CF[6] 0.374057f
C136 CF[4] SWP[3] 0.048285f
C137 x2/net4 DOUT[6] 0.023038f
C138 SWP[4] SWP[3] 0.578805f
C139 SWP[6] SWN[6] 0.275196f
C140 x2/net11 x2/TRIG2 0.052753f
C141 CF[0] SWP[2] 0.118489f
C142 SWP[8] SWP[7] 2.04122f
C143 x2/net13 SWN[2] 0.2195f
C144 CF[0] CF[5] 0.045581f
C145 SWP[1] CLKS 1.11109f
C146 VDDD SWN[3] 2.0913f
C147 CLKS CF[8] 0.936053f
C148 SWP[1] CF[8] 0.088345f
C149 EN CKO 0.107593f
C150 SWN[1] SWN[2] 0.486568f
C151 CF[9] CF[2] 0.321543f
C152 clknet_1_0__leaf_CLK SWP[3] 0.358502f
C153 CF[3] CF[4] 0.607457f
C154 VDDD CF[4] 2.46997f
C155 VDDD DOUT[2] 0.911187f
C156 COMP_N DOUT[5] 0.06647f
C157 x2/TRIG2 DOUT[7] 0.018462f
C158 x3/COMP_BUF_N EN 1.04605f
C159 CF[3] SWP[4] 0.024539f
C160 VDDD SWN[7] 1.38654f
C161 VDDD SWP[4] 2.24314f
C162 x2/net10 SWN[0] 0.016182f
C163 FINAL CF[3] 0.11438f
C164 CF[4] CF[7] 0.019657f
C165 clknet_1_0__leaf_CLK CF[3] 0.535504f
C166 CF[5] SWP[6] 0.022823f
C167 SWP[2] SWP[6] 0.047914f
C168 FINAL VDDD 2.12817f
C169 SWP[2] CLK 0.021818f
C170 SWP[5] CF[4] 1.8157f
C171 SWP[2] COMP_P 0.208997f
C172 clknet_1_0__leaf_CLK VDDD 4.28697f
C173 x2/net9 EN 0.217771f
C174 SWP[4] CF[7] 0.019468f
C175 clknet_0_CLK VDDD 2.63092f
C176 EN SWN[0] 0.720487f
C177 x2/net7 EN 0.024817f
C178 SWP[5] SWP[4] 0.4532f
C179 SWP[3] CF[9] 0.023384f
C180 CKO CF[4] 0.177601f
C181 clknet_1_1__leaf_CLK VDDD 6.42383f
C182 EN SWP[0] 0.083803f
C183 FINAL SWP[5] 0.028139f
C184 clknet_1_0__leaf_CLK CF[7] 0.429896f
C185 SWP[6] SWN[9] 0.014471f
C186 clknet_0_CLK CF[7] 0.219607f
C187 CKO SWP[4] 0.216079f
C188 x3/COMP_BUF_N CF[4] 0.085047f
C189 EN SWP[9] 0.018599f
C190 FINAL CKO 0.100541f
C191 clknet_1_0__leaf_CLK CKO 0.25605f
C192 SWP[3] CF[2] 0.065428f
C193 DOUT[9] SWN[6] 0.058104f
C194 CF[3] CF[9] 0.022881f
C195 CF[5] CF[1] 0.076172f
C196 SWP[2] CF[1] 0.047826f
C197 x3/COMP_BUF_N SWP[4] 0.374729f
C198 SWN[0] SWN[3] 0.038449f
C199 x2/net7 SWN[3] 0.064419f
C200 clknet_0_CLK CKO 0.020985f
C201 x2/net5 VDDD 0.436352f
C202 EN DOUT[4] 0.049569f
C203 VDDD CF[9] 3.05718f
C204 VDDD DOUT[8] 1.32961f
C205 DOUT[6] DOUT[3] 0.058953f
C206 x3/COMP_BUF_N FINAL 0.079385f
C207 VDDD COMP_N 1.3547f
C208 clkload0.X VDDD 0.756718f
C209 clknet_0_CLK x3/COMP_BUF_N 0.08933f
C210 SWP[0] CF[4] 0.025128f
C211 CF[9] CF[7] 0.336327f
C212 CLKS CF[5] 1.06387f
C213 SWP[1] SWP[2] 0.638919f
C214 CLKS SWP[2] 0.425127f
C215 COMP_N CLKSB 0.224871f
C216 SWP[1] CF[5] 0.033805f
C217 SWP[5] CF[9] 0.062184f
C218 CF[5] CF[8] 0.01532f
C219 CF[3] CF[2] 0.176269f
C220 SWP[2] CF[8] 0.020775f
C221 SWP[8] SWP[6] 0.258475f
C222 VDDD CF[2] 1.9956f
C223 x2/net10 SWN[1] 0.014076f
C224 VDDD DOUT[5] 1.05245f
C225 SWP[0] SWN[7] 0.01583f
C226 x2/net12 SWN[3] 0.036846f
C227 x2/TRIG2 SWN[2] 0.060043f
C228 SWP[0] SWP[4] 0.031427f
C229 x2/net4 EN 0.236925f
C230 SWP[9] CF[4] 0.494976f
C231 SWP[7] SWN[5] 0.01892f
C232 CKO CF[9] 0.193093f
C233 x3/COMP_BUF_P CF[0] 0.204923f
C234 CLKS SWN[9] 0.145958f
C235 clknet_1_1__leaf_CLK x2/net9 0.23047f
C236 CF[8] SWN[9] 0.400094f
C237 clknet_1_0__leaf_CLK SWP[0] 0.353713f
C238 CF[2] CF[7] 0.025957f
C239 EN SWN[1] 0.2277f
C240 SWP[5] CF[2] 0.017492f
C241 SWP[9] SWP[4] 0.044127f
C242 SWN[4] SWP[6] 0.062807f
C243 DOUT[7] DOUT[9] 0.633679f
C244 CKO COMP_N 0.080269f
C245 DOUT[2] DOUT[4] 1.3712f
C246 x2/net1 SWN[1] 0.053512f
C247 clknet_1_1__leaf_CLK x2/net7 0.097418f
C248 clkload0.X CKO 0.0163f
C249 clknet_1_1__leaf_CLK SWN[0] 0.451859f
C250 clknet_0_CLK SWP[0] 0.045258f
C251 x2/net3 x2/net11 0.159517f
C252 CF[0] CF[6] 0.026023f
C253 x3/COMP_BUF_N CF[9] 0.09783f
C254 FINAL SWP[9] 0.020132f
C255 SWP[6] SWN[2] 0.154514f
C256 COMP_P DOUT[6] 0.726518f
C257 CKO DOUT[5] 0.093707f
C258 x3/COMP_BUF_N clkload0.X 0.024086f
C259 x3/COMP_BUF_N COMP_N 0.012131f
C260 CF[3] SWP[3] 0.418991f
C261 SWN[8] SWN[9] 0.173118f
C262 VDDD SWP[3] 2.98632f
C263 EN SWP[7] 0.215752f
C264 x2/net13 SWN[3] 0.034937f
C265 x3/COMP_BUF_P SWP[6] 0.303049f
C266 x2/net9 DOUT[8] 0.017763f
C267 SWN[3] SWN[1] 0.17609f
C268 x3/COMP_BUF_N DOUT[5] 0.139406f
C269 DOUT[8] SWN[0] 0.032323f
C270 SWP[0] CF[9] 0.69914f
C271 SWP[3] CF[7] 0.02345f
C272 CLKS SWP[8] 0.136267f
C273 SWP[1] SWP[8] 0.069683f
C274 DOUT[7] SWN[6] 0.046916f
C275 SWP[5] SWP[3] 0.107526f
C276 SWP[8] CF[8] 0.08049f
C277 VDDD CF[3] 2.5081f
C278 x2/net6 SWN[2] 0.102433f
C279 COMP_N SWP[0] 0.024254f
C280 SWP[4] SWN[1] 0.13218f
C281 SWP[9] CF[9] 0.067153f
C282 SWP[8] DOUT[9] 0.018251f
C283 CKO SWP[3] 0.10161f
C284 VDDD CLKSB 0.367406f
C285 FINAL SWN[1] 0.025405f
C286 SWP[0] CF[2] 0.037279f
C287 CLKS SWN[4] 0.058823f
C288 CF[3] CF[7] 0.023444f
C289 x3/COMP_BUF_P CF[1] 0.934921f
C290 clknet_1_1__leaf_CLK x2/net4 0.143772f
C291 SWP[2] CF[5] 0.095478f
C292 VDDD CF[7] 1.75228f
C293 VDDD SWP[5] 1.86243f
C294 CLKS SWN[2] 0.777035f
C295 CLKS DOUT[6] 0.024449f
C296 COMP_N DOUT[4] 0.029996f
C297 DOUT[1] COMP_P 0.049955f
C298 EN DOUT[3] 0.413468f
C299 SWP[7] SWN[7] 0.713537f
C300 SWP[9] CF[2] 0.268968f
C301 clknet_1_1__leaf_CLK SWN[1] 0.354484f
C302 SWP[7] SWP[4] 0.059439f
C303 DOUT[9] SWN[4] 0.052338f
C304 CF[6] CF[1] 0.019931f
C305 CKO CF[3] 0.938675f
C306 VDDD CKO 7.42588f
C307 x2/TRIG1 EN 0.08758f
C308 SWP[5] CF[7] 0.017355f
C309 DOUT[9] SWN[2] 0.041276f
C310 x3/COMP_BUF_P SWP[1] 0.146774f
C311 x3/COMP_BUF_P CLKS 0.635905f
C312 EN CF[0] 0.013561f
C313 x3/COMP_BUF_P CF[8] 0.135365f
C314 DOUT[5] DOUT[4] 0.241837f
C315 SWP[8] SWN[6] 0.076729f
C316 x2/TRIG2 EN 1.1719f
C317 SWP[1] CF[6] 0.045934f
C318 SWP[0] SWP[3] 0.02043f
C319 CLKS CF[6] 0.571925f
C320 x3/COMP_BUF_N VDDD 4.65431f
C321 CF[6] CF[8] 0.018487f
C322 CKO SWP[5] 0.343635f
C323 DOUT[8] SWN[1] 0.029429f
C324 x2/net9 VDDD 1.08017f
C325 SWN[4] SWN[6] 0.201194f
C326 SWP[9] SWP[3] 0.041226f
C327 x3/COMP_BUF_N CF[7] 0.352679f
C328 DOUT[2] DOUT[3] 0.248577f
C329 EN CLK 0.431408f
C330 x3/COMP_BUF_N SWP[5] 0.044282f
C331 EN COMP_P 0.089435f
C332 x2/net7 VDDD 1.02412f
C333 VDDD SWN[0] 1.06477f
C334 x2/TRIG2 SWN[3] 0.01936f
C335 SWP[0] CF[3] 0.037476f
C336 DOUT[1] DOUT[0] 0.519039f
C337 CF[0] CF[4] 0.034114f
C338 VDDD SWP[0] 3.17338f
C339 SWP[8] SWP[2] 0.043558f
C340 x3/COMP_BUF_N CKO 0.111072f
C341 CF[0] SWP[4] 0.165705f
C342 SWP[8] DOUT[7] 0.185126f
C343 VDDD SWP[9] 1.36372f
C344 SWP[0] CF[7] 0.173895f
C345 FINAL CF[0] 0.271769f
C346 SWP[0] SWP[5] 0.02513f
C347 x2/net12 VDDD 0.588705f
C348 SWP[8] SWN[9] 0.068367f
C349 clknet_1_0__leaf_CLK CF[0] 0.224351f
C350 x2/net11 DOUT[6] 0.024879f
C351 VDDD DOUT[4] 0.720282f
C352 x2/net6 EN 0.447872f
C353 clknet_0_CLK CF[0] 0.19475f
C354 SWP[9] CF[7] 0.022508f
C355 x2/net2 x2/net3 0.030818f
C356 CF[4] SWP[6] 0.057766f
C357 DOUT[7] SWN[4] 0.03589f
C358 CKO SWP[0] 0.059067f
C359 SWP[5] SWP[9] 0.778272f
C360 SWP[2] DOUT[6] 0.133444f
C361 SWN[5] DOUT[9] 0.018675f
C362 DOUT[2] COMP_P 0.053238f
C363 clknet_1_1__leaf_CLK x2/TRIG2 0.289214f
C364 DOUT[7] SWN[2] 0.034971f
C365 SWP[6] SWP[4] 0.116164f
C366 x3/COMP_BUF_P SWP[2] 0.112413f
C367 x3/COMP_BUF_P CF[5] 0.083154f
C368 x2/net5 DOUT[3] 0.027711f
C369 CKO SWP[9] 0.037108f
C370 x3/COMP_BUF_N SWP[0] 0.054965f
C371 EN SWP[1] 0.650903f
C372 EN CLKS 0.105082f
C373 FINAL CLK 0.086438f
C374 x2/net4 VDDD 0.456021f
C375 clknet_1_0__leaf_CLK CLK 0.021107f
C376 COMP_N DOUT[3] 0.036631f
C377 x2/net13 VDDD 0.902092f
C378 x2/net6 SWN[3] 0.066246f
C379 CF[5] CF[6] 0.409172f
C380 CF[0] CF[9] 0.06305f
C381 SWP[2] CF[6] 0.257441f
C382 SWP[7] SWP[3] 0.043107f
C383 x2/net7 SWN[0] 0.173771f
C384 x3/COMP_BUF_N SWP[9] 0.228718f
C385 EN DOUT[9] 1.5946f
C386 VDDD SWN[1] 2.72394f
C387 x2/TRIG2 DOUT[8] 0.014937f
C388 CF[4] CF[1] 0.044459f
C389 SWN[5] SWN[6] 0.177435f
C390 CLKS SWN[3] 0.012758f
C391 SWP[4] CF[1] 0.033362f
C392 SWP[5] SWN[1] 0.747975f
C393 CF[0] CF[2] 0.101787f
C394 DOUT[0] DOUT[2] 0.063033f
C395 x2/net3 EN 0.112364f
C396 VDDD SWP[7] 1.16442f
C397 FINAL CF[1] 0.026569f
C398 CLKS CF[4] 0.325599f
C399 SWP[1] CF[4] 0.024758f
C400 clknet_1_0__leaf_CLK CF[1] 0.126129f
C401 SWP[0] SWP[9] 0.042861f
C402 CLKS DOUT[2] 0.043561f
C403 CF[4] CF[8] 0.01535f
C404 SWN[3] DOUT[9] 0.035946f
C405 CKO SWN[1] 0.027956f
C406 clknet_0_CLK CF[1] 0.458088f
C407 CLKS SWN[7] 0.193965f
C408 CLKS SWP[4] 1.97232f
C409 SWP[1] SWP[4] 0.031058f
C410 EN SWN[6] 0.150227f
C411 COMP_N COMP_P 0.433165f
C412 SWP[4] CF[8] 0.023113f
C413 SWP[7] SWP[5] 0.041798f
C414 x3/COMP_BUF_P SWP[8] 0.202291f
C415 FINAL CLKS 0.756376f
C416 clknet_1_0__leaf_CLK CLKS 0.876917f
C417 clknet_1_0__leaf_CLK SWP[1] 0.150001f
C418 x3/COMP_BUF_N SWN[1] 0.047192f
C419 clknet_1_0__leaf_CLK CF[8] 0.128649f
C420 SWN[4] SWN[2] 0.125583f
C421 DOUT[7] SWN[5] 0.128494f
C422 clknet_0_CLK CLKS 0.099932f
C423 clknet_0_CLK SWP[1] 0.019278f
C424 clknet_0_CLK CF[8] 0.015934f
C425 CKO SWP[7] 0.010641f
C426 CF[0] SWP[3] 0.040093f
C427 SWN[8] SWN[7] 0.161017f
C428 x2/net9 SWN[1] 0.051513f
C429 x2/net11 EN 0.179583f
C430 CF[1] CF[9] 0.127123f
C431 SWN[0] SWN[1] 0.463249f
C432 VDDD DOUT[3] 1.25371f
C433 x3/COMP_BUF_P DOUT[6] 0.011864f
C434 clknet_1_1__leaf_CLK DOUT[9] 0.344782f
C435 CF[0] CF[3] 1.37253f
C436 x2/TRIG1 VDDD 0.484796f
C437 EN DOUT[7] 0.791273f
C438 VDDD CF[0] 2.16811f
C439 CLKS CF[9] 0.306593f
C440 SWP[1] CF[9] 0.06501f
C441 CF[1] CF[2] 1.12944f
C442 SWN[6] SWN[7] 0.308281f
C443 CF[9] CF[8] 0.374014f
C444 x2/net12 x2/net13 0.474603f
C445 SWP[6] SWP[3] 0.044662f
C446 CLK SWP[3] 0.019063f
C447 COMP_N DOUT[0] 0.061261f
C448 x2/TRIG2 VDDD 0.535876f
C449 SWP[1] COMP_N 0.046763f
C450 clkload0.X CLKS 0.049202f
C451 clknet_1_1__leaf_CLK x2/net3 0.07351f
C452 SWP[0] SWP[7] 0.049409f
C453 CF[0] CF[7] 0.019135f
C454 x3/COMP_BUF_P CF[6] 0.694709f
C455 DOUT[8] DOUT[9] 0.356538f
C456 CF[0] SWP[5] 0.083255f
C457 SWP[8] SWN[5] 0.021139f
C458 CLKS CF[2] 0.038574f
C459 SWP[1] CF[2] 0.042285f
C460 CF[8] CF[2] 0.024382f
C461 CLKS DOUT[5] 0.153911f
C462 CF[5] CF[4] 0.340043f
C463 CF[3] CLK 0.022117f
C464 SWP[2] CF[4] 0.036131f
C465 SWN[3] DOUT[7] 0.034845f
C466 VDDD SWP[6] 2.11804f
C467 VDDD CLK 0.622641f
C468 CKO CF[0] 0.052657f
C469 VDDD COMP_P 0.999956f
C470 x2/net8 SWN[2] 0.051959f
C471 CF[5] SWP[4] 0.041719f
C472 SWN[5] SWN[4] 0.163342f
C473 SWP[2] SWP[4] 0.052824f
C474 SWP[3] CF[1] 0.132757f
C475 FINAL CF[5] 0.016965f
C476 SWP[6] CF[7] 0.200687f
C477 x2/net13 SWN[1] 0.015124f
C478 x3/COMP_BUF_N CF[0] 0.028307f
C479 clknet_1_0__leaf_CLK SWP[2] 1.47177f
C480 clknet_1_0__leaf_CLK CF[5] 0.752642f
C481 EN SWP[8] 0.614322f
C482 SWP[5] SWP[6] 0.491833f
C483 clknet_1_1__leaf_CLK x2/net11 0.302258f
C484 SWN[7] SWN[9] 0.130328f
C485 CLKS SWP[3] 0.380036f
C486 x2/net3 DOUT[5] 0.03729f
C487 SWP[1] SWP[3] 0.019802f
C488 CKO CLK 0.298934f
C489 CKO SWP[6] 0.083123f
C490 SWP[3] CF[8] 0.024592f
C491 CKO COMP_P 0.30089f
C492 CF[3] CF[1] 0.039958f
C493 x2/net6 VDDD 0.960719f
C494 VDDD CF[1] 1.50883f
C495 EN SWN[4] 0.056712f
C496 clknet_1_1__leaf_CLK DOUT[7] 0.055485f
C497 x2/TRIG2 x2/net7 0.018389f
C498 SWP[0] CF[0] 0.404727f
C499 x2/TRIG2 SWN[0] 0.025291f
C500 EN SWN[2] 0.18966f
C501 x2/net5 x2/net11 0.021886f
C502 x3/COMP_BUF_N SWP[6] 0.191989f
C503 EN DOUT[6] 0.167239f
C504 VDDD DOUT[0] 0.594659f
C505 CF[1] CF[7] 0.015359f
C506 DOUT[4] DOUT[3] 2.2149f
C507 SWP[1] CF[3] 0.024632f
C508 CLKS CF[3] 0.987838f
C509 SWP[5] CF[1] 0.020141f
C510 CF[5] CF[9] 0.027656f
C511 SWP[2] CF[9] 0.019698f
C512 CF[3] CF[8] 0.024572f
C513 VDDD CLKS 11.8564f
C514 VDDD SWP[1] 2.63298f
C515 VDDD CF[8] 4.578f
C516 x3/COMP_BUF_P EN 0.285508f
C517 CLKS CLKSB 0.312614f
C518 SWP[8] SWP[4] 0.048743f
C519 SWN[3] SWN[4] 0.480097f
C520 DOUT[8] DOUT[7] 2.46101f
C521 x2/net11 DOUT[5] 0.024213f
C522 VDDD DOUT[9] 1.63252f
C523 CLKS CF[7] 0.881462f
C524 SWP[1] CF[7] 0.085603f
C525 CF[8] CF[7] 0.329745f
C526 SWP[0] CLK 0.018331f
C527 SWP[0] SWP[6] 0.039648f
C528 SWP[1] SWP[5] 0.025096f
C529 SWP[0] COMP_P 0.065604f
C530 CLKS SWP[5] 0.330238f
C531 CF[5] CF[2] 0.200155f
C532 SWP[5] CF[8] 0.019214f
C533 SWP[2] CF[2] 0.050614f
C534 SWN[3] SWN[2] 0.486898f
C535 VDDD SWN[8] 0.442783f
C536 SWP[9] SWP[6] 0.085052f
C537 CKO SWP[1] 0.085925f
C538 CKO CLKS 0.935833f
C539 x2/net3 VDDD 1.20538f
C540 x2/net2 EN 0.03168f
C541 SWP[4] SWN[2] 0.025013f
C542 DOUT[6] SWP[4] 0.454543f
C543 COMP_P DOUT[4] 0.046075f
C544 x3/COMP_BUF_P CF[4] 0.047913f
C545 CKO DOUT[9] 0.361718f
C546 x2/TRIG1 SWN[1] 0.025457f
C547 x2/net6 SWN[0] 0.035769f
C548 x2/net6 x2/net7 0.109841f
C549 CF[0] SWN[1] 0.216263f
C550 x3/COMP_BUF_N SWP[1] 0.010828f
C551 x3/COMP_BUF_N CLKS 1.55149f
C552 x3/COMP_BUF_N CF[8] 0.452996f
C553 VDDD SWN[6] 1.02098f
C554 x2/net8 EN 0.072432f
C555 x3/COMP_BUF_P SWP[4] 0.262781f
C556 SWP[0] CF[1] 0.046901f
C557 x2/TRIG2 SWN[1] 0.028475f
C558 CF[4] CF[6] 0.902529f
C559 CF[5] SWP[3] 0.061453f
C560 SWP[2] SWP[3] 2.03044f
C561 x3/COMP_BUF_P FINAL 0.031828f
C562 EN SWN[5] 0.463474f
C563 clknet_1_1__leaf_CLK SWN[2] 0.098414f
C564 clknet_1_1__leaf_CLK DOUT[6] 0.015237f
C565 SWP[9] CF[1] 0.053398f
C566 clknet_0_CLK x3/COMP_BUF_P 1.32062f
C567 x2/net6 x2/net12 0.14998f
C568 x2/net9 DOUT[9] 0.030129f
C569 SWP[1] SWP[0] 4.69417f
C570 SWP[0] CLKS 0.405401f
C571 SWP[0] CF[8] 0.083319f
C572 x2/net11 VDDD 2.51174f
C573 clknet_1_0__leaf_CLK CF[6] 0.15192f
C574 SWP[6] SWN[1] 0.031321f
C575 x2/net10 EN 0.272337f
C576 x2/net7 DOUT[9] 0.023015f
C577 DOUT[8] SWN[4] 0.048105f
C578 SWN[0] DOUT[9] 0.1491f
C579 CKO SWN[6] 0.150426f
C580 CF[3] CF[5] 0.043261f
C581 CF[3] SWP[2] 0.091601f
C582 x2/net10 x2/net1 0.015525f
C583 x2/net8 SWN[3] 0.052986f
C584 VDDD CF[5] 4.04704f
C585 VDDD SWP[2] 2.47449f
C586 SWP[1] SWP[9] 0.032644f
C587 CLKS SWP[9] 1.05486f
C588 x2/net5 DOUT[6] 0.048038f
C589 DOUT[1] DOUT[2] 0.33988f
C590 SWP[9] CF[8] 0.036314f
C591 DOUT[8] SWN[2] 0.029632f
C592 VDDD DOUT[7] 0.715152f
C593 x2/net1 EN 0.166882f
C594 CLKS DOUT[4] 0.413541f
C595 clkload0.X DOUT[6] 0.11079f
C596 COMP_N DOUT[6] 0.044231f
C597 CF[5] CF[7] 0.02083f
C598 SWP[2] CF[7] 0.023158f
C599 x3/COMP_BUF_P CF[9] 0.112133f
C600 SWP[7] SWP[6] 0.349701f
C601 CF[5] SWP[5] 0.209199f
C602 SWP[2] SWP[5] 0.047772f
C603 VDDD SWN[9] 0.745797f
C604 SWN[9] VSSD 1.14869f
C605 CF[7] VSSD 5.53496f
C606 SWN[7] VSSD 1.16356f
C607 SWN[2] VSSD 1.83093f
C608 SWN[8] VSSD 1.38987f
C609 CF[2] VSSD 3.73077f
C610 CF[8] VSSD 3.048668f
C611 CF[9] VSSD 3.224304f
C612 CF[1] VSSD 4.63515f
C613 SWN[1] VSSD 4.729379f
C614 CF[6] VSSD 3.41792f
C615 SWN[6] VSSD 1.23244f
C616 DOUT[3] VSSD 3.111028f
C617 SWP[3] VSSD 7.407114f
C618 CLK VSSD 2.77574f
C619 DOUT[4] VSSD 3.113709f
C620 SWP[4] VSSD 4.500352f
C621 DOUT[6] VSSD 4.749067f
C622 SWP[6] VSSD 3.788809f
C623 CF[4] VSSD 3.226725f
C624 SWN[4] VSSD 1.23717f
C625 DOUT[9] VSSD 1.61305f
C626 SWP[9] VSSD 4.05661f
C627 DOUT[5] VSSD 2.89282f
C628 SWN[5] VSSD 2.18352f
C629 DOUT[7] VSSD 4.413061f
C630 COMP_P VSSD 1.69997f
C631 SWP[5] VSSD 3.26489f
C632 CF[5] VSSD 2.977226f
C633 SWP[7] VSSD 4.04492f
C634 CLKSB VSSD 0.993378f
C635 DOUT[2] VSSD 1.61598f
C636 SWP[2] VSSD 7.276391f
C637 CF[3] VSSD 5.184036f
C638 SWN[3] VSSD 4.082685f
C639 CF[0] VSSD 7.498019f
C640 SWN[0] VSSD 1.75901f
C641 DOUT[8] VSSD 3.359154f
C642 SWP[8] VSSD 5.213109f
C643 DOUT[0] VSSD 1.11428f
C644 CLKS VSSD 27.17558f
C645 SWP[0] VSSD 7.841119f
C646 COMP_N VSSD 1.94556f
C647 DOUT[1] VSSD 0.93513f
C648 SWP[1] VSSD 8.039521f
C649 CKO VSSD 7.278111f
C650 EN VSSD 20.513067f
C651 VDDD VSSD 0.458585p
C652 FINAL VSSD 1.560651f
C653 clkload0.X VSSD 0.544346f
C654 clknet_1_0__leaf_CLK VSSD 4.837007f
C655 x3/COMP_BUF_P VSSD 5.464219f
C656 x3/COMP_BUF_N VSSD 6.077292f
C657 x2/net13 VSSD 1.36127f
C658 clknet_0_CLK VSSD 3.660447f
C659 x2/net12 VSSD 0.720534f
C660 x2/net7 VSSD 0.440933f
C661 x2/net6 VSSD 0.79435f
C662 x2/TRIG2 VSSD 2.97343f
C663 x2/net11 VSSD 2.096697f
C664 x2/net5 VSSD 0.512639f
C665 x2/net4 VSSD 0.574721f
C666 x2/net8 VSSD 0.63756f
C667 x2/net3 VSSD 0.463739f
C668 x2/net1 VSSD 0.403119f
C669 x2/net2 VSSD 0.354111f
C670 x2/net9 VSSD 0.36708f
C671 x2/TRIG1 VSSD 0.807423f
C672 x2/net10 VSSD 0.503742f
C673 clknet_1_1__leaf_CLK VSSD 6.15894f
C674 SWN[3].n0 VSSD 0.013612f
C675 SWN[3].n1 VSSD 0.018377f
C676 SWN[3].t1 VSSD 0.010471f
C677 SWN[3].n2 VSSD 0.151096f
C678 SWN[3].t0 VSSD 0.010471f
C679 SWN[3].n3 VSSD 0.020941f
C680 SWP[2].t5 VSSD 0.018879f
C681 SWP[2].t4 VSSD 0.020782f
C682 SWP[2].n0 VSSD 0.058855f
C683 SWP[2].t0 VSSD 0.015031f
C684 SWP[2].t1 VSSD 0.015031f
C685 SWP[2].n1 VSSD 0.030092f
C686 SWP[2].n3 VSSD 0.01954f
C687 SWP[2].n4 VSSD 0.024014f
C688 SWP[2].n6 VSSD 0.700772f
C689 SWP[1].t5 VSSD 0.029387f
C690 SWP[1].t4 VSSD 0.03235f
C691 SWP[1].n0 VSSD 0.091617f
C692 SWP[1].t1 VSSD 0.023397f
C693 SWP[1].t0 VSSD 0.023397f
C694 SWP[1].n1 VSSD 0.046843f
C695 SWP[1].t2 VSSD 0.015208f
C696 SWP[1].t3 VSSD 0.015208f
C697 SWP[1].n3 VSSD 0.030417f
C698 SWP[1].n4 VSSD 0.037381f
C699 SWP[1].n6 VSSD 1.9137f
C700 DOUT[7].n0 VSSD 0.017413f
C701 DOUT[7].n1 VSSD 0.020785f
C702 DOUT[7].t1 VSSD 0.013395f
C703 DOUT[7].t0 VSSD 0.013395f
C704 DOUT[7].n3 VSSD 0.026789f
C705 DOUT[7].n5 VSSD 0.030982f
C706 DOUT[3].n0 VSSD 0.019147f
C707 DOUT[3].n1 VSSD 0.022854f
C708 DOUT[3].t1 VSSD 0.014728f
C709 DOUT[3].t0 VSSD 0.014728f
C710 DOUT[3].n3 VSSD 0.029456f
C711 DOUT[3].n5 VSSD 0.405227f
C712 DOUT[6].n0 VSSD 0.012515f
C713 DOUT[6].n1 VSSD 0.016896f
C714 DOUT[6].n3 VSSD 0.019254f
C715 DOUT[6].n4 VSSD 0.379709f
C716 CF[5].t9 VSSD 0.018173f
C717 CF[5].t6 VSSD 0.027163f
C718 CF[5].n0 VSSD 0.050203f
C719 CF[5].t1 VSSD 0.016734f
C720 CF[5].t0 VSSD 0.016734f
C721 CF[5].t3 VSSD 0.010877f
C722 CF[5].t2 VSSD 0.010877f
C723 CF[5].n1 VSSD 0.021754f
C724 CF[5].n2 VSSD 0.027947f
C725 CF[5].n3 VSSD 0.010536f
C726 CF[5].n4 VSSD 0.033467f
C727 CF[5].n6 VSSD 0.016246f
C728 CF[5].n7 VSSD 0.23529f
C729 CF[5].t8 VSSD 0.021017f
C730 CF[5].t4 VSSD 0.023136f
C731 CF[5].n8 VSSD 0.066164f
C732 CF[5].n9 VSSD 0.066661f
C733 CF[5].n10 VSSD 0.669164f
C734 CF[5].t7 VSSD 0.018173f
C735 CF[5].t5 VSSD 0.027163f
C736 CF[5].n11 VSSD 0.050203f
C737 CF[5].n12 VSSD 0.030659f
C738 CF[5].n13 VSSD 0.970208f
C739 CF[5].n14 VSSD 0.325822f
C740 DOUT[8].n0 VSSD 0.019259f
C741 DOUT[8].n1 VSSD 0.026001f
C742 DOUT[8].t1 VSSD 0.014815f
C743 DOUT[8].n2 VSSD 0.440628f
C744 DOUT[8].t0 VSSD 0.014815f
C745 DOUT[8].n3 VSSD 0.029629f
C746 SWP[4].t5 VSSD 0.010753f
C747 SWP[4].t4 VSSD 0.011837f
C748 SWP[4].n0 VSSD 0.03385f
C749 SWP[4].n2 VSSD 0.017122f
C750 SWP[4].n4 VSSD 0.011129f
C751 SWP[4].n5 VSSD 0.014298f
C752 SWP[4].n6 VSSD 0.603061f
C753 SWP[4].n7 VSSD 0.433906f
C754 SWP[7].t5 VSSD 0.012413f
C755 SWP[7].t4 VSSD 0.013674f
C756 SWP[7].n0 VSSD 0.039159f
C757 SWP[7].n1 VSSD 0.019885f
C758 SWP[7].n3 VSSD 0.012912f
C759 SWP[7].n4 VSSD 0.015868f
C760 SWP[7].n6 VSSD 0.603418f
C761 SWN[1].n0 VSSD 0.015693f
C762 SWN[1].n1 VSSD 0.021186f
C763 SWN[1].t1 VSSD 0.012071f
C764 SWN[1].t0 VSSD 0.012071f
C765 SWN[1].n2 VSSD 0.024167f
C766 SWP[6].t5 VSSD 0.011576f
C767 SWP[6].t4 VSSD 0.012744f
C768 SWP[6].n0 VSSD 0.036443f
C769 SWP[6].n1 VSSD 0.011982f
C770 SWP[6].n2 VSSD 0.016176f
C771 SWP[6].n4 VSSD 0.018434f
C772 SWP[6].n6 VSSD 0.511904f
C773 SWP[6].n7 VSSD 0.272415f
C774 SWP[0].t4 VSSD 0.032557f
C775 SWP[0].t5 VSSD 0.035839f
C776 SWP[0].n0 VSSD 0.10249f
C777 SWP[0].t0 VSSD 0.025921f
C778 SWP[0].t1 VSSD 0.025921f
C779 SWP[0].t2 VSSD 0.016849f
C780 SWP[0].t3 VSSD 0.016849f
C781 SWP[0].n1 VSSD 0.033697f
C782 SWP[0].n2 VSSD 0.04329f
C783 SWP[0].n3 VSSD 0.016321f
C784 SWP[0].n4 VSSD 0.051842f
C785 SWP[0].n5 VSSD 0.01224f
C786 SWP[0].n7 VSSD 1.73651f
C787 SWP[0].n8 VSSD 0.586018f
C788 FINAL.t1 VSSD 0.018311f
C789 FINAL.t3 VSSD 0.018311f
C790 FINAL.n0 VSSD 0.039051f
C791 FINAL.t2 VSSD 0.018311f
C792 FINAL.t4 VSSD 0.018311f
C793 FINAL.n1 VSSD 0.039051f
C794 FINAL.t0 VSSD 0.018311f
C795 FINAL.t5 VSSD 0.018311f
C796 FINAL.n2 VSSD 0.040382f
C797 FINAL.t17 VSSD 0.020081f
C798 FINAL.t19 VSSD 0.013799f
C799 FINAL.n3 VSSD 0.058353f
C800 FINAL.n5 VSSD 0.074806f
C801 FINAL.t16 VSSD 0.013799f
C802 FINAL.t18 VSSD 0.020081f
C803 FINAL.n6 VSSD 0.058353f
C804 FINAL.n7 VSSD 0.014622f
C805 FINAL.n8 VSSD 0.33183f
C806 FINAL.n9 VSSD 0.119081f
C807 FINAL.n10 VSSD 0.07251f
C808 FINAL.n11 VSSD 0.071588f
C809 FINAL.t12 VSSD 0.011902f
C810 FINAL.t14 VSSD 0.011902f
C811 FINAL.n12 VSSD 0.025008f
C812 FINAL.t13 VSSD 0.011902f
C813 FINAL.t15 VSSD 0.011902f
C814 FINAL.n13 VSSD 0.025008f
C815 FINAL.t11 VSSD 0.011902f
C816 FINAL.t8 VSSD 0.011902f
C817 FINAL.n14 VSSD 0.035707f
C818 FINAL.n15 VSSD 0.093193f
C819 FINAL.n16 VSSD 0.055751f
C820 FINAL.t10 VSSD 0.011902f
C821 FINAL.t9 VSSD 0.011902f
C822 FINAL.n17 VSSD 0.025511f
C823 FINAL.n18 VSSD 0.045726f
C824 FINAL.n19 VSSD 0.027202f
C825 FINAL.t7 VSSD 0.018311f
C826 FINAL.t6 VSSD 0.018311f
C827 FINAL.n20 VSSD 0.039051f
C828 x3/COMP_BUF_N.t0 VSSD 0.013983f
C829 x3/COMP_BUF_N.t2 VSSD 0.013983f
C830 x3/COMP_BUF_N.n0 VSSD 0.029821f
C831 x3/COMP_BUF_N.n1 VSSD 0.019097f
C832 x3/COMP_BUF_N.n2 VSSD 0.019097f
C833 x3/COMP_BUF_N.n3 VSSD 0.027267f
C834 x3/COMP_BUF_N.n4 VSSD 0.071165f
C835 x3/COMP_BUF_N.n5 VSSD 0.042573f
C836 x3/COMP_BUF_N.n6 VSSD 0.019481f
C837 x3/COMP_BUF_N.n7 VSSD 0.034918f
C838 x3/COMP_BUF_N.t6 VSSD 0.013983f
C839 x3/COMP_BUF_N.t3 VSSD 0.013983f
C840 x3/COMP_BUF_N.n8 VSSD 0.029821f
C841 x3/COMP_BUF_N.t1 VSSD 0.013983f
C842 x3/COMP_BUF_N.t5 VSSD 0.013983f
C843 x3/COMP_BUF_N.n9 VSSD 0.030837f
C844 x3/COMP_BUF_N.t32 VSSD 0.017476f
C845 x3/COMP_BUF_N.t31 VSSD 0.01925f
C846 x3/COMP_BUF_N.n10 VSSD 0.055129f
C847 x3/COMP_BUF_N.t23 VSSD 0.017476f
C848 x3/COMP_BUF_N.t28 VSSD 0.01925f
C849 x3/COMP_BUF_N.n11 VSSD 0.05486f
C850 x3/COMP_BUF_N.t34 VSSD 0.017476f
C851 x3/COMP_BUF_N.t33 VSSD 0.01925f
C852 x3/COMP_BUF_N.n12 VSSD 0.054948f
C853 x3/COMP_BUF_N.n13 VSSD 0.067706f
C854 x3/COMP_BUF_N.n14 VSSD 0.252147f
C855 x3/COMP_BUF_N.t25 VSSD 0.017476f
C856 x3/COMP_BUF_N.t21 VSSD 0.01925f
C857 x3/COMP_BUF_N.n15 VSSD 0.054948f
C858 x3/COMP_BUF_N.n16 VSSD 0.094223f
C859 x3/COMP_BUF_N.t35 VSSD 0.017476f
C860 x3/COMP_BUF_N.t22 VSSD 0.01925f
C861 x3/COMP_BUF_N.n17 VSSD 0.055129f
C862 x3/COMP_BUF_N.t16 VSSD 0.017476f
C863 x3/COMP_BUF_N.t29 VSSD 0.01925f
C864 x3/COMP_BUF_N.n18 VSSD 0.054948f
C865 x3/COMP_BUF_N.n19 VSSD 0.076482f
C866 x3/COMP_BUF_N.t27 VSSD 0.017476f
C867 x3/COMP_BUF_N.t26 VSSD 0.01925f
C868 x3/COMP_BUF_N.n20 VSSD 0.055129f
C869 x3/COMP_BUF_N.n21 VSSD 0.451968f
C870 x3/COMP_BUF_N.n22 VSSD 0.140827f
C871 x3/COMP_BUF_N.n23 VSSD 0.264362f
C872 x3/COMP_BUF_N.t18 VSSD 0.017476f
C873 x3/COMP_BUF_N.t17 VSSD 0.01925f
C874 x3/COMP_BUF_N.n24 VSSD 0.05486f
C875 x3/COMP_BUF_N.n25 VSSD 0.178933f
C876 x3/COMP_BUF_N.n26 VSSD 0.142238f
C877 x3/COMP_BUF_N.t20 VSSD 0.017476f
C878 x3/COMP_BUF_N.t30 VSSD 0.01925f
C879 x3/COMP_BUF_N.n27 VSSD 0.05486f
C880 x3/COMP_BUF_N.n28 VSSD 0.291269f
C881 x3/COMP_BUF_N.n29 VSSD 0.383689f
C882 x3/COMP_BUF_N.t19 VSSD 0.017476f
C883 x3/COMP_BUF_N.t24 VSSD 0.01925f
C884 x3/COMP_BUF_N.n30 VSSD 0.055129f
C885 x3/COMP_BUF_N.n31 VSSD 0.179767f
C886 x3/COMP_BUF_N.n32 VSSD 0.055605f
C887 x3/COMP_BUF_N.t7 VSSD 0.013983f
C888 x3/COMP_BUF_N.t4 VSSD 0.013983f
C889 x3/COMP_BUF_N.n33 VSSD 0.029821f
C890 x3/COMP_BUF_N.n34 VSSD 0.055371f
C891 x3/COMP_BUF_N.n35 VSSD 0.054667f
C892 x3/COMP_BUF_N.n36 VSSD 0.020772f
C893 CKO.t9 VSSD 0.020089f
C894 CKO.t21 VSSD 0.030026f
C895 CKO.n0 VSSD 0.055495f
C896 CKO.n1 VSSD 0.017125f
C897 CKO.t23 VSSD 0.030026f
C898 CKO.t11 VSSD 0.020089f
C899 CKO.n2 VSSD 0.054869f
C900 CKO.n4 VSSD 0.063929f
C901 CKO.t10 VSSD 0.020089f
C902 CKO.t22 VSSD 0.030026f
C903 CKO.n5 VSSD 0.055495f
C904 CKO.n6 VSSD 0.016305f
C905 CKO.n7 VSSD 0.269074f
C906 CKO.t16 VSSD 0.030026f
C907 CKO.t5 VSSD 0.020089f
C908 CKO.n8 VSSD 0.054869f
C909 CKO.n9 VSSD 0.016305f
C910 CKO.n10 VSSD 0.267522f
C911 CKO.t12 VSSD 0.020089f
C912 CKO.t4 VSSD 0.030026f
C913 CKO.n11 VSSD 0.055495f
C914 CKO.n12 VSSD 0.01915f
C915 CKO.t20 VSSD 0.030026f
C916 CKO.t6 VSSD 0.020089f
C917 CKO.n13 VSSD 0.054869f
C918 CKO.n15 VSSD 0.078668f
C919 CKO.t19 VSSD 0.020089f
C920 CKO.t13 VSSD 0.030026f
C921 CKO.n16 VSSD 0.055495f
C922 CKO.n17 VSSD 0.016305f
C923 CKO.n18 VSSD 0.212354f
C924 CKO.t8 VSSD 0.030026f
C925 CKO.t15 VSSD 0.020089f
C926 CKO.n19 VSSD 0.054869f
C927 CKO.n20 VSSD 0.016305f
C928 CKO.n21 VSSD 0.368072f
C929 CKO.t18 VSSD 0.030026f
C930 CKO.t7 VSSD 0.020089f
C931 CKO.n22 VSSD 0.054869f
C932 CKO.n24 VSSD 0.055697f
C933 CKO.n25 VSSD 0.377716f
C934 CKO.n26 VSSD 0.38534f
C935 CKO.n27 VSSD 0.278857f
C936 CKO.t14 VSSD 0.030026f
C937 CKO.t17 VSSD 0.020089f
C938 CKO.n28 VSSD 0.054869f
C939 CKO.n30 VSSD 0.041416f
C940 CKO.n31 VSSD 0.211876f
C941 CKO.n32 VSSD 0.123306f
C942 CKO.t2 VSSD 0.045244f
C943 CKO.n33 VSSD 0.014168f
C944 CKO.n34 VSSD 0.016072f
C945 CKO.t0 VSSD 0.0322f
C946 CKO.n35 VSSD 0.098009f
C947 CKO.n36 VSSD 0.018594f
C948 CKO.n37 VSSD 0.034318f
C949 CKO.t1 VSSD 0.0322f
C950 CKO.n38 VSSD 0.098116f
C951 CKO.t3 VSSD 0.045244f
C952 CKO.n39 VSSD 0.025753f
C953 CKO.n40 VSSD 0.018004f
C954 CKO.n41 VSSD 0.013236f
C955 CKO.n42 VSSD 0.065103f
C956 CKO.n43 VSSD 0.38365f
C957 SWP[8].t4 VSSD 0.023052f
C958 SWP[8].t5 VSSD 0.025391f
C959 SWP[8].n0 VSSD 0.072362f
C960 SWP[8].t1 VSSD 0.018444f
C961 SWP[8].t0 VSSD 0.018444f
C962 SWP[8].t2 VSSD 0.011989f
C963 SWP[8].t3 VSSD 0.011989f
C964 SWP[8].n1 VSSD 0.023977f
C965 SWP[8].n2 VSSD 0.030803f
C966 SWP[8].n3 VSSD 0.011613f
C967 SWP[8].n4 VSSD 0.036888f
C968 SWP[8].n6 VSSD 0.115073f
C969 SWP[8].n7 VSSD 1.43153f
C970 CF[3].t6 VSSD 0.017704f
C971 CF[3].t8 VSSD 0.011845f
C972 CF[3].n0 VSSD 0.032352f
C973 CF[3].n2 VSSD 0.214654f
C974 CF[3].t7 VSSD 0.011845f
C975 CF[3].t5 VSSD 0.017704f
C976 CF[3].n3 VSSD 0.032721f
C977 CF[3].n4 VSSD 0.090857f
C978 CF[3].n5 VSSD 0.623344f
C979 CF[3].t4 VSSD 0.013631f
C980 CF[3].t9 VSSD 0.015015f
C981 CF[3].n6 VSSD 0.042859f
C982 CF[3].n7 VSSD 0.048066f
C983 CF[3].n8 VSSD 0.25894f
C984 CF[3].t1 VSSD 0.010907f
C985 CF[3].t2 VSSD 0.010907f
C986 CF[3].n10 VSSD 0.021813f
C987 CF[3].n12 VSSD 0.014179f
C988 CF[3].n13 VSSD 0.018215f
C989 CF[3].n14 VSSD 0.24377f
C990 x3/COMP_BUF_P.t5 VSSD 0.018765f
C991 x3/COMP_BUF_P.t2 VSSD 0.018765f
C992 x3/COMP_BUF_P.n0 VSSD 0.04002f
C993 x3/COMP_BUF_P.t6 VSSD 0.018765f
C994 x3/COMP_BUF_P.t0 VSSD 0.018765f
C995 x3/COMP_BUF_P.n1 VSSD 0.04002f
C996 x3/COMP_BUF_P.t4 VSSD 0.018765f
C997 x3/COMP_BUF_P.t3 VSSD 0.018765f
C998 x3/COMP_BUF_P.n2 VSSD 0.050402f
C999 x3/COMP_BUF_P.n3 VSSD 0.128547f
C1000 x3/COMP_BUF_P.n4 VSSD 0.073363f
C1001 x3/COMP_BUF_P.t8 VSSD 0.012197f
C1002 x3/COMP_BUF_P.t13 VSSD 0.012197f
C1003 x3/COMP_BUF_P.n5 VSSD 0.025628f
C1004 x3/COMP_BUF_P.t9 VSSD 0.012197f
C1005 x3/COMP_BUF_P.t11 VSSD 0.012197f
C1006 x3/COMP_BUF_P.n6 VSSD 0.025628f
C1007 x3/COMP_BUF_P.t15 VSSD 0.012197f
C1008 x3/COMP_BUF_P.t14 VSSD 0.012197f
C1009 x3/COMP_BUF_P.n7 VSSD 0.036592f
C1010 x3/COMP_BUF_P.n8 VSSD 0.095505f
C1011 x3/COMP_BUF_P.n9 VSSD 0.057133f
C1012 x3/COMP_BUF_P.t10 VSSD 0.012197f
C1013 x3/COMP_BUF_P.t12 VSSD 0.012197f
C1014 x3/COMP_BUF_P.n10 VSSD 0.026144f
C1015 x3/COMP_BUF_P.n11 VSSD 0.04686f
C1016 x3/COMP_BUF_P.t19 VSSD 0.023569f
C1017 x3/COMP_BUF_P.t30 VSSD 0.025945f
C1018 x3/COMP_BUF_P.n12 VSSD 0.073598f
C1019 x3/COMP_BUF_P.n13 VSSD 0.095978f
C1020 x3/COMP_BUF_P.t20 VSSD 0.023453f
C1021 x3/COMP_BUF_P.t32 VSSD 0.025834f
C1022 x3/COMP_BUF_P.n14 VSSD 0.073983f
C1023 x3/COMP_BUF_P.t22 VSSD 0.023453f
C1024 x3/COMP_BUF_P.t21 VSSD 0.025834f
C1025 x3/COMP_BUF_P.n15 VSSD 0.073983f
C1026 x3/COMP_BUF_P.n16 VSSD 0.344166f
C1027 x3/COMP_BUF_P.t16 VSSD 0.023453f
C1028 x3/COMP_BUF_P.t25 VSSD 0.025834f
C1029 x3/COMP_BUF_P.n17 VSSD 0.073983f
C1030 x3/COMP_BUF_P.t28 VSSD 0.023569f
C1031 x3/COMP_BUF_P.t35 VSSD 0.025945f
C1032 x3/COMP_BUF_P.n18 VSSD 0.073598f
C1033 x3/COMP_BUF_P.n19 VSSD 0.089612f
C1034 x3/COMP_BUF_P.n20 VSSD 0.567733f
C1035 x3/COMP_BUF_P.n21 VSSD 0.229123f
C1036 x3/COMP_BUF_P.t27 VSSD 0.023453f
C1037 x3/COMP_BUF_P.t26 VSSD 0.025834f
C1038 x3/COMP_BUF_P.n22 VSSD 0.073983f
C1039 x3/COMP_BUF_P.n23 VSSD 0.276122f
C1040 x3/COMP_BUF_P.t18 VSSD 0.023569f
C1041 x3/COMP_BUF_P.t31 VSSD 0.025945f
C1042 x3/COMP_BUF_P.n24 VSSD 0.074553f
C1043 x3/COMP_BUF_P.n25 VSSD 0.139186f
C1044 x3/COMP_BUF_P.n26 VSSD 0.287206f
C1045 x3/COMP_BUF_P.n27 VSSD 0.357688f
C1046 x3/COMP_BUF_P.t33 VSSD 0.023569f
C1047 x3/COMP_BUF_P.t17 VSSD 0.025945f
C1048 x3/COMP_BUF_P.n28 VSSD 0.073478f
C1049 x3/COMP_BUF_P.t24 VSSD 0.023453f
C1050 x3/COMP_BUF_P.t23 VSSD 0.025834f
C1051 x3/COMP_BUF_P.n29 VSSD 0.073622f
C1052 x3/COMP_BUF_P.n30 VSSD 0.465175f
C1053 x3/COMP_BUF_P.t29 VSSD 0.023569f
C1054 x3/COMP_BUF_P.t34 VSSD 0.025945f
C1055 x3/COMP_BUF_P.n31 VSSD 0.073598f
C1056 x3/COMP_BUF_P.n32 VSSD 0.075622f
C1057 x3/COMP_BUF_P.n33 VSSD 0.305405f
C1058 x3/COMP_BUF_P.t7 VSSD 0.018765f
C1059 x3/COMP_BUF_P.t1 VSSD 0.018765f
C1060 x3/COMP_BUF_P.n34 VSSD 0.04002f
C1061 DOUT[4].t0 VSSD 0.015356f
C1062 DOUT[4].t1 VSSD 0.015356f
C1063 DOUT[4].n0 VSSD 0.019962f
C1064 DOUT[4].n1 VSSD 0.02695f
C1065 DOUT[4].n3 VSSD 0.030711f
C1066 DOUT[4].n4 VSSD 0.365275f
C1067 SWP[3].t5 VSSD 0.021478f
C1068 SWP[3].t4 VSSD 0.023643f
C1069 SWP[3].n0 VSSD 0.067614f
C1070 SWP[3].n1 VSSD 0.331727f
C1071 SWP[3].t0 VSSD 0.0171f
C1072 SWP[3].t1 VSSD 0.0171f
C1073 SWP[3].t3 VSSD 0.011115f
C1074 SWP[3].t2 VSSD 0.011115f
C1075 SWP[3].n2 VSSD 0.02223f
C1076 SWP[3].n3 VSSD 0.028559f
C1077 SWP[3].n4 VSSD 0.010767f
C1078 SWP[3].n5 VSSD 0.034201f
C1079 SWP[3].n8 VSSD 0.493402f
C1080 clknet_1_0__leaf_CLK.n0 VSSD 0.021098f
C1081 clknet_1_0__leaf_CLK.n1 VSSD 0.024953f
C1082 clknet_1_0__leaf_CLK.n2 VSSD 0.018177f
C1083 clknet_1_0__leaf_CLK.n3 VSSD 0.011686f
C1084 clknet_1_0__leaf_CLK.n4 VSSD 0.073839f
C1085 clknet_1_0__leaf_CLK.n5 VSSD 0.011686f
C1086 clknet_1_0__leaf_CLK.n6 VSSD 0.044383f
C1087 clknet_1_0__leaf_CLK.n7 VSSD 0.011693f
C1088 clknet_1_0__leaf_CLK.n8 VSSD 0.045782f
C1089 clknet_1_0__leaf_CLK.n9 VSSD 0.011686f
C1090 clknet_1_0__leaf_CLK.n10 VSSD 0.044383f
C1091 clknet_1_0__leaf_CLK.n11 VSSD 0.011686f
C1092 clknet_1_0__leaf_CLK.n12 VSSD 0.044605f
C1093 clknet_1_0__leaf_CLK.n13 VSSD 0.011686f
C1094 clknet_1_0__leaf_CLK.n14 VSSD 0.038315f
C1095 clknet_1_0__leaf_CLK.n15 VSSD 0.011375f
C1096 clknet_1_0__leaf_CLK.t53 VSSD 0.012764f
C1097 clknet_1_0__leaf_CLK.t47 VSSD 0.019077f
C1098 clknet_1_0__leaf_CLK.n16 VSSD 0.035259f
C1099 clknet_1_0__leaf_CLK.n17 VSSD 0.0112f
C1100 clknet_1_0__leaf_CLK.t39 VSSD 0.017172f
C1101 clknet_1_0__leaf_CLK.t36 VSSD 0.017172f
C1102 clknet_1_0__leaf_CLK.n18 VSSD 0.039201f
C1103 clknet_1_0__leaf_CLK.n19 VSSD 0.062882f
C1104 clknet_1_0__leaf_CLK.n20 VSSD 0.077368f
C1105 clknet_1_0__leaf_CLK.t40 VSSD 0.019077f
C1106 clknet_1_0__leaf_CLK.t41 VSSD 0.012764f
C1107 clknet_1_0__leaf_CLK.n21 VSSD 0.034861f
C1108 clknet_1_0__leaf_CLK.n22 VSSD 0.24247f
C1109 clknet_1_0__leaf_CLK.t54 VSSD 0.012764f
C1110 clknet_1_0__leaf_CLK.t44 VSSD 0.019077f
C1111 clknet_1_0__leaf_CLK.n23 VSSD 0.035259f
C1112 clknet_1_0__leaf_CLK.n24 VSSD 0.015083f
C1113 clknet_1_0__leaf_CLK.n25 VSSD 0.08275f
C1114 clknet_1_0__leaf_CLK.t37 VSSD 0.019077f
C1115 clknet_1_0__leaf_CLK.t43 VSSD 0.012764f
C1116 clknet_1_0__leaf_CLK.n26 VSSD 0.034861f
C1117 clknet_1_0__leaf_CLK.n27 VSSD 0.101329f
C1118 clknet_1_0__leaf_CLK.t46 VSSD 0.019077f
C1119 clknet_1_0__leaf_CLK.t32 VSSD 0.012764f
C1120 clknet_1_0__leaf_CLK.n28 VSSD 0.034861f
C1121 clknet_1_0__leaf_CLK.n29 VSSD 0.01036f
C1122 clknet_1_0__leaf_CLK.t49 VSSD 0.019077f
C1123 clknet_1_0__leaf_CLK.t33 VSSD 0.012764f
C1124 clknet_1_0__leaf_CLK.n30 VSSD 0.034861f
C1125 clknet_1_0__leaf_CLK.n31 VSSD 0.01036f
C1126 clknet_1_0__leaf_CLK.t50 VSSD 0.019077f
C1127 clknet_1_0__leaf_CLK.t34 VSSD 0.012764f
C1128 clknet_1_0__leaf_CLK.n32 VSSD 0.034861f
C1129 clknet_1_0__leaf_CLK.n33 VSSD 0.01036f
C1130 clknet_1_0__leaf_CLK.t35 VSSD 0.012764f
C1131 clknet_1_0__leaf_CLK.t55 VSSD 0.019077f
C1132 clknet_1_0__leaf_CLK.n34 VSSD 0.034949f
C1133 clknet_1_0__leaf_CLK.n35 VSSD 0.034805f
C1134 clknet_1_0__leaf_CLK.t52 VSSD 0.012764f
C1135 clknet_1_0__leaf_CLK.t45 VSSD 0.019077f
C1136 clknet_1_0__leaf_CLK.n36 VSSD 0.034949f
C1137 clknet_1_0__leaf_CLK.n37 VSSD 0.015604f
C1138 clknet_1_0__leaf_CLK.n38 VSSD 0.15533f
C1139 clknet_1_0__leaf_CLK.n39 VSSD 0.207604f
C1140 clknet_1_0__leaf_CLK.n40 VSSD 0.09593f
C1141 clknet_1_0__leaf_CLK.t42 VSSD 0.012764f
C1142 clknet_1_0__leaf_CLK.t38 VSSD 0.019077f
C1143 clknet_1_0__leaf_CLK.n41 VSSD 0.035259f
C1144 clknet_1_0__leaf_CLK.n42 VSSD 0.015083f
C1145 clknet_1_0__leaf_CLK.n43 VSSD 0.130909f
C1146 clknet_1_0__leaf_CLK.n44 VSSD 0.107315f
C1147 clknet_1_0__leaf_CLK.n45 VSSD 0.106923f
C1148 clknet_1_0__leaf_CLK.t17 VSSD 0.012188f
C1149 clknet_1_0__leaf_CLK.t24 VSSD 0.012188f
C1150 clknet_1_0__leaf_CLK.n46 VSSD 0.024376f
C1151 clknet_1_0__leaf_CLK.n47 VSSD 0.017589f
C1152 clknet_1_0__leaf_CLK.t29 VSSD 0.012188f
C1153 clknet_1_0__leaf_CLK.t1 VSSD 0.012188f
C1154 clknet_1_0__leaf_CLK.n48 VSSD 0.02569f
C1155 clknet_1_0__leaf_CLK.t26 VSSD 0.012188f
C1156 clknet_1_0__leaf_CLK.t31 VSSD 0.012188f
C1157 clknet_1_0__leaf_CLK.n49 VSSD 0.02569f
C1158 clknet_1_0__leaf_CLK.t12 VSSD 0.012188f
C1159 clknet_1_0__leaf_CLK.t8 VSSD 0.012188f
C1160 clknet_1_0__leaf_CLK.n50 VSSD 0.03096f
C1161 clknet_1_0__leaf_CLK.t21 VSSD 0.012188f
C1162 clknet_1_0__leaf_CLK.t15 VSSD 0.012188f
C1163 clknet_1_0__leaf_CLK.n51 VSSD 0.02569f
C1164 clknet_1_0__leaf_CLK.n52 VSSD 0.117079f
C1165 clknet_1_0__leaf_CLK.t13 VSSD 0.012188f
C1166 clknet_1_0__leaf_CLK.t11 VSSD 0.012188f
C1167 clknet_1_0__leaf_CLK.n53 VSSD 0.02569f
C1168 clknet_1_0__leaf_CLK.n54 VSSD 0.067442f
C1169 clknet_1_0__leaf_CLK.t3 VSSD 0.012188f
C1170 clknet_1_0__leaf_CLK.t0 VSSD 0.012188f
C1171 clknet_1_0__leaf_CLK.n55 VSSD 0.02569f
C1172 clknet_1_0__leaf_CLK.n56 VSSD 0.067129f
C1173 clknet_1_0__leaf_CLK.n57 VSSD 0.067129f
C1174 clknet_1_0__leaf_CLK.n58 VSSD 0.067442f
C1175 clknet_1_0__leaf_CLK.n59 VSSD 0.031316f
C1176 clknet_1_0__leaf_CLK.t10 VSSD 0.012188f
C1177 clknet_1_0__leaf_CLK.t19 VSSD 0.012188f
C1178 clknet_1_0__leaf_CLK.n60 VSSD 0.025335f
C1179 x2/net11.t3 VSSD 0.02245f
C1180 x2/net11.t2 VSSD 0.02245f
C1181 x2/net11.n0 VSSD 0.044899f
C1182 x2/net11.n1 VSSD 0.060617f
C1183 x2/net11.t0 VSSD 0.034538f
C1184 x2/net11.t1 VSSD 0.034538f
C1185 x2/net11.t5 VSSD 0.035731f
C1186 x2/net11.t4 VSSD 0.057213f
C1187 x2/net11.n2 VSSD 0.107196f
C1188 x2/net11.n3 VSSD 0.03182f
C1189 x2/net11.n4 VSSD 0.726032f
C1190 x2/net11.n5 VSSD 0.069076f
C1191 x2/net11.n6 VSSD 0.021746f
C1192 clknet_0_CLK.n0 VSSD 0.015649f
C1193 clknet_0_CLK.n1 VSSD 0.010061f
C1194 clknet_0_CLK.n2 VSSD 0.063572f
C1195 clknet_0_CLK.n3 VSSD 0.010061f
C1196 clknet_0_CLK.n4 VSSD 0.038211f
C1197 clknet_0_CLK.n5 VSSD 0.010067f
C1198 clknet_0_CLK.n6 VSSD 0.039416f
C1199 clknet_0_CLK.n7 VSSD 0.010061f
C1200 clknet_0_CLK.n8 VSSD 0.038211f
C1201 clknet_0_CLK.t40 VSSD 0.014784f
C1202 clknet_0_CLK.t33 VSSD 0.014784f
C1203 clknet_0_CLK.t45 VSSD 0.014784f
C1204 clknet_0_CLK.t34 VSSD 0.014784f
C1205 clknet_0_CLK.n10 VSSD 0.033751f
C1206 clknet_0_CLK.n11 VSSD 0.044454f
C1207 clknet_0_CLK.n12 VSSD 0.044454f
C1208 clknet_0_CLK.n13 VSSD 0.054138f
C1209 clknet_0_CLK.n14 VSSD 0.103343f
C1210 clknet_0_CLK.t35 VSSD 0.014784f
C1211 clknet_0_CLK.t36 VSSD 0.014784f
C1212 clknet_0_CLK.t37 VSSD 0.014784f
C1213 clknet_0_CLK.t39 VSSD 0.014784f
C1214 clknet_0_CLK.n15 VSSD 0.033751f
C1215 clknet_0_CLK.n16 VSSD 0.044454f
C1216 clknet_0_CLK.n17 VSSD 0.044454f
C1217 clknet_0_CLK.n18 VSSD 0.053991f
C1218 clknet_0_CLK.n19 VSSD 0.010336f
C1219 clknet_0_CLK.n20 VSSD 0.463294f
C1220 clknet_0_CLK.n21 VSSD 0.015024f
C1221 clknet_0_CLK.n22 VSSD 0.024644f
C1222 clknet_0_CLK.n23 VSSD 0.010061f
C1223 clknet_0_CLK.n24 VSSD 0.032987f
C1224 clknet_0_CLK.n26 VSSD 0.043864f
C1225 clknet_0_CLK.t11 VSSD 0.010493f
C1226 clknet_0_CLK.t0 VSSD 0.010493f
C1227 clknet_0_CLK.n27 VSSD 0.022118f
C1228 clknet_0_CLK.t12 VSSD 0.010493f
C1229 clknet_0_CLK.t13 VSSD 0.010493f
C1230 clknet_0_CLK.n28 VSSD 0.022118f
C1231 clknet_0_CLK.t1 VSSD 0.010493f
C1232 clknet_0_CLK.t4 VSSD 0.010493f
C1233 clknet_0_CLK.n29 VSSD 0.026655f
C1234 clknet_0_CLK.t6 VSSD 0.010493f
C1235 clknet_0_CLK.t8 VSSD 0.010493f
C1236 clknet_0_CLK.n30 VSSD 0.022118f
C1237 clknet_0_CLK.n31 VSSD 0.100799f
C1238 clknet_0_CLK.t10 VSSD 0.010493f
C1239 clknet_0_CLK.t5 VSSD 0.010493f
C1240 clknet_0_CLK.n32 VSSD 0.022118f
C1241 clknet_0_CLK.n33 VSSD 0.058065f
C1242 clknet_0_CLK.t7 VSSD 0.010493f
C1243 clknet_0_CLK.t9 VSSD 0.010493f
C1244 clknet_0_CLK.n34 VSSD 0.022118f
C1245 clknet_0_CLK.n35 VSSD 0.057795f
C1246 clknet_0_CLK.t14 VSSD 0.010493f
C1247 clknet_0_CLK.t15 VSSD 0.010493f
C1248 clknet_0_CLK.n36 VSSD 0.022118f
C1249 clknet_0_CLK.n37 VSSD 0.057795f
C1250 clknet_0_CLK.n38 VSSD 0.058065f
C1251 clknet_0_CLK.n39 VSSD 0.050039f
C1252 clknet_0_CLK.t2 VSSD 0.010493f
C1253 clknet_0_CLK.t3 VSSD 0.010493f
C1254 clknet_0_CLK.n40 VSSD 0.021812f
C1255 CF[9].t1 VSSD 0.016871f
C1256 CF[9].t0 VSSD 0.016871f
C1257 CF[9].n0 VSSD 0.033777f
C1258 CF[9].n1 VSSD 0.010623f
C1259 CF[9].t2 VSSD 0.010966f
C1260 CF[9].t3 VSSD 0.010966f
C1261 CF[9].n2 VSSD 0.021933f
C1262 CF[9].n3 VSSD 0.026955f
C1263 CF[9].n4 VSSD 0.016284f
C1264 CF[9].t7 VSSD 0.018323f
C1265 CF[9].t5 VSSD 0.027386f
C1266 CF[9].n5 VSSD 0.05017f
C1267 CF[9].n6 VSSD 0.13282f
C1268 CF[9].t4 VSSD 0.027386f
C1269 CF[9].t8 VSSD 0.018323f
C1270 CF[9].n7 VSSD 0.050044f
C1271 CF[9].n8 VSSD 0.014872f
C1272 CF[9].n9 VSSD 0.553394f
C1273 CF[9].t9 VSSD 0.02119f
C1274 CF[9].t6 VSSD 0.023326f
C1275 CF[9].n10 VSSD 0.066708f
C1276 CF[9].n11 VSSD 0.067209f
C1277 CF[9].n12 VSSD 0.599106f
C1278 CF[9].n13 VSSD 0.167943f
C1279 CF[8].t2 VSSD 0.021803f
C1280 CF[8].t3 VSSD 0.021803f
C1281 CF[8].t0 VSSD 0.014172f
C1282 CF[8].t1 VSSD 0.014172f
C1283 CF[8].n0 VSSD 0.028344f
C1284 CF[8].n1 VSSD 0.036413f
C1285 CF[8].n2 VSSD 0.013728f
C1286 CF[8].n3 VSSD 0.043607f
C1287 CF[8].n4 VSSD 0.010296f
C1288 CF[8].t5 VSSD 0.023679f
C1289 CF[8].t9 VSSD 0.035392f
C1290 CF[8].n6 VSSD 0.064836f
C1291 CF[8].n7 VSSD 0.12389f
C1292 CF[8].t4 VSSD 0.023679f
C1293 CF[8].t7 VSSD 0.035392f
C1294 CF[8].n8 VSSD 0.065412f
C1295 CF[8].n9 VSSD 0.064038f
C1296 CF[8].n10 VSSD 1.04821f
C1297 CF[8].t6 VSSD 0.027385f
C1298 CF[8].t8 VSSD 0.030146f
C1299 CF[8].n11 VSSD 0.086209f
C1300 CF[8].n12 VSSD 0.086857f
C1301 CF[8].n13 VSSD 0.964449f
C1302 CF[8].n14 VSSD 0.309545f
C1303 CF[4].t1 VSSD 0.011346f
C1304 CF[4].t3 VSSD 0.011346f
C1305 CF[4].n0 VSSD 0.022716f
C1306 CF[4].n2 VSSD 0.01475f
C1307 CF[4].n3 VSSD 0.018128f
C1308 CF[4].n4 VSSD 0.013629f
C1309 CF[4].t6 VSSD 0.018418f
C1310 CF[4].t8 VSSD 0.012323f
C1311 CF[4].n5 VSSD 0.033656f
C1312 CF[4].n7 VSSD 0.258172f
C1313 CF[4].t5 VSSD 0.012323f
C1314 CF[4].t4 VSSD 0.018418f
C1315 CF[4].n8 VSSD 0.033741f
C1316 CF[4].n9 VSSD 0.015065f
C1317 CF[4].n10 VSSD 0.223351f
C1318 CF[4].t9 VSSD 0.014251f
C1319 CF[4].t7 VSSD 0.015688f
C1320 CF[4].n11 VSSD 0.044863f
C1321 CF[4].n12 VSSD 0.0452f
C1322 CF[4].n13 VSSD 0.351016f
C1323 CF[4].n14 VSSD 0.177456f
C1324 CF[6].t0 VSSD 0.011787f
C1325 CF[6].t1 VSSD 0.011787f
C1326 CF[6].n0 VSSD 0.015324f
C1327 CF[6].n1 VSSD 0.019686f
C1328 CF[6].n3 VSSD 0.023575f
C1329 CF[6].t7 VSSD 0.019134f
C1330 CF[6].t9 VSSD 0.012802f
C1331 CF[6].n6 VSSD 0.034965f
C1332 CF[6].n7 VSSD 0.01039f
C1333 CF[6].t5 VSSD 0.019134f
C1334 CF[6].t6 VSSD 0.012802f
C1335 CF[6].n8 VSSD 0.034965f
C1336 CF[6].n10 VSSD 0.122592f
C1337 CF[6].n11 VSSD 0.611504f
C1338 CF[6].t4 VSSD 0.014805f
C1339 CF[6].t8 VSSD 0.016298f
C1340 CF[6].n12 VSSD 0.046607f
C1341 CF[6].n13 VSSD 0.046957f
C1342 CF[6].n14 VSSD 0.382457f
C1343 CF[6].n15 VSSD 0.194739f
C1344 EN.t11 VSSD 0.010639f
C1345 EN.n4 VSSD 0.020752f
C1346 EN.n5 VSSD 0.010998f
C1347 EN.n7 VSSD 0.024943f
C1348 EN.t48 VSSD 0.012222f
C1349 EN.n8 VSSD 0.021702f
C1350 EN.n9 VSSD 0.027895f
C1351 EN.t60 VSSD 0.012222f
C1352 EN.n11 VSSD 0.021702f
C1353 EN.n12 VSSD 0.029635f
C1354 EN.t32 VSSD 0.010639f
C1355 EN.n14 VSSD 0.020752f
C1356 EN.n15 VSSD 0.010998f
C1357 EN.n17 VSSD 0.016143f
C1358 EN.t2 VSSD 0.010639f
C1359 EN.n22 VSSD 0.020752f
C1360 EN.n23 VSSD 0.010998f
C1361 EN.n25 VSSD 0.029635f
C1362 EN.t73 VSSD 0.012222f
C1363 EN.n26 VSSD 0.020964f
C1364 EN.n27 VSSD 0.016978f
C1365 EN.n31 VSSD 0.016143f
C1366 EN.t5 VSSD 0.010639f
C1367 EN.n34 VSSD 0.020752f
C1368 EN.n35 VSSD 0.010998f
C1369 EN.n37 VSSD 0.029635f
C1370 EN.t75 VSSD 0.012222f
C1371 EN.n38 VSSD 0.020964f
C1372 EN.n39 VSSD 0.016978f
C1373 EN.n43 VSSD 0.070141f
C1374 EN.t14 VSSD 0.012222f
C1375 EN.n44 VSSD 0.021702f
C1376 EN.n45 VSSD 0.027895f
C1377 EN.t21 VSSD 0.010639f
C1378 EN.n50 VSSD 0.020752f
C1379 EN.n51 VSSD 0.010998f
C1380 EN.n53 VSSD 0.024943f
C1381 EN.n54 VSSD 0.057288f
C1382 EN.n56 VSSD 0.203308f
C1383 EN.n57 VSSD 0.264704f
C1384 EN.t3 VSSD 0.012222f
C1385 EN.n58 VSSD 0.021676f
C1386 EN.t46 VSSD 0.010639f
C1387 EN.n61 VSSD 0.020752f
C1388 EN.n65 VSSD 0.030424f
C1389 EN.n66 VSSD 0.024316f
C1390 EN.t36 VSSD 0.012222f
C1391 EN.n67 VSSD 0.021676f
C1392 EN.t4 VSSD 0.010639f
C1393 EN.n70 VSSD 0.020752f
C1394 EN.n74 VSSD 0.030424f
C1395 EN.n75 VSSD 0.024316f
C1396 EN.t59 VSSD 0.010639f
C1397 EN.n77 VSSD 0.020752f
C1398 EN.n81 VSSD 0.030424f
C1399 EN.t88 VSSD 0.012222f
C1400 EN.n82 VSSD 0.021676f
C1401 EN.n83 VSSD 0.024316f
C1402 EN.t24 VSSD 0.012222f
C1403 EN.n85 VSSD 0.021676f
C1404 EN.n86 VSSD 0.024316f
C1405 EN.n87 VSSD 0.030424f
C1406 EN.t26 VSSD 0.010639f
C1407 EN.n90 VSSD 0.020752f
C1408 EN.n93 VSSD 0.044103f
C1409 EN.t81 VSSD 0.010639f
C1410 EN.n95 VSSD 0.020752f
C1411 EN.n99 VSSD 0.028368f
C1412 EN.t87 VSSD 0.012222f
C1413 EN.n100 VSSD 0.021676f
C1414 EN.n101 VSSD 0.024316f
C1415 EN.n102 VSSD 0.026204f
C1416 EN.n103 VSSD 0.059519f
C1417 EN.n105 VSSD 0.148087f
C1418 EN.t44 VSSD 0.010639f
C1419 EN.n107 VSSD 0.020752f
C1420 EN.n111 VSSD 0.030424f
C1421 EN.t53 VSSD 0.012222f
C1422 EN.n112 VSSD 0.021676f
C1423 EN.n113 VSSD 0.024316f
C1424 EN.t34 VSSD 0.010639f
C1425 EN.n116 VSSD 0.020752f
C1426 EN.n120 VSSD 0.028368f
C1427 EN.t79 VSSD 0.012222f
C1428 EN.n121 VSSD 0.021676f
C1429 EN.n122 VSSD 0.024316f
C1430 EN.n123 VSSD 0.026204f
C1431 EN.n124 VSSD 0.059519f
C1432 EN.t74 VSSD 0.010514f
C1433 EN.n126 VSSD 0.030213f
C1434 EN.n127 VSSD 0.063748f
C1435 EN.t1 VSSD 0.010639f
C1436 EN.n129 VSSD 0.020752f
C1437 EN.n133 VSSD 0.028368f
C1438 EN.t35 VSSD 0.012222f
C1439 EN.n134 VSSD 0.021676f
C1440 EN.n135 VSSD 0.024316f
C1441 EN.n136 VSSD 0.015321f
C1442 EN.n137 VSSD 0.028424f
C1443 EN.n139 VSSD 0.092067f
C1444 EN.n140 VSSD 0.072397f
C1445 EN.t61 VSSD 0.010639f
C1446 EN.n143 VSSD 0.020752f
C1447 EN.n147 VSSD 0.028368f
C1448 EN.t7 VSSD 0.012222f
C1449 EN.n148 VSSD 0.021676f
C1450 EN.n149 VSSD 0.024316f
C1451 EN.n150 VSSD 0.026204f
C1452 EN.n151 VSSD 0.059519f
C1453 EN.n153 VSSD 0.085077f
C1454 EN.t76 VSSD 0.012222f
C1455 EN.n156 VSSD 0.020964f
C1456 EN.t16 VSSD 0.010639f
C1457 EN.n158 VSSD 0.020752f
C1458 EN.n162 VSSD 0.027903f
C1459 EN.n164 VSSD 0.016978f
C1460 EN.n167 VSSD 0.047218f
C1461 EN.t20 VSSD 0.012222f
C1462 EN.n170 VSSD 0.020964f
C1463 EN.t18 VSSD 0.010639f
C1464 EN.n173 VSSD 0.020752f
C1465 EN.n177 VSSD 0.027903f
C1466 EN.n179 VSSD 0.016978f
C1467 EN.n182 VSSD 0.077441f
C1468 EN.t13 VSSD 0.012222f
C1469 EN.n185 VSSD 0.020964f
C1470 EN.t19 VSSD 0.010639f
C1471 EN.n188 VSSD 0.020752f
C1472 EN.n192 VSSD 0.027903f
C1473 EN.n194 VSSD 0.016978f
C1474 EN.n196 VSSD 0.020211f
C1475 EN.n197 VSSD 0.117453f
C1476 EN.n198 VSSD 0.107044f
C1477 EN.n199 VSSD 0.127062f
C1478 EN.t10 VSSD 0.012222f
C1479 EN.n202 VSSD 0.020964f
C1480 EN.t72 VSSD 0.010639f
C1481 EN.n205 VSSD 0.020752f
C1482 EN.n209 VSSD 0.027903f
C1483 EN.n211 VSSD 0.016978f
C1484 EN.n214 VSSD 0.084492f
C1485 EN.n215 VSSD 0.171048f
C1486 EN.t54 VSSD 0.012222f
C1487 EN.n217 VSSD 0.021702f
C1488 EN.n218 VSSD 0.029635f
C1489 EN.t69 VSSD 0.010639f
C1490 EN.n220 VSSD 0.020752f
C1491 EN.n221 VSSD 0.010998f
C1492 EN.n223 VSSD 0.136876f
C1493 EN.n224 VSSD 0.1318f
C1494 EN.n225 VSSD 0.107047f
C1495 EN.n226 VSSD 0.116327f
C1496 EN.t31 VSSD 0.010639f
C1497 EN.n229 VSSD 0.020752f
C1498 EN.n232 VSSD 0.030424f
C1499 EN.t33 VSSD 0.012222f
C1500 EN.n233 VSSD 0.021676f
C1501 EN.n234 VSSD 0.024316f
C1502 EN.n235 VSSD 0.049501f
C1503 EN.t40 VSSD 0.010639f
C1504 EN.n238 VSSD 0.020752f
C1505 EN.n242 VSSD 0.028368f
C1506 EN.t12 VSSD 0.012222f
C1507 EN.n243 VSSD 0.021676f
C1508 EN.n244 VSSD 0.024316f
C1509 EN.n245 VSSD 0.015321f
C1510 EN.n246 VSSD 0.028424f
C1511 EN.n248 VSSD 0.043099f
C1512 EN.n249 VSSD 0.043662f
C1513 EN.t63 VSSD 0.010639f
C1514 EN.n251 VSSD 0.020752f
C1515 EN.n255 VSSD 0.030424f
C1516 EN.t77 VSSD 0.012222f
C1517 EN.n256 VSSD 0.021676f
C1518 EN.n257 VSSD 0.024316f
C1519 EN.n258 VSSD 0.06473f
C1520 EN.n259 VSSD 0.019811f
C1521 EN.n260 VSSD 0.057288f
C1522 CF[0].t8 VSSD 0.011843f
C1523 CF[0].n0 VSSD 0.021695f
C1524 CF[0].n1 VSSD 0.010209f
C1525 CF[0].t10 VSSD 0.011843f
C1526 CF[0].n2 VSSD 0.021641f
C1527 CF[0].n4 VSSD 0.067494f
C1528 CF[0].t9 VSSD 0.012146f
C1529 CF[0].t6 VSSD 0.011592f
C1530 CF[0].n5 VSSD 0.014324f
C1531 CF[0].t7 VSSD 0.011592f
C1532 CF[0].n6 VSSD 0.016294f
C1533 CF[0].n11 VSSD 0.021989f
C1534 CF[0].n12 VSSD 0.013315f
C1535 CF[0].n13 VSSD 0.244631f
C1536 CF[0].n14 VSSD 0.27455f
C1537 CF[0].n15 VSSD 0.014606f
C1538 CF[0].n18 VSSD 0.011656f
C1539 CF[0].n20 VSSD 0.34767f
C1540 CLKS.t104 VSSD 0.011237f
C1541 CLKS.n4 VSSD 0.02192f
C1542 CLKS.n5 VSSD 0.011617f
C1543 CLKS.n7 VSSD 0.022515f
C1544 CLKS.t94 VSSD 0.01291f
C1545 CLKS.n8 VSSD 0.022924f
C1546 CLKS.n9 VSSD 0.029465f
C1547 CLKS.t60 VSSD 0.01291f
C1548 CLKS.n10 VSSD 0.022924f
C1549 CLKS.n11 VSSD 0.029465f
C1550 CLKS.t103 VSSD 0.011237f
C1551 CLKS.n14 VSSD 0.02192f
C1552 CLKS.n15 VSSD 0.011617f
C1553 CLKS.n17 VSSD 0.011019f
C1554 CLKS.n18 VSSD 0.016719f
C1555 CLKS.n19 VSSD 0.025972f
C1556 CLKS.t123 VSSD 0.01291f
C1557 CLKS.n20 VSSD 0.022924f
C1558 CLKS.n21 VSSD 0.029465f
C1559 CLKS.t135 VSSD 0.011237f
C1560 CLKS.n26 VSSD 0.02192f
C1561 CLKS.n27 VSSD 0.011617f
C1562 CLKS.n29 VSSD 0.026347f
C1563 CLKS.n30 VSSD 0.060512f
C1564 CLKS.n32 VSSD 0.083079f
C1565 CLKS.t66 VSSD 0.01291f
C1566 CLKS.n34 VSSD 0.022924f
C1567 CLKS.n35 VSSD 0.031303f
C1568 CLKS.t137 VSSD 0.011237f
C1569 CLKS.n39 VSSD 0.02192f
C1570 CLKS.n40 VSSD 0.011617f
C1571 CLKS.t50 VSSD 0.01291f
C1572 CLKS.n42 VSSD 0.022896f
C1573 CLKS.t49 VSSD 0.011237f
C1574 CLKS.n45 VSSD 0.02192f
C1575 CLKS.n46 VSSD 0.011617f
C1576 CLKS.n48 VSSD 0.031303f
C1577 CLKS.n49 VSSD 0.052538f
C1578 CLKS.n50 VSSD 0.063722f
C1579 CLKS.t34 VSSD 0.01291f
C1580 CLKS.n51 VSSD 0.022924f
C1581 CLKS.n52 VSSD 0.029518f
C1582 CLKS.t106 VSSD 0.011237f
C1583 CLKS.n57 VSSD 0.02192f
C1584 CLKS.n58 VSSD 0.011617f
C1585 CLKS.n60 VSSD 0.029335f
C1586 CLKS.n61 VSSD 0.017856f
C1587 CLKS.n62 VSSD 0.048441f
C1588 CLKS.n63 VSSD 0.017856f
C1589 CLKS.n64 VSSD 0.017856f
C1590 CLKS.n65 VSSD 0.011891f
C1591 CLKS.n66 VSSD 0.011891f
C1592 CLKS.n67 VSSD 0.011891f
C1593 CLKS.n68 VSSD 0.011891f
C1594 CLKS.n69 VSSD 0.040647f
C1595 CLKS.n70 VSSD 0.035608f
C1596 CLKS.n71 VSSD 0.035608f
C1597 CLKS.n72 VSSD 0.040902f
C1598 CLKS.n73 VSSD 0.048598f
C1599 CLKS.n74 VSSD 0.046618f
C1600 CLKS.n75 VSSD 0.023673f
C1601 CLKS.n76 VSSD 0.016129f
C1602 CLKS.n77 VSSD 0.02214f
C1603 CLKS.t74 VSSD 0.01291f
C1604 CLKS.n78 VSSD 0.022904f
C1605 CLKS.n79 VSSD 0.037839f
C1606 CLKS.t19 VSSD 0.011237f
C1607 CLKS.n84 VSSD 0.02192f
C1608 CLKS.n85 VSSD 0.011617f
C1609 CLKS.n87 VSSD 0.030179f
C1610 CLKS.n88 VSSD 0.071073f
C1611 CLKS.n90 VSSD 0.07805f
C1612 CLKS.n91 VSSD 0.017052f
C1613 CLKS.t82 VSSD 0.011237f
C1614 CLKS.n94 VSSD 0.02192f
C1615 CLKS.n95 VSSD 0.011617f
C1616 CLKS.n97 VSSD 0.031303f
C1617 CLKS.t130 VSSD 0.01291f
C1618 CLKS.n98 VSSD 0.022143f
C1619 CLKS.n99 VSSD 0.017933f
C1620 CLKS.n103 VSSD 0.049885f
C1621 CLKS.t119 VSSD 0.01291f
C1622 CLKS.n104 VSSD 0.022924f
C1623 CLKS.n105 VSSD 0.029465f
C1624 CLKS.t117 VSSD 0.011237f
C1625 CLKS.n110 VSSD 0.02192f
C1626 CLKS.n111 VSSD 0.011617f
C1627 CLKS.n113 VSSD 0.022515f
C1628 CLKS.n114 VSSD 0.049564f
C1629 CLKS.n116 VSSD 0.099857f
C1630 CLKS.n117 VSSD 0.10344f
C1631 CLKS.t56 VSSD 0.01291f
C1632 CLKS.n118 VSSD 0.022904f
C1633 CLKS.n119 VSSD 0.037839f
C1634 CLKS.t89 VSSD 0.011237f
C1635 CLKS.n122 VSSD 0.02192f
C1636 CLKS.n123 VSSD 0.011617f
C1637 CLKS.n125 VSSD 0.030179f
C1638 CLKS.n126 VSSD 0.071073f
C1639 CLKS.n128 VSSD 0.132608f
C1640 CLKS.n129 VSSD 0.017052f
C1641 CLKS.t101 VSSD 0.011237f
C1642 CLKS.n132 VSSD 0.02192f
C1643 CLKS.n133 VSSD 0.011617f
C1644 CLKS.n135 VSSD 0.031303f
C1645 CLKS.t70 VSSD 0.01291f
C1646 CLKS.n136 VSSD 0.022143f
C1647 CLKS.n137 VSSD 0.017933f
C1648 CLKS.t21 VSSD 0.011237f
C1649 CLKS.n145 VSSD 0.02192f
C1650 CLKS.n146 VSSD 0.011617f
C1651 CLKS.t23 VSSD 0.01291f
C1652 CLKS.n148 VSSD 0.022924f
C1653 CLKS.n149 VSSD 0.031759f
C1654 CLKS.n151 VSSD 0.070333f
C1655 CLKS.t24 VSSD 0.01291f
C1656 CLKS.n153 VSSD 0.022896f
C1657 CLKS.n154 VSSD 0.025684f
C1658 CLKS.n155 VSSD 0.032136f
C1659 CLKS.t81 VSSD 0.011237f
C1660 CLKS.n158 VSSD 0.02192f
C1661 CLKS.n160 VSSD 0.012926f
C1662 CLKS.t51 VSSD 0.013306f
C1663 CLKS.n161 VSSD 0.025061f
C1664 CLKS.n162 VSSD 0.02441f
C1665 CLKS.n163 VSSD 0.167703f
C1666 CLKS.t120 VSSD 0.011237f
C1667 CLKS.n166 VSSD 0.02192f
C1668 CLKS.n170 VSSD 0.029964f
C1669 CLKS.t93 VSSD 0.01291f
C1670 CLKS.n171 VSSD 0.022896f
C1671 CLKS.n172 VSSD 0.025684f
C1672 CLKS.n173 VSSD 0.016184f
C1673 CLKS.n174 VSSD 0.030024f
C1674 CLKS.t52 VSSD 0.01291f
C1675 CLKS.n177 VSSD 0.022896f
C1676 CLKS.n178 VSSD 0.025684f
C1677 CLKS.n179 VSSD 0.032136f
C1678 CLKS.t20 VSSD 0.011237f
C1679 CLKS.n182 VSSD 0.02192f
C1680 CLKS.n184 VSSD 0.042721f
C1681 CLKS.t30 VSSD 0.01291f
C1682 CLKS.n185 VSSD 0.022896f
C1683 CLKS.t58 VSSD 0.011237f
C1684 CLKS.n190 VSSD 0.02192f
C1685 CLKS.n191 VSSD 0.011617f
C1686 CLKS.n193 VSSD 0.031303f
C1687 CLKS.n194 VSSD 0.08484f
C1688 CLKS.n195 VSSD 0.086251f
C1689 CLKS.n196 VSSD 0.021268f
C1690 CLKS.n198 VSSD 0.028107f
C1691 CLKS.t76 VSSD 0.01291f
C1692 CLKS.n199 VSSD 0.022896f
C1693 CLKS.t111 VSSD 0.011237f
C1694 CLKS.n204 VSSD 0.02192f
C1695 CLKS.n205 VSSD 0.011617f
C1696 CLKS.n207 VSSD 0.031303f
C1697 CLKS.n208 VSSD 0.13862f
C1698 CLKS.n209 VSSD 0.02128f
C1699 CLKS.n211 VSSD 0.171247f
C1700 CLKS.n212 VSSD 0.156678f
C1701 CLKS.n213 VSSD 0.076752f
C1702 CLKS.n214 VSSD 0.08105f
C1703 CLKS.t18 VSSD 0.011237f
C1704 CLKS.n216 VSSD 0.02192f
C1705 CLKS.n220 VSSD 0.029964f
C1706 CLKS.t91 VSSD 0.01291f
C1707 CLKS.n221 VSSD 0.022896f
C1708 CLKS.n222 VSSD 0.025684f
C1709 CLKS.n223 VSSD 0.027679f
C1710 CLKS.n224 VSSD 0.062868f
C1711 CLKS.n226 VSSD 0.059624f
C1712 CLKS.t112 VSSD 0.01291f
C1713 CLKS.n227 VSSD 0.022896f
C1714 CLKS.n228 VSSD 0.025684f
C1715 CLKS.n229 VSSD 0.032136f
C1716 CLKS.t115 VSSD 0.011237f
C1717 CLKS.n232 VSSD 0.02192f
C1718 CLKS.n236 VSSD 0.044965f
C1719 CLKS.t31 VSSD 0.01291f
C1720 CLKS.n238 VSSD 0.022896f
C1721 CLKS.n239 VSSD 0.025684f
C1722 CLKS.n240 VSSD 0.032136f
C1723 CLKS.t32 VSSD 0.011237f
C1724 CLKS.n243 VSSD 0.02192f
C1725 CLKS.n246 VSSD 0.134786f
C1726 CLKS.n247 VSSD 0.103623f
C1727 CLKS.t36 VSSD 0.011237f
C1728 CLKS.n249 VSSD 0.02192f
C1729 CLKS.n253 VSSD 0.029964f
C1730 CLKS.t107 VSSD 0.01291f
C1731 CLKS.n254 VSSD 0.022896f
C1732 CLKS.n255 VSSD 0.025684f
C1733 CLKS.n256 VSSD 0.027679f
C1734 CLKS.n257 VSSD 0.062868f
C1735 CLKS.n259 VSSD 0.058382f
C1736 CLKS.t33 VSSD 0.011237f
C1737 CLKS.n261 VSSD 0.02192f
C1738 CLKS.n265 VSSD 0.029964f
C1739 CLKS.t105 VSSD 0.01291f
C1740 CLKS.n266 VSSD 0.022896f
C1741 CLKS.n267 VSSD 0.025684f
C1742 CLKS.n268 VSSD 0.027679f
C1743 CLKS.n269 VSSD 0.062868f
C1744 CLKS.n271 VSSD 0.017052f
C1745 CLKS.t98 VSSD 0.011237f
C1746 CLKS.n274 VSSD 0.02192f
C1747 CLKS.n275 VSSD 0.011617f
C1748 CLKS.n277 VSSD 0.031303f
C1749 CLKS.t55 VSSD 0.01291f
C1750 CLKS.n278 VSSD 0.022143f
C1751 CLKS.n279 VSSD 0.017933f
C1752 CLKS.n282 VSSD 0.033904f
C1753 CLKS.t85 VSSD 0.01291f
C1754 CLKS.n284 VSSD 0.022896f
C1755 CLKS.n285 VSSD 0.025684f
C1756 CLKS.n286 VSSD 0.032136f
C1757 CLKS.t86 VSSD 0.011237f
C1758 CLKS.n289 VSSD 0.02192f
C1759 CLKS.n293 VSSD 0.20624f
C1760 CLKS.n294 VSSD 0.108778f
C1761 CLKS.t48 VSSD 0.011237f
C1762 CLKS.n297 VSSD 0.02192f
C1763 CLKS.n301 VSSD 0.029964f
C1764 CLKS.t46 VSSD 0.01291f
C1765 CLKS.n302 VSSD 0.022896f
C1766 CLKS.n303 VSSD 0.025684f
C1767 CLKS.n304 VSSD 0.027679f
C1768 CLKS.n305 VSSD 0.062868f
C1769 CLKS.n307 VSSD 0.042678f
C1770 CLKS.t140 VSSD 0.01291f
C1771 CLKS.n308 VSSD 0.022896f
C1772 CLKS.n309 VSSD 0.025684f
C1773 CLKS.n310 VSSD 0.032136f
C1774 CLKS.t68 VSSD 0.011237f
C1775 CLKS.n312 VSSD 0.02192f
C1776 CLKS.n316 VSSD 0.036971f
C1777 CLKS.n317 VSSD 0.113798f
C1778 CLKS.n318 VSSD 0.135758f
C1779 CLKS.t109 VSSD 0.01291f
C1780 CLKS.n320 VSSD 0.022896f
C1781 CLKS.n321 VSSD 0.025684f
C1782 CLKS.n322 VSSD 0.032136f
C1783 CLKS.t78 VSSD 0.011237f
C1784 CLKS.n325 VSSD 0.02192f
C1785 CLKS.n328 VSSD 0.037548f
C1786 CLKS.n329 VSSD 0.15959f
C1787 CLKS.n330 VSSD 0.122142f
C1788 CLKS.t16 VSSD 0.011237f
C1789 CLKS.n331 VSSD 0.02192f
C1790 CLKS.t90 VSSD 0.01291f
C1791 CLKS.n335 VSSD 0.022896f
C1792 CLKS.n336 VSSD 0.025684f
C1793 CLKS.n337 VSSD 0.032136f
C1794 CLKS.n338 VSSD 0.028408f
C1795 CLKS.n339 VSSD 0.050019f
C1796 CLKS.n340 VSSD 0.107547f
C1797 CLKS.n341 VSSD 0.051776f
C1798 CLKS.t38 VSSD 0.011237f
C1799 CLKS.n347 VSSD 0.02192f
C1800 CLKS.n348 VSSD 0.011617f
C1801 CLKS.n350 VSSD 0.031303f
C1802 CLKS.t87 VSSD 0.01291f
C1803 CLKS.n351 VSSD 0.022143f
C1804 CLKS.n352 VSSD 0.017933f
C1805 CLKS.n355 VSSD 0.011091f
C1806 CLKS.n356 VSSD 0.13476f
C1807 CLKS.n357 VSSD 0.14485f
C1808 CLKS.t127 VSSD 0.011237f
C1809 CLKS.n361 VSSD 0.02192f
C1810 CLKS.n362 VSSD 0.011617f
C1811 CLKS.n364 VSSD 0.031303f
C1812 CLKS.t57 VSSD 0.01291f
C1813 CLKS.n365 VSSD 0.022143f
C1814 CLKS.n366 VSSD 0.017933f
C1815 CLKS.n370 VSSD 0.040125f
C1816 CLKS.n371 VSSD 0.011084f
C1817 CLKS.n372 VSSD 0.049564f
C1818 clknet_1_1__leaf_CLK.t4 VSSD 0.015383f
C1819 clknet_1_1__leaf_CLK.t11 VSSD 0.015383f
C1820 clknet_1_1__leaf_CLK.n0 VSSD 0.039077f
C1821 clknet_1_1__leaf_CLK.t0 VSSD 0.015383f
C1822 clknet_1_1__leaf_CLK.t2 VSSD 0.015383f
C1823 clknet_1_1__leaf_CLK.n1 VSSD 0.032425f
C1824 clknet_1_1__leaf_CLK.n2 VSSD 0.147771f
C1825 clknet_1_1__leaf_CLK.t10 VSSD 0.015383f
C1826 clknet_1_1__leaf_CLK.t14 VSSD 0.015383f
C1827 clknet_1_1__leaf_CLK.n3 VSSD 0.032425f
C1828 clknet_1_1__leaf_CLK.n4 VSSD 0.085123f
C1829 clknet_1_1__leaf_CLK.t9 VSSD 0.015383f
C1830 clknet_1_1__leaf_CLK.t13 VSSD 0.015383f
C1831 clknet_1_1__leaf_CLK.n5 VSSD 0.032425f
C1832 clknet_1_1__leaf_CLK.n6 VSSD 0.084727f
C1833 clknet_1_1__leaf_CLK.t8 VSSD 0.015383f
C1834 clknet_1_1__leaf_CLK.t3 VSSD 0.015383f
C1835 clknet_1_1__leaf_CLK.n7 VSSD 0.032425f
C1836 clknet_1_1__leaf_CLK.n8 VSSD 0.084727f
C1837 clknet_1_1__leaf_CLK.t37 VSSD 0.01611f
C1838 clknet_1_1__leaf_CLK.t35 VSSD 0.024079f
C1839 clknet_1_1__leaf_CLK.n9 VSSD 0.044503f
C1840 clknet_1_1__leaf_CLK.n10 VSSD 0.013075f
C1841 clknet_1_1__leaf_CLK.t47 VSSD 0.01611f
C1842 clknet_1_1__leaf_CLK.t40 VSSD 0.024079f
C1843 clknet_1_1__leaf_CLK.n11 VSSD 0.044503f
C1844 clknet_1_1__leaf_CLK.n12 VSSD 0.01642f
C1845 clknet_1_1__leaf_CLK.n13 VSSD 0.08278f
C1846 clknet_1_1__leaf_CLK.t33 VSSD 0.024079f
C1847 clknet_1_1__leaf_CLK.t32 VSSD 0.01611f
C1848 clknet_1_1__leaf_CLK.n14 VSSD 0.044f
C1849 clknet_1_1__leaf_CLK.n15 VSSD 0.013075f
C1850 clknet_1_1__leaf_CLK.t44 VSSD 0.01611f
C1851 clknet_1_1__leaf_CLK.t38 VSSD 0.024079f
C1852 clknet_1_1__leaf_CLK.n16 VSSD 0.044111f
C1853 clknet_1_1__leaf_CLK.n17 VSSD 0.079682f
C1854 clknet_1_1__leaf_CLK.n18 VSSD 0.322945f
C1855 clknet_1_1__leaf_CLK.t45 VSSD 0.024079f
C1856 clknet_1_1__leaf_CLK.t43 VSSD 0.01611f
C1857 clknet_1_1__leaf_CLK.n19 VSSD 0.044f
C1858 clknet_1_1__leaf_CLK.n20 VSSD 0.013075f
C1859 clknet_1_1__leaf_CLK.n21 VSSD 0.135286f
C1860 clknet_1_1__leaf_CLK.t48 VSSD 0.024079f
C1861 clknet_1_1__leaf_CLK.t46 VSSD 0.01611f
C1862 clknet_1_1__leaf_CLK.n22 VSSD 0.044f
C1863 clknet_1_1__leaf_CLK.n23 VSSD 0.013075f
C1864 clknet_1_1__leaf_CLK.t39 VSSD 0.024079f
C1865 clknet_1_1__leaf_CLK.t42 VSSD 0.01611f
C1866 clknet_1_1__leaf_CLK.n24 VSSD 0.044f
C1867 clknet_1_1__leaf_CLK.n26 VSSD 0.040292f
C1868 clknet_1_1__leaf_CLK.t41 VSSD 0.01611f
C1869 clknet_1_1__leaf_CLK.t36 VSSD 0.024079f
C1870 clknet_1_1__leaf_CLK.n27 VSSD 0.044111f
C1871 clknet_1_1__leaf_CLK.n28 VSSD 0.020133f
C1872 clknet_1_1__leaf_CLK.n29 VSSD 0.224038f
C1873 clknet_1_1__leaf_CLK.t34 VSSD 0.024079f
C1874 clknet_1_1__leaf_CLK.t49 VSSD 0.01611f
C1875 clknet_1_1__leaf_CLK.n30 VSSD 0.044f
C1876 clknet_1_1__leaf_CLK.n31 VSSD 0.013075f
C1877 clknet_1_1__leaf_CLK.t55 VSSD 0.01611f
C1878 clknet_1_1__leaf_CLK.t51 VSSD 0.024079f
C1879 clknet_1_1__leaf_CLK.n32 VSSD 0.044503f
C1880 clknet_1_1__leaf_CLK.n33 VSSD 0.117161f
C1881 clknet_1_1__leaf_CLK.n34 VSSD 0.30967f
C1882 clknet_1_1__leaf_CLK.n35 VSSD 0.118273f
C1883 clknet_1_1__leaf_CLK.n36 VSSD 0.349868f
C1884 clknet_1_1__leaf_CLK.t53 VSSD 0.024079f
C1885 clknet_1_1__leaf_CLK.t52 VSSD 0.01611f
C1886 clknet_1_1__leaf_CLK.n37 VSSD 0.044f
C1887 clknet_1_1__leaf_CLK.n38 VSSD 0.013075f
C1888 clknet_1_1__leaf_CLK.n39 VSSD 0.234317f
C1889 clknet_1_1__leaf_CLK.n40 VSSD 0.15751f
C1890 clknet_1_1__leaf_CLK.n41 VSSD 0.131831f
C1891 clknet_1_1__leaf_CLK.t54 VSSD 0.01611f
C1892 clknet_1_1__leaf_CLK.t50 VSSD 0.024079f
C1893 clknet_1_1__leaf_CLK.n42 VSSD 0.044111f
C1894 clknet_1_1__leaf_CLK.n43 VSSD 0.062931f
C1895 clknet_1_1__leaf_CLK.n44 VSSD 0.246453f
C1896 clknet_1_1__leaf_CLK.t5 VSSD 0.015383f
C1897 clknet_1_1__leaf_CLK.t12 VSSD 0.015383f
C1898 clknet_1_1__leaf_CLK.n45 VSSD 0.030766f
C1899 clknet_1_1__leaf_CLK.n46 VSSD 0.032542f
C1900 clknet_1_1__leaf_CLK.n47 VSSD 0.05129f
C1901 clknet_1_1__leaf_CLK.t1 VSSD 0.015383f
C1902 clknet_1_1__leaf_CLK.t7 VSSD 0.015383f
C1903 clknet_1_1__leaf_CLK.n48 VSSD 0.032425f
C1904 clknet_1_1__leaf_CLK.n49 VSSD 0.073111f
C1905 clknet_1_1__leaf_CLK.t15 VSSD 0.015383f
C1906 clknet_1_1__leaf_CLK.t6 VSSD 0.015383f
C1907 clknet_1_1__leaf_CLK.n50 VSSD 0.032004f
C1908 clknet_1_1__leaf_CLK.n51 VSSD 0.100676f
C1909 clknet_1_1__leaf_CLK.n52 VSSD 0.022942f
C1910 clknet_1_1__leaf_CLK.n53 VSSD 0.014749f
C1911 clknet_1_1__leaf_CLK.n54 VSSD 0.093196f
C1912 clknet_1_1__leaf_CLK.n55 VSSD 0.014749f
C1913 clknet_1_1__leaf_CLK.n56 VSSD 0.056018f
C1914 clknet_1_1__leaf_CLK.n57 VSSD 0.014758f
C1915 clknet_1_1__leaf_CLK.n58 VSSD 0.057784f
C1916 clknet_1_1__leaf_CLK.n59 VSSD 0.014749f
C1917 clknet_1_1__leaf_CLK.n60 VSSD 0.056018f
C1918 clknet_1_1__leaf_CLK.n61 VSSD 0.014749f
C1919 clknet_1_1__leaf_CLK.n62 VSSD 0.056298f
C1920 clknet_1_1__leaf_CLK.n63 VSSD 0.014749f
C1921 clknet_1_1__leaf_CLK.n64 VSSD 0.048359f
C1922 clknet_1_1__leaf_CLK.n65 VSSD 0.014238f
C1923 clknet_1_1__leaf_CLK.n66 VSSD 0.046786f
C1924 VDDD.t2047 VSSD 0.011775f
C1925 VDDD.t1998 VSSD 0.081647f
C1926 VDDD.n5 VSSD 0.038136f
C1927 VDDD.t2059 VSSD 0.081647f
C1928 VDDD.n12 VSSD 0.038136f
C1929 VDDD.n15 VSSD 0.014016f
C1930 VDDD.n26 VSSD 0.138631f
C1931 VDDD.n34 VSSD 0.013708f
C1932 VDDD.t2036 VSSD 0.023382f
C1933 VDDD.n41 VSSD 0.138631f
C1934 VDDD.t2048 VSSD 0.011775f
C1935 VDDD.n51 VSSD 0.017816f
C1936 VDDD.t2092 VSSD 0.081647f
C1937 VDDD.t2029 VSSD 0.081647f
C1938 VDDD.n74 VSSD 0.038136f
C1939 VDDD.n107 VSSD 0.038136f
C1940 VDDD.n113 VSSD 0.149079f
C1941 VDDD.t2007 VSSD 0.081647f
C1942 VDDD.n123 VSSD 0.038136f
C1943 VDDD.t2072 VSSD 0.011775f
C1944 VDDD.t1853 VSSD 0.032961f
C1945 VDDD.t1027 VSSD 0.132808f
C1946 VDDD.t981 VSSD 0.132808f
C1947 VDDD.t508 VSSD 0.035247f
C1948 VDDD.n129 VSSD 0.035054f
C1949 VDDD.n131 VSSD 0.015264f
C1950 VDDD.t2099 VSSD 0.011775f
C1951 VDDD.n133 VSSD 0.017816f
C1952 VDDD.n134 VSSD 0.014638f
C1953 VDDD.n139 VSSD 0.013974f
C1954 VDDD.n142 VSSD 0.017816f
C1955 VDDD.n143 VSSD 0.014638f
C1956 VDDD.t2027 VSSD 0.081647f
C1957 VDDD.n174 VSSD 0.038136f
C1958 VDDD.n205 VSSD 0.140415f
C1959 VDDD.n207 VSSD 0.244388f
C1960 VDDD.t2013 VSSD 0.081647f
C1961 VDDD.t2060 VSSD 0.081647f
C1962 VDDD.n225 VSSD 0.038136f
C1963 VDDD.t1003 VSSD 0.058119f
C1964 VDDD.n233 VSSD 0.026834f
C1965 VDDD.n234 VSSD 0.018019f
C1966 VDDD.t2002 VSSD 0.042267f
C1967 VDDD.n236 VSSD 0.076191f
C1968 VDDD.n237 VSSD 0.022234f
C1969 VDDD.n246 VSSD 0.011268f
C1970 VDDD.n248 VSSD 0.016244f
C1971 VDDD.n249 VSSD 0.01711f
C1972 VDDD.n253 VSSD 0.024266f
C1973 VDDD.n254 VSSD 0.018019f
C1974 VDDD.n255 VSSD 0.029567f
C1975 VDDD.t1984 VSSD 0.040373f
C1976 VDDD.n256 VSSD 0.049034f
C1977 VDDD.n257 VSSD 0.018973f
C1978 VDDD.n258 VSSD 0.011892f
C1979 VDDD.t1987 VSSD 0.011988f
C1980 VDDD.n260 VSSD 0.030737f
C1981 VDDD.n261 VSSD 0.016743f
C1982 VDDD.t2052 VSSD 0.011988f
C1983 VDDD.n264 VSSD 0.030737f
C1984 VDDD.n265 VSSD 0.016743f
C1985 VDDD.n266 VSSD 0.013794f
C1986 VDDD.n267 VSSD 0.022897f
C1987 VDDD.n268 VSSD 0.042531f
C1988 VDDD.t1856 VSSD 0.084633f
C1989 VDDD.t1079 VSSD 0.071906f
C1990 VDDD.t565 VSSD 0.045604f
C1991 VDDD.t563 VSSD 0.030757f
C1992 VDDD.t1365 VSSD 0.050483f
C1993 VDDD.t1866 VSSD 0.040726f
C1994 VDDD.t561 VSSD 0.040726f
C1995 VDDD.t1368 VSSD 0.036059f
C1996 VDDD.t1509 VSSD 0.032029f
C1997 VDDD.t1758 VSSD 0.020999f
C1998 VDDD.t1903 VSSD 0.048998f
C1999 VDDD.t1591 VSSD 0.062361f
C2000 VDDD.t678 VSSD 0.050271f
C2001 VDDD.t1508 VSSD 0.041362f
C2002 VDDD.t83 VSSD 0.028848f
C2003 VDDD.t1195 VSSD 0.076149f
C2004 VDDD.t1454 VSSD 0.074452f
C2005 VDDD.t135 VSSD 0.031605f
C2006 VDDD.t1138 VSSD 0.015909f
C2007 VDDD.n269 VSSD 0.013532f
C2008 VDDD.n270 VSSD 0.010882f
C2009 VDDD.n282 VSSD 0.019037f
C2010 VDDD.t2097 VSSD 0.011988f
C2011 VDDD.n284 VSSD 0.030737f
C2012 VDDD.n285 VSSD 0.016743f
C2013 VDDD.t2028 VSSD 0.042035f
C2014 VDDD.n286 VSSD 0.070387f
C2015 VDDD.n287 VSSD 0.014424f
C2016 VDDD.n288 VSSD 0.026923f
C2017 VDDD.n289 VSSD 0.039466f
C2018 VDDD.t2094 VSSD 0.023588f
C2019 VDDD.n291 VSSD 0.04098f
C2020 VDDD.n292 VSSD 0.023515f
C2021 VDDD.t2074 VSSD 0.011988f
C2022 VDDD.n294 VSSD 0.030737f
C2023 VDDD.n295 VSSD 0.016743f
C2024 VDDD.t2001 VSSD 0.011988f
C2025 VDDD.n297 VSSD 0.030737f
C2026 VDDD.n298 VSSD 0.016743f
C2027 VDDD.n300 VSSD 0.013785f
C2028 VDDD.n301 VSSD 0.02207f
C2029 VDDD.n305 VSSD 0.015017f
C2030 VDDD.n313 VSSD 0.012503f
C2031 VDDD.n329 VSSD 0.011873f
C2032 VDDD.n336 VSSD 0.014873f
C2033 VDDD.n341 VSSD 0.244388f
C2034 VDDD.t2091 VSSD 0.081647f
C2035 VDDD.n362 VSSD 0.138631f
C2036 VDDD.t1986 VSSD 0.023382f
C2037 VDDD.n376 VSSD 0.013148f
C2038 VDDD.t2062 VSSD 0.081647f
C2039 VDDD.t2018 VSSD 0.023382f
C2040 VDDD.t490 VSSD 0.058119f
C2041 VDDD.t1328 VSSD 0.032878f
C2042 VDDD.t50 VSSD 0.020999f
C2043 VDDD.t139 VSSD 0.032029f
C2044 VDDD.t177 VSSD 0.031817f
C2045 VDDD.t900 VSSD 0.01909f
C2046 VDDD.t217 VSSD 0.013787f
C2047 VDDD.t784 VSSD 0.017817f
C2048 VDDD.t1911 VSSD 0.017817f
C2049 VDDD.t1924 VSSD 0.045604f
C2050 VDDD.t835 VSSD 0.056634f
C2051 VDDD.t1243 VSSD 0.017817f
C2052 VDDD.t837 VSSD 0.019514f
C2053 VDDD.t693 VSSD 0.027787f
C2054 VDDD.t1262 VSSD 0.041362f
C2055 VDDD.t94 VSSD 0.050271f
C2056 VDDD.t1868 VSSD 0.062361f
C2057 VDDD.t1935 VSSD 0.048998f
C2058 VDDD.t1141 VSSD 0.020999f
C2059 VDDD.t1261 VSSD 0.032029f
C2060 VDDD.t200 VSSD 0.036059f
C2061 VDDD.t13 VSSD 0.040726f
C2062 VDDD.t1864 VSSD 0.040726f
C2063 VDDD.t119 VSSD 0.050483f
C2064 VDDD.t1654 VSSD 0.030757f
C2065 VDDD.t1652 VSSD 0.019939f
C2066 VDDD.t1764 VSSD 0.027787f
C2067 VDDD.t499 VSSD 0.042976f
C2068 VDDD.n394 VSSD 0.012834f
C2069 VDDD.t2078 VSSD 0.012029f
C2070 VDDD.n395 VSSD 0.021885f
C2071 VDDD.n397 VSSD 0.021823f
C2072 VDDD.t2084 VSSD 0.011988f
C2073 VDDD.n399 VSSD 0.030737f
C2074 VDDD.n400 VSSD 0.016743f
C2075 VDDD.t2064 VSSD 0.011988f
C2076 VDDD.n402 VSSD 0.030737f
C2077 VDDD.n403 VSSD 0.016743f
C2078 VDDD.n404 VSSD 0.013794f
C2079 VDDD.n411 VSSD 0.021149f
C2080 VDDD.n413 VSSD 0.01711f
C2081 VDDD.n414 VSSD 0.011268f
C2082 VDDD.n416 VSSD 0.016244f
C2083 VDDD.n428 VSSD 0.038136f
C2084 VDDD.n455 VSSD 0.011099f
C2085 VDDD.n471 VSSD 0.021149f
C2086 VDDD.n472 VSSD 0.013033f
C2087 VDDD.n474 VSSD 0.013752f
C2088 VDDD.n475 VSSD 0.011522f
C2089 VDDD.n479 VSSD 0.017987f
C2090 VDDD.t2010 VSSD 0.011988f
C2091 VDDD.n481 VSSD 0.030737f
C2092 VDDD.n482 VSSD 0.016743f
C2093 VDDD.n496 VSSD 0.014424f
C2094 VDDD.t1988 VSSD 0.042035f
C2095 VDDD.n497 VSSD 0.070387f
C2096 VDDD.n498 VSSD 0.018492f
C2097 VDDD.n500 VSSD 0.011438f
C2098 VDDD.n503 VSSD 0.017135f
C2099 VDDD.t2034 VSSD 0.012068f
C2100 VDDD.n504 VSSD 0.019643f
C2101 VDDD.n506 VSSD 0.015041f
C2102 VDDD.n509 VSSD 0.016365f
C2103 VDDD.t2005 VSSD 0.042191f
C2104 VDDD.n510 VSSD 0.052548f
C2105 VDDD.n511 VSSD 0.023078f
C2106 VDDD.n513 VSSD 0.013464f
C2107 VDDD.n515 VSSD 0.01367f
C2108 VDDD.n518 VSSD 0.014295f
C2109 VDDD.t2016 VSSD 0.023382f
C2110 VDDD.n522 VSSD 0.021181f
C2111 VDDD.n524 VSSD 0.015644f
C2112 VDDD.n525 VSSD 0.013913f
C2113 VDDD.n539 VSSD 0.011567f
C2114 VDDD.n540 VSSD 0.014239f
C2115 VDDD.n541 VSSD 0.011472f
C2116 VDDD.n542 VSSD 0.010239f
C2117 VDDD.n545 VSSD 0.011021f
C2118 VDDD.n548 VSSD 0.01557f
C2119 VDDD.n552 VSSD 0.013033f
C2120 VDDD.n553 VSSD 0.017188f
C2121 VDDD.n554 VSSD 0.013558f
C2122 VDDD.n561 VSSD 0.171505f
C2123 VDDD.n562 VSSD 0.33981f
C2124 VDDD.n564 VSSD 0.221962f
C2125 VDDD.t2057 VSSD 0.041456f
C2126 VDDD.n574 VSSD 0.019389f
C2127 VDDD.n577 VSSD 0.02077f
C2128 VDDD.t2103 VSSD 0.042046f
C2129 VDDD.n578 VSSD 0.063281f
C2130 VDDD.n579 VSSD 0.013486f
C2131 VDDD.n581 VSSD 0.01681f
C2132 VDDD.n595 VSSD 0.010305f
C2133 VDDD.n616 VSSD 0.013558f
C2134 VDDD.n617 VSSD 0.019992f
C2135 VDDD.n620 VSSD 0.021637f
C2136 VDDD.n621 VSSD 0.039466f
C2137 VDDD.n622 VSSD 0.030897f
C2138 VDDD.n626 VSSD 0.221962f
C2139 VDDD.t2014 VSSD 0.011988f
C2140 VDDD.n634 VSSD 0.030737f
C2141 VDDD.n635 VSSD 0.015201f
C2142 VDDD.n636 VSSD 0.01426f
C2143 VDDD.n637 VSSD 0.018492f
C2144 VDDD.t2113 VSSD 0.042035f
C2145 VDDD.n638 VSSD 0.070387f
C2146 VDDD.n639 VSSD 0.014424f
C2147 VDDD.n640 VSSD 0.021661f
C2148 VDDD.n642 VSSD 0.013386f
C2149 VDDD.n647 VSSD 0.010704f
C2150 VDDD.t1790 VSSD 0.058119f
C2151 VDDD.t2104 VSSD 0.011988f
C2152 VDDD.n671 VSSD 0.030737f
C2153 VDDD.n672 VSSD 0.016743f
C2154 VDDD.t2067 VSSD 0.011988f
C2155 VDDD.n674 VSSD 0.030737f
C2156 VDDD.n675 VSSD 0.016743f
C2157 VDDD.n676 VSSD 0.014164f
C2158 VDDD.t2038 VSSD 0.023382f
C2159 VDDD.n679 VSSD 0.021149f
C2160 VDDD.n680 VSSD 0.016544f
C2161 VDDD.t2065 VSSD 0.081647f
C2162 VDDD.n723 VSSD 0.038045f
C2163 VDDD.n749 VSSD 0.33981f
C2164 VDDD.t2009 VSSD 0.081647f
C2165 VDDD.n759 VSSD 0.038136f
C2166 VDDD.t1796 VSSD 0.058119f
C2167 VDDD.t2063 VSSD 0.011988f
C2168 VDDD.n775 VSSD 0.030737f
C2169 VDDD.n776 VSSD 0.016743f
C2170 VDDD.t2031 VSSD 0.011988f
C2171 VDDD.n778 VSSD 0.030737f
C2172 VDDD.n779 VSSD 0.016743f
C2173 VDDD.n780 VSSD 0.013794f
C2174 VDDD.n784 VSSD 0.02077f
C2175 VDDD.t2077 VSSD 0.042046f
C2176 VDDD.n786 VSSD 0.063281f
C2177 VDDD.n787 VSSD 0.013486f
C2178 VDDD.n797 VSSD 0.019389f
C2179 VDDD.n798 VSSD 0.016432f
C2180 VDDD.n799 VSSD 0.01711f
C2181 VDDD.n800 VSSD 0.01206f
C2182 VDDD.n803 VSSD 0.021637f
C2183 VDDD.n804 VSSD 0.039466f
C2184 VDDD.n805 VSSD 0.026923f
C2185 VDDD.t2105 VSSD 0.042035f
C2186 VDDD.n806 VSSD 0.070387f
C2187 VDDD.n807 VSSD 0.014424f
C2188 VDDD.n809 VSSD 0.025461f
C2189 VDDD.n810 VSSD 0.062674f
C2190 VDDD.t1112 VSSD 0.077846f
C2191 VDDD.t994 VSSD 0.027787f
C2192 VDDD.t1310 VSSD 0.039453f
C2193 VDDD.t1289 VSSD 0.050271f
C2194 VDDD.t356 VSSD 0.030969f
C2195 VDDD.t1476 VSSD 0.040726f
C2196 VDDD.t1287 VSSD 0.040726f
C2197 VDDD.t371 VSSD 0.036059f
C2198 VDDD.t1701 VSSD 0.039241f
C2199 VDDD.t1901 VSSD 0.033302f
C2200 VDDD.t1843 VSSD 0.041786f
C2201 VDDD.t1259 VSSD 0.050059f
C2202 VDDD.t811 VSSD 0.050271f
C2203 VDDD.t1230 VSSD 0.050695f
C2204 VDDD.t583 VSSD 0.031181f
C2205 VDDD.t1192 VSSD 0.019727f
C2206 VDDD.t423 VSSD 0.024181f
C2207 VDDD.t1442 VSSD 0.035635f
C2208 VDDD.t421 VSSD 0.02206f
C2209 VDDD.t1699 VSSD 0.017817f
C2210 VDDD.t1957 VSSD 0.017817f
C2211 VDDD.t190 VSSD 0.017817f
C2212 VDDD.t1959 VSSD 0.013787f
C2213 VDDD.n811 VSSD 0.021059f
C2214 VDDD.n815 VSSD 0.010242f
C2215 VDDD.n828 VSSD 0.012412f
C2216 VDDD.n861 VSSD 0.012549f
C2217 VDDD.t2080 VSSD 0.032941f
C2218 VDDD.n877 VSSD 0.013558f
C2219 VDDD.n908 VSSD 0.013708f
C2220 VDDD.t1199 VSSD 0.019514f
C2221 VDDD.t927 VSSD 0.021424f
C2222 VDDD.t365 VSSD 0.014212f
C2223 VDDD.t1955 VSSD 0.018242f
C2224 VDDD.t359 VSSD 0.017817f
C2225 VDDD.t923 VSSD 0.018242f
C2226 VDDD.t434 VSSD 0.017817f
C2227 VDDD.t1197 VSSD 0.018242f
C2228 VDDD.t432 VSSD 0.017817f
C2229 VDDD.t925 VSSD 0.018242f
C2230 VDDD.t1530 VSSD 0.030332f
C2231 VDDD.t436 VSSD 0.036484f
C2232 VDDD.t1526 VSSD 0.027363f
C2233 VDDD.t1306 VSSD 0.018242f
C2234 VDDD.t430 VSSD 0.017817f
C2235 VDDD.t1308 VSSD 0.018242f
C2236 VDDD.t1528 VSSD 0.027787f
C2237 VDDD.t1409 VSSD 0.036059f
C2238 VDDD.t385 VSSD 0.035635f
C2239 VDDD.t1899 VSSD 0.03415f
C2240 VDDD.t715 VSSD 0.022908f
C2241 VDDD.t543 VSSD 0.017817f
C2242 VDDD.t1556 VSSD 0.017817f
C2243 VDDD.t1102 VSSD 0.024817f
C2244 VDDD.t219 VSSD 0.039029f
C2245 VDDD.t243 VSSD 0.020999f
C2246 VDDD.t931 VSSD 0.017817f
C2247 VDDD.t670 VSSD 0.040514f
C2248 VDDD.t1558 VSSD 0.024181f
C2249 VDDD.t672 VSSD 0.017817f
C2250 VDDD.t411 VSSD 0.020575f
C2251 VDDD.t1519 VSSD 0.018242f
C2252 VDDD.t114 VSSD 0.029696f
C2253 VDDD.t222 VSSD 0.020999f
C2254 VDDD.t79 VSSD 0.020999f
C2255 VDDD.t1101 VSSD 0.034999f
C2256 VDDD.t817 VSSD 0.026302f
C2257 VDDD.t668 VSSD 0.027363f
C2258 VDDD.t929 VSSD 0.049847f
C2259 VDDD.t220 VSSD 0.029696f
C2260 VDDD.t884 VSSD 0.017817f
C2261 VDDD.t1521 VSSD 0.020999f
C2262 VDDD.t410 VSSD 0.013787f
C2263 VDDD.t795 VSSD 0.015909f
C2264 VDDD.n909 VSSD 0.032725f
C2265 VDDD.t112 VSSD 0.04518f
C2266 VDDD.t1965 VSSD 0.031605f
C2267 VDDD.t1012 VSSD 0.019514f
C2268 VDDD.t799 VSSD 0.024393f
C2269 VDDD.t440 VSSD 0.032453f
C2270 VDDD.t41 VSSD 0.022484f
C2271 VDDD.t1953 VSSD 0.017817f
C2272 VDDD.t1897 VSSD 0.019514f
C2273 VDDD.t1604 VSSD 0.038605f
C2274 VDDD.t1879 VSSD 0.039029f
C2275 VDDD.t416 VSSD 0.029696f
C2276 VDDD.t144 VSSD 0.019514f
C2277 VDDD.t1266 VSSD 0.020575f
C2278 VDDD.t1674 VSSD 0.020999f
C2279 VDDD.t1939 VSSD 0.037968f
C2280 VDDD.t713 VSSD 0.033514f
C2281 VDDD.t557 VSSD 0.020575f
C2282 VDDD.t1660 VSSD 0.020999f
C2283 VDDD.t442 VSSD 0.022484f
C2284 VDDD.t1603 VSSD 0.036059f
C2285 VDDD.t1886 VSSD 0.019302f
C2286 VDDD.t1940 VSSD 0.022484f
C2287 VDDD.t1896 VSSD 0.021424f
C2288 VDDD.t259 VSSD 0.018242f
C2289 VDDD.t451 VSSD 0.035635f
C2290 VDDD.t9 VSSD 0.040726f
C2291 VDDD.t1666 VSSD 0.027787f
C2292 VDDD.t1888 VSSD 0.017817f
C2293 VDDD.t1400 VSSD 0.017817f
C2294 VDDD.t1884 VSSD 0.045604f
C2295 VDDD.t11 VSSD 0.054725f
C2296 VDDD.t7 VSSD 0.015696f
C2297 VDDD.t1015 VSSD 0.058543f
C2298 VDDD.t447 VSSD 0.032878f
C2299 VDDD.t1066 VSSD 0.017817f
C2300 VDDD.t943 VSSD 0.046029f
C2301 VDDD.t1579 VSSD 0.06024f
C2302 VDDD.t1535 VSSD 0.017817f
C2303 VDDD.t642 VSSD 0.017817f
C2304 VDDD.t755 VSSD 0.022908f
C2305 VDDD.t445 VSSD 0.02609f
C2306 VDDD.t726 VSSD 0.036059f
C2307 VDDD.t425 VSSD 0.019514f
C2308 VDDD.t17 VSSD 0.01909f
C2309 VDDD.t1870 VSSD 0.019727f
C2310 VDDD.t617 VSSD 0.022908f
C2311 VDDD.t1933 VSSD 0.038817f
C2312 VDDD.t1534 VSSD 0.020787f
C2313 VDDD.t1253 VSSD 0.018242f
C2314 VDDD.t105 VSSD 0.020575f
C2315 VDDD.t1916 VSSD 0.020999f
C2316 VDDD.t1267 VSSD 0.029696f
C2317 VDDD.t684 VSSD 0.034999f
C2318 VDDD.t685 VSSD 0.027787f
C2319 VDDD.t1593 VSSD 0.019514f
C2320 VDDD.t1213 VSSD 0.020575f
C2321 VDDD.t121 VSSD 0.037544f
C2322 VDDD.t1402 VSSD 0.048786f
C2323 VDDD.t682 VSSD 0.020999f
C2324 VDDD.t598 VSSD 0.017817f
C2325 VDDD.t188 VSSD 0.019514f
C2326 VDDD.t986 VSSD 0.03415f
C2327 VDDD.t103 VSSD 0.01909f
C2328 VDDD.t1523 VSSD 0.024393f
C2329 VDDD.n910 VSSD 0.038452f
C2330 VDDD.t2069 VSSD 0.023382f
C2331 VDDD.n915 VSSD 0.02096f
C2332 VDDD.t2050 VSSD 0.023382f
C2333 VDDD.n937 VSSD 0.021149f
C2334 VDDD.t1993 VSSD 0.011988f
C2335 VDDD.n939 VSSD 0.030737f
C2336 VDDD.n940 VSSD 0.016743f
C2337 VDDD.t2101 VSSD 0.011988f
C2338 VDDD.n942 VSSD 0.030737f
C2339 VDDD.n943 VSSD 0.016743f
C2340 VDDD.n944 VSSD 0.014113f
C2341 VDDD.n948 VSSD 0.018289f
C2342 VDDD.n949 VSSD 0.016338f
C2343 VDDD.n950 VSSD 0.019389f
C2344 VDDD.n956 VSSD 0.010653f
C2345 VDDD.n958 VSSD 0.013224f
C2346 VDDD.n985 VSSD 0.01681f
C2347 VDDD.n990 VSSD 0.012221f
C2348 VDDD.n1000 VSSD 0.011873f
C2349 VDDD.n1037 VSSD 0.017188f
C2350 VDDD.n1038 VSSD 0.017188f
C2351 VDDD.n1039 VSSD 0.013558f
C2352 VDDD.n1040 VSSD 0.036216f
C2353 VDDD.n1073 VSSD 0.013708f
C2354 VDDD.n1083 VSSD 0.011236f
C2355 VDDD.n1092 VSSD 0.19393f
C2356 VDDD.n1093 VSSD 0.676845f
C2357 VDDD.n1095 VSSD 0.199537f
C2358 VDDD.n1101 VSSD 0.021474f
C2359 VDDD.t2083 VSSD 0.023382f
C2360 VDDD.n1117 VSSD 0.019449f
C2361 VDDD.t2106 VSSD 0.023382f
C2362 VDDD.n1132 VSSD 0.021149f
C2363 VDDD.n1142 VSSD 0.138631f
C2364 VDDD.t1980 VSSD 0.081647f
C2365 VDDD.n1150 VSSD 0.037547f
C2366 VDDD.n1153 VSSD 0.014872f
C2367 VDDD.t738 VSSD 0.023333f
C2368 VDDD.t1575 VSSD 0.018878f
C2369 VDDD.t1569 VSSD 0.02312f
C2370 VDDD.t1571 VSSD 0.035635f
C2371 VDDD.t196 VSSD 0.022484f
C2372 VDDD.t1173 VSSD 0.017817f
C2373 VDDD.t148 VSSD 0.030969f
C2374 VDDD.t192 VSSD 0.019727f
C2375 VDDD.t150 VSSD 0.019514f
C2376 VDDD.t1631 VSSD 0.014212f
C2377 VDDD.t194 VSSD 0.017817f
C2378 VDDD.t1389 VSSD 0.017817f
C2379 VDDD.t152 VSSD 0.025454f
C2380 VDDD.t1249 VSSD 0.035635f
C2381 VDDD.t146 VSSD 0.031181f
C2382 VDDD.t1949 VSSD 0.032878f
C2383 VDDD.t844 VSSD 0.035635f
C2384 VDDD.t1683 VSSD 0.034575f
C2385 VDDD.t1695 VSSD 0.040726f
C2386 VDDD.t1162 VSSD 0.020575f
C2387 VDDD.t397 VSSD 0.032878f
C2388 VDDD.t1324 VSSD 0.039453f
C2389 VDDD.t1682 VSSD 0.039241f
C2390 VDDD.t843 VSSD 0.036059f
C2391 VDDD.t1107 VSSD 0.040726f
C2392 VDDD.t305 VSSD 0.040726f
C2393 VDDD.t1641 VSSD 0.024817f
C2394 VDDD.t487 VSSD 0.045604f
C2395 VDDD.t1103 VSSD 0.056422f
C2396 VDDD.t1105 VSSD 0.04921f
C2397 VDDD.t1030 VSSD 0.058543f
C2398 VDDD.t1071 VSSD 0.234173f
C2399 VDDD.t1041 VSSD 0.234173f
C2400 VDDD.n1155 VSSD 0.057543f
C2401 VDDD.t2030 VSSD 0.081647f
C2402 VDDD.t1994 VSSD 0.081647f
C2403 VDDD.n1159 VSSD 0.075101f
C2404 VDDD.n1161 VSSD 0.014343f
C2405 VDDD.t2045 VSSD 0.081647f
C2406 VDDD.t2006 VSSD 0.081647f
C2407 VDDD.n1166 VSSD 0.075101f
C2408 VDDD.n1168 VSSD 0.014343f
C2409 VDDD.t2096 VSSD 0.011988f
C2410 VDDD.n1172 VSSD 0.030737f
C2411 VDDD.n1173 VSSD 0.016743f
C2412 VDDD.t2058 VSSD 0.011988f
C2413 VDDD.n1175 VSSD 0.030737f
C2414 VDDD.n1176 VSSD 0.016743f
C2415 VDDD.n1178 VSSD 0.014115f
C2416 VDDD.n1182 VSSD 0.013875f
C2417 VDDD.n1183 VSSD 0.014343f
C2418 VDDD.n1184 VSSD 0.014343f
C2419 VDDD.n1188 VSSD 0.014343f
C2420 VDDD.n1189 VSSD 0.014343f
C2421 VDDD.n1190 VSSD 0.010523f
C2422 VDDD.n1193 VSSD 0.010991f
C2423 VDDD.n1194 VSSD 0.014343f
C2424 VDDD.n1195 VSSD 0.013875f
C2425 VDDD.n1202 VSSD 0.013875f
C2426 VDDD.n1203 VSSD 0.014343f
C2427 VDDD.n1204 VSSD 0.014343f
C2428 VDDD.n1208 VSSD 0.014343f
C2429 VDDD.n1209 VSSD 0.014343f
C2430 VDDD.n1210 VSSD 0.010523f
C2431 VDDD.n1213 VSSD 0.010991f
C2432 VDDD.n1214 VSSD 0.014343f
C2433 VDDD.n1215 VSSD 0.013875f
C2434 VDDD.n1222 VSSD 0.019206f
C2435 VDDD.n1224 VSSD 0.012594f
C2436 VDDD.n1237 VSSD 0.138631f
C2437 VDDD.n1243 VSSD 0.016544f
C2438 VDDD.t2095 VSSD 0.041456f
C2439 VDDD.n1244 VSSD 0.017377f
C2440 VDDD.t2108 VSSD 0.023382f
C2441 VDDD.n1247 VSSD 0.033916f
C2442 VDDD.n1259 VSSD 0.017377f
C2443 VDDD.t2088 VSSD 0.011988f
C2444 VDDD.n1262 VSSD 0.030737f
C2445 VDDD.n1263 VSSD 0.015201f
C2446 VDDD.t2043 VSSD 0.032941f
C2447 VDDD.n1281 VSSD 0.138631f
C2448 VDDD.n1293 VSSD 0.011885f
C2449 VDDD.t56 VSSD 0.058119f
C2450 VDDD.t2026 VSSD 0.011988f
C2451 VDDD.n1298 VSSD 0.030737f
C2452 VDDD.n1299 VSSD 0.016743f
C2453 VDDD.t2090 VSSD 0.011988f
C2454 VDDD.n1301 VSSD 0.030737f
C2455 VDDD.n1302 VSSD 0.016743f
C2456 VDDD.n1303 VSSD 0.014164f
C2457 VDDD.n1330 VSSD 0.012503f
C2458 VDDD.n1335 VSSD 0.014424f
C2459 VDDD.t2049 VSSD 0.042035f
C2460 VDDD.n1337 VSSD 0.070387f
C2461 VDDD.n1338 VSSD 0.018492f
C2462 VDDD.t2040 VSSD 0.023382f
C2463 VDDD.n1386 VSSD 0.011427f
C2464 VDDD.n1387 VSSD 0.012663f
C2465 VDDD.n1389 VSSD 0.021149f
C2466 VDDD.n1397 VSSD 0.015516f
C2467 VDDD.t1050 VSSD 0.058119f
C2468 VDDD.t955 VSSD 0.016333f
C2469 VDDD.n1437 VSSD 0.013276f
C2470 VDDD.n1438 VSSD 0.010513f
C2471 VDDD.t2023 VSSD 0.011988f
C2472 VDDD.n1440 VSSD 0.030737f
C2473 VDDD.n1441 VSSD 0.016743f
C2474 VDDD.t1991 VSSD 0.011988f
C2475 VDDD.n1443 VSSD 0.030737f
C2476 VDDD.n1444 VSSD 0.016743f
C2477 VDDD.n1445 VSSD 0.013922f
C2478 VDDD.t2079 VSSD 0.023382f
C2479 VDDD.n1450 VSSD 0.011511f
C2480 VDDD.n1454 VSSD 0.011873f
C2481 VDDD.n1468 VSSD 0.011152f
C2482 VDDD.n1473 VSSD 0.013033f
C2483 VDDD.n1474 VSSD 0.01841f
C2484 VDDD.n1481 VSSD 0.013175f
C2485 VDDD.n1482 VSSD 0.021474f
C2486 VDDD.t595 VSSD 0.022696f
C2487 VDDD.t1540 VSSD 0.045604f
C2488 VDDD.t1009 VSSD 0.017817f
C2489 VDDD.t1676 VSSD 0.028211f
C2490 VDDD.t593 VSSD 0.027575f
C2491 VDDD.t1883 VSSD 0.027787f
C2492 VDDD.t1413 VSSD 0.018242f
C2493 VDDD.t853 VSSD 0.017817f
C2494 VDDD.t1417 VSSD 0.020999f
C2495 VDDD.t1697 VSSD 0.045604f
C2496 VDDD.t1430 VSSD 0.041786f
C2497 VDDD.t279 VSSD 0.017817f
C2498 VDDD.t1225 VSSD 0.020575f
C2499 VDDD.t635 VSSD 0.022908f
C2500 VDDD.t1415 VSSD 0.029696f
C2501 VDDD.t852 VSSD 0.017817f
C2502 VDDD.t247 VSSD 0.020999f
C2503 VDDD.t1882 VSSD 0.018242f
C2504 VDDD.t810 VSSD 0.019514f
C2505 VDDD.t213 VSSD 0.020999f
C2506 VDDD.t1245 VSSD 0.045817f
C2507 VDDD.t1478 VSSD 0.052604f
C2508 VDDD.t742 VSSD 0.020575f
C2509 VDDD.t1909 VSSD 0.017817f
C2510 VDDD.t367 VSSD 0.021848f
C2511 VDDD.t1724 VSSD 0.028848f
C2512 VDDD.t1712 VSSD 0.040514f
C2513 VDDD.t154 VSSD 0.055362f
C2514 VDDD.t989 VSSD 0.056634f
C2515 VDDD.t1722 VSSD 0.038605f
C2516 VDDD.t780 VSSD 0.031605f
C2517 VDDD.t1383 VSSD 0.015909f
C2518 VDDD.t1082 VSSD 0.039877f
C2519 VDDD.t654 VSSD 0.024817f
C2520 VDDD.t337 VSSD 0.040726f
C2521 VDDD.t1385 VSSD 0.037968f
C2522 VDDD.t1504 VSSD 0.017817f
C2523 VDDD.t1908 VSSD 0.018242f
C2524 VDDD.t1506 VSSD 0.018242f
C2525 VDDD.t1485 VSSD 0.018242f
C2526 VDDD.t1316 VSSD 0.020999f
C2527 VDDD.t1377 VSSD 0.018242f
C2528 VDDD.t235 VSSD 0.030969f
C2529 VDDD.t183 VSSD 0.02906f
C2530 VDDD.t315 VSSD 0.018242f
C2531 VDDD.t233 VSSD 0.020575f
C2532 VDDD.t660 VSSD 0.018242f
C2533 VDDD.t179 VSSD 0.023333f
C2534 VDDD.t181 VSSD 0.024605f
C2535 VDDD.t611 VSSD 0.01803f
C2536 VDDD.t963 VSSD 0.020999f
C2537 VDDD.t142 VSSD 0.018242f
C2538 VDDD.t967 VSSD 0.019514f
C2539 VDDD.t414 VSSD 0.018242f
C2540 VDDD.t1500 VSSD 0.025878f
C2541 VDDD.t237 VSSD 0.036484f
C2542 VDDD.t965 VSSD 0.030757f
C2543 VDDD.t1725 VSSD 0.018242f
C2544 VDDD.t1498 VSSD 0.017817f
C2545 VDDD.t569 VSSD 0.018242f
C2546 VDDD.t1314 VSSD 0.019302f
C2547 VDDD.t1554 VSSD 0.034999f
C2548 VDDD.t1496 VSSD 0.022484f
C2549 VDDD.t1494 VSSD 0.021424f
C2550 VDDD.t621 VSSD 0.018242f
C2551 VDDD.t854 VSSD 0.017605f
C2552 VDDD.t828 VSSD 0.021424f
C2553 VDDD.t623 VSSD 0.035635f
C2554 VDDD.t1678 VSSD 0.01803f
C2555 VDDD.t241 VSSD 0.042058f
C2556 VDDD.n1483 VSSD 0.01268f
C2557 VDDD.n1487 VSSD 0.016621f
C2558 VDDD.n1488 VSSD 0.013558f
C2559 VDDD.n1490 VSSD 0.01426f
C2560 VDDD.n1491 VSSD 0.013193f
C2561 VDDD.n1492 VSSD 0.011265f
C2562 VDDD.n1493 VSSD 0.018357f
C2563 VDDD.n1517 VSSD 0.19393f
C2564 VDDD.n1533 VSSD 0.011885f
C2565 VDDD.t2004 VSSD 0.032941f
C2566 VDDD.t2081 VSSD 0.032941f
C2567 VDDD.n1535 VSSD 0.018563f
C2568 VDDD.n1536 VSSD 0.018563f
C2569 VDDD.n1537 VSSD 0.031352f
C2570 VDDD.n1541 VSSD 0.032409f
C2571 VDDD.n1542 VSSD 0.032409f
C2572 VDDD.n1543 VSSD 0.087162f
C2573 VDDD.n1561 VSSD 0.216356f
C2574 VDDD.n1562 VSSD 0.676845f
C2575 VDDD.n1564 VSSD 0.277262f
C2576 VDDD.n1569 VSSD 0.029437f
C2577 VDDD.t2003 VSSD 0.040409f
C2578 VDDD.n1570 VSSD 0.018019f
C2579 VDDD.n1573 VSSD 0.011873f
C2580 VDDD.t2061 VSSD 0.042267f
C2581 VDDD.n1597 VSSD 0.076191f
C2582 VDDD.n1598 VSSD 0.022234f
C2583 VDDD.n1600 VSSD 0.014449f
C2584 VDDD.n1601 VSSD 0.013558f
C2585 VDDD.n1633 VSSD 0.214062f
C2586 VDDD.t2044 VSSD 0.032941f
C2587 VDDD.n1644 VSSD 0.012305f
C2588 VDDD.t1512 VSSD 0.015909f
C2589 VDDD.n1655 VSSD 0.018492f
C2590 VDDD.t2100 VSSD 0.042035f
C2591 VDDD.n1656 VSSD 0.070387f
C2592 VDDD.n1657 VSSD 0.014424f
C2593 VDDD.n1662 VSSD 0.011866f
C2594 VDDD.t484 VSSD 0.058119f
C2595 VDDD.t1989 VSSD 0.011988f
C2596 VDDD.n1692 VSSD 0.030737f
C2597 VDDD.n1693 VSSD 0.016743f
C2598 VDDD.t2053 VSSD 0.011988f
C2599 VDDD.n1695 VSSD 0.030737f
C2600 VDDD.n1696 VSSD 0.016743f
C2601 VDDD.n1697 VSSD 0.014164f
C2602 VDDD.t2012 VSSD 0.023382f
C2603 VDDD.n1702 VSSD 0.016544f
C2604 VDDD.t2032 VSSD 0.081647f
C2605 VDDD.n1709 VSSD 0.037547f
C2606 VDDD.t2109 VSSD 0.081647f
C2607 VDDD.n1730 VSSD 0.038136f
C2608 VDDD.n1735 VSSD 0.010774f
C2609 VDDD.n1785 VSSD 0.011502f
C2610 VDDD.n1790 VSSD 0.013033f
C2611 VDDD.n1791 VSSD 0.021149f
C2612 VDDD.n1793 VSSD 0.017775f
C2613 VDDD.n1794 VSSD 0.042483f
C2614 VDDD.t1739 VSSD 0.028211f
C2615 VDDD.t1605 VSSD 0.032878f
C2616 VDDD.t1342 VSSD 0.05218f
C2617 VDDD.t463 VSSD 0.063422f
C2618 VDDD.t399 VSSD 0.040726f
C2619 VDDD.t1344 VSSD 0.040726f
C2620 VDDD.t612 VSSD 0.030332f
C2621 VDDD.t1778 VSSD 0.018242f
C2622 VDDD.t1459 VSSD 0.026726f
C2623 VDDD.t1355 VSSD 0.062786f
C2624 VDDD.t307 VSSD 0.062361f
C2625 VDDD.t231 VSSD 0.042423f
C2626 VDDD.t1458 VSSD 0.028848f
C2627 VDDD.t345 VSSD 0.040514f
C2628 VDDD.t906 VSSD 0.076149f
C2629 VDDD.t1456 VSSD 0.074452f
C2630 VDDD.t577 VSSD 0.018242f
C2631 VDDD.t520 VSSD 0.013787f
C2632 VDDD.t354 VSSD 0.04815f
C2633 VDDD.t766 VSSD 0.036484f
C2634 VDDD.t764 VSSD 0.036484f
C2635 VDDD.t1607 VSSD 0.031181f
C2636 VDDD.t1975 VSSD 0.015909f
C2637 VDDD.t1047 VSSD 0.058543f
C2638 VDDD.t1468 VSSD 0.031605f
C2639 VDDD.t1538 VSSD 0.01909f
C2640 VDDD.t514 VSSD 0.056634f
C2641 VDDD.t1729 VSSD 0.074876f
C2642 VDDD.t1332 VSSD 0.040514f
C2643 VDDD.t601 VSSD 0.048786f
C2644 VDDD.t1423 VSSD 0.01909f
C2645 VDDD.t25 VSSD 0.028635f
C2646 VDDD.t27 VSSD 0.031181f
C2647 VDDD.t770 VSSD 0.018242f
C2648 VDDD.t29 VSSD 0.020999f
C2649 VDDD.t1537 VSSD 0.018242f
C2650 VDDD.t35 VSSD 0.018242f
C2651 VDDD.t1333 VSSD 0.018242f
C2652 VDDD.t352 VSSD 0.017817f
C2653 VDDD.t625 VSSD 0.018242f
C2654 VDDD.t648 VSSD 0.021211f
C2655 VDDD.t652 VSSD 0.019939f
C2656 VDDD.t732 VSSD 0.018242f
C2657 VDDD.t768 VSSD 0.017817f
C2658 VDDD.t1686 VSSD 0.018242f
C2659 VDDD.t646 VSSD 0.035211f
C2660 VDDD.t650 VSSD 0.028635f
C2661 VDDD.t740 VSSD 0.018242f
C2662 VDDD.t346 VSSD 0.017817f
C2663 VDDD.t627 VSSD 0.018242f
C2664 VDDD.t350 VSSD 0.026302f
C2665 VDDD.t1977 VSSD 0.019302f
C2666 VDDD.t1609 VSSD 0.035211f
C2667 VDDD.t348 VSSD 0.025878f
C2668 VDDD.n1795 VSSD 0.021898f
C2669 VDDD.n1796 VSSD 0.013589f
C2670 VDDD.n1807 VSSD 0.011199f
C2671 VDDD.n1809 VSSD 0.011507f
C2672 VDDD.t1997 VSSD 0.081647f
C2673 VDDD.n1824 VSSD 0.037275f
C2674 VDDD.t1999 VSSD 0.011988f
C2675 VDDD.n1828 VSSD 0.030737f
C2676 VDDD.n1829 VSSD 0.016743f
C2677 VDDD.n1832 VSSD 0.010792f
C2678 VDDD.n1833 VSSD 0.019362f
C2679 VDDD.n1882 VSSD 0.216356f
C2680 VDDD.n1883 VSSD 0.214062f
C2681 VDDD.n1887 VSSD 0.011504f
C2682 VDDD.t997 VSSD 0.058119f
C2683 VDDD.t2087 VSSD 0.011988f
C2684 VDDD.n1891 VSSD 0.030737f
C2685 VDDD.n1892 VSSD 0.016743f
C2686 VDDD.t2017 VSSD 0.011988f
C2687 VDDD.n1894 VSSD 0.030737f
C2688 VDDD.n1895 VSSD 0.016743f
C2689 VDDD.n1896 VSSD 0.014164f
C2690 VDDD.n1900 VSSD 0.013262f
C2691 VDDD.n1902 VSSD 0.011542f
C2692 VDDD.t2054 VSSD 0.023588f
C2693 VDDD.n1933 VSSD 0.04098f
C2694 VDDD.n1934 VSSD 0.023515f
C2695 VDDD.n1935 VSSD 0.019829f
C2696 VDDD.n1936 VSSD 0.014261f
C2697 VDDD.t2076 VSSD 0.033523f
C2698 VDDD.n1937 VSSD 0.050791f
C2699 VDDD.n1938 VSSD 0.032898f
C2700 VDDD.n1940 VSSD 0.018199f
C2701 VDDD.t2039 VSSD 0.081647f
C2702 VDDD.n1972 VSSD 0.038136f
C2703 VDDD.n1975 VSSD 0.010064f
C2704 VDDD.n1977 VSSD 0.012867f
C2705 VDDD.t2042 VSSD 0.041456f
C2706 VDDD.n1978 VSSD 0.012305f
C2707 VDDD.n1980 VSSD 0.013033f
C2708 VDDD.t1091 VSSD 0.058119f
C2709 VDDD.n1982 VSSD 0.020665f
C2710 VDDD.t2086 VSSD 0.011988f
C2711 VDDD.n1984 VSSD 0.030737f
C2712 VDDD.n1985 VSSD 0.016743f
C2713 VDDD.t2008 VSSD 0.011988f
C2714 VDDD.n1988 VSSD 0.030737f
C2715 VDDD.n1989 VSSD 0.016743f
C2716 VDDD.t1979 VSSD 0.011988f
C2717 VDDD.n1991 VSSD 0.030737f
C2718 VDDD.n1992 VSSD 0.016743f
C2719 VDDD.n1993 VSSD 0.014164f
C2720 VDDD.t2102 VSSD 0.081647f
C2721 VDDD.n2008 VSSD 0.038136f
C2722 VDDD.n2020 VSSD 0.024579f
C2723 VDDD.n2021 VSSD 0.055038f
C2724 VDDD.t1379 VSSD 0.039029f
C2725 VDDD.t1153 VSSD 0.017817f
C2726 VDDD.t1381 VSSD 0.02312f
C2727 VDDD.t89 VSSD 0.050483f
C2728 VDDD.t395 VSSD 0.040726f
C2729 VDDD.t1387 VSSD 0.040726f
C2730 VDDD.t779 VSSD 0.036059f
C2731 VDDD.t1891 VSSD 0.032029f
C2732 VDDD.t475 VSSD 0.020999f
C2733 VDDD.t1720 VSSD 0.048998f
C2734 VDDD.t303 VSSD 0.062361f
C2735 VDDD.t383 VSSD 0.050271f
C2736 VDDD.t1890 VSSD 0.041362f
C2737 VDDD.t778 VSSD 0.028848f
C2738 VDDD.t801 VSSD 0.076149f
C2739 VDDD.t1688 VSSD 0.074452f
C2740 VDDD.t1448 VSSD 0.031605f
C2741 VDDD.t1770 VSSD 0.01909f
C2742 VDDD.t1799 VSSD 0.097996f
C2743 VDDD.n2022 VSSD 0.024534f
C2744 VDDD.n2023 VSSD 0.018467f
C2745 VDDD.n2026 VSSD 0.017278f
C2746 VDDD.t1983 VSSD 0.081647f
C2747 VDDD.t2025 VSSD 0.023382f
C2748 VDDD.n2055 VSSD 0.023952f
C2749 VDDD.n2056 VSSD 0.012594f
C2750 VDDD.n2076 VSSD 0.011438f
C2751 VDDD.t2066 VSSD 0.012068f
C2752 VDDD.n2078 VSSD 0.019643f
C2753 VDDD.n2079 VSSD 0.015041f
C2754 VDDD.t2114 VSSD 0.081647f
C2755 VDDD.n2108 VSSD 0.038136f
C2756 VDDD.t1992 VSSD 0.081647f
C2757 VDDD.n2131 VSSD 0.036549f
C2758 VDDD.n2137 VSSD 0.014872f
C2759 VDDD.n2143 VSSD 0.010064f
C2760 VDDD.n2146 VSSD 0.017532f
C2761 VDDD.n2147 VSSD 0.022614f
C2762 VDDD.n2148 VSSD 0.013484f
C2763 VDDD.n2155 VSSD 0.214062f
C2764 VDDD.t2070 VSSD 0.011988f
C2765 VDDD.n2161 VSSD 0.030737f
C2766 VDDD.n2162 VSSD 0.016743f
C2767 VDDD.n2163 VSSD 0.01603f
C2768 VDDD.t2073 VSSD 0.081647f
C2769 VDDD.n2170 VSSD 0.038136f
C2770 VDDD.n2197 VSSD 0.012922f
C2771 VDDD.n2198 VSSD 0.03791f
C2772 VDDD.n2199 VSSD 0.012594f
C2773 VDDD.n2216 VSSD 0.010064f
C2774 VDDD.n2217 VSSD 0.012867f
C2775 VDDD.t2110 VSSD 0.041456f
C2776 VDDD.n2218 VSSD 0.058912f
C2777 VDDD.n2219 VSSD 0.017024f
C2778 VDDD.n2223 VSSD 0.023376f
C2779 VDDD.n2224 VSSD 0.022614f
C2780 VDDD.n2225 VSSD 0.012305f
C2781 VDDD.n2226 VSSD 0.016441f
C2782 VDDD.t2015 VSSD 0.081647f
C2783 VDDD.t1985 VSSD 0.081647f
C2784 VDDD.n2231 VSSD 0.075101f
C2785 VDDD.n2233 VSSD 0.014343f
C2786 VDDD.t2033 VSSD 0.081647f
C2787 VDDD.t1996 VSSD 0.081647f
C2788 VDDD.n2238 VSSD 0.075101f
C2789 VDDD.n2240 VSSD 0.014343f
C2790 VDDD.t2082 VSSD 0.011988f
C2791 VDDD.n2244 VSSD 0.030737f
C2792 VDDD.n2245 VSSD 0.016743f
C2793 VDDD.t2051 VSSD 0.011988f
C2794 VDDD.n2247 VSSD 0.030737f
C2795 VDDD.n2248 VSSD 0.016743f
C2796 VDDD.n2250 VSSD 0.014115f
C2797 VDDD.n2254 VSSD 0.013875f
C2798 VDDD.n2255 VSSD 0.014343f
C2799 VDDD.n2256 VSSD 0.014343f
C2800 VDDD.n2260 VSSD 0.014343f
C2801 VDDD.n2261 VSSD 0.014343f
C2802 VDDD.n2262 VSSD 0.010523f
C2803 VDDD.n2265 VSSD 0.010991f
C2804 VDDD.n2266 VSSD 0.014343f
C2805 VDDD.n2267 VSSD 0.013875f
C2806 VDDD.n2274 VSSD 0.013875f
C2807 VDDD.n2275 VSSD 0.014343f
C2808 VDDD.n2276 VSSD 0.014343f
C2809 VDDD.n2280 VSSD 0.014343f
C2810 VDDD.n2281 VSSD 0.014343f
C2811 VDDD.n2282 VSSD 0.010523f
C2812 VDDD.n2285 VSSD 0.010991f
C2813 VDDD.n2286 VSSD 0.014343f
C2814 VDDD.n2287 VSSD 0.013875f
C2815 VDDD.n2291 VSSD 0.020887f
C2816 VDDD.t47 VSSD 0.058543f
C2817 VDDD.t1787 VSSD 0.234173f
C2818 VDDD.t1750 VSSD 0.234173f
C2819 VDDD.n2292 VSSD 0.042127f
C2820 VDDD.t1807 VSSD 0.110935f
C2821 VDDD.t1817 VSSD 0.099693f
C2822 VDDD.t704 VSSD 0.039453f
C2823 VDDD.t751 VSSD 0.063422f
C2824 VDDD.t229 VSSD 0.063422f
C2825 VDDD.t297 VSSD 0.038181f
C2826 VDDD.t702 VSSD 0.020363f
C2827 VDDD.t1880 VSSD 0.036059f
C2828 VDDD.t735 VSSD 0.039241f
C2829 VDDD.t223 VSSD 0.062786f
C2830 VDDD.t1241 VSSD 0.051332f
C2831 VDDD.t1118 VSSD 0.020575f
C2832 VDDD.t43 VSSD 0.040726f
C2833 VDDD.t734 VSSD 0.050695f
C2834 VDDD.t1484 VSSD 0.040514f
C2835 VDDD.t1727 VSSD 0.061513f
C2836 VDDD.t736 VSSD 0.02312f
C2837 VDDD.t1109 VSSD 0.017817f
C2838 VDDD.t797 VSSD 0.015909f
C2839 VDDD.n2293 VSSD 0.046341f
C2840 VDDD.t1767 VSSD 0.093542f
C2841 VDDD.t1276 VSSD 0.078058f
C2842 VDDD.t1830 VSSD 0.017817f
C2843 VDDD.t1280 VSSD 0.046029f
C2844 VDDD.t1302 VSSD 0.063422f
C2845 VDDD.t293 VSSD 0.040726f
C2846 VDDD.t1278 VSSD 0.040726f
C2847 VDDD.t1327 VSSD 0.036059f
C2848 VDDD.t553 VSSD 0.018666f
C2849 VDDD.t753 VSSD 0.062361f
C2850 VDDD.t331 VSSD 0.062361f
C2851 VDDD.t808 VSSD 0.048574f
C2852 VDDD.t1804 VSSD 0.029696f
C2853 VDDD.t554 VSSD 0.022696f
C2854 VDDD.t1326 VSSD 0.040514f
C2855 VDDD.t61 VSSD 0.076149f
C2856 VDDD.t555 VSSD 0.074452f
C2857 VDDD.t631 VSSD 0.024393f
C2858 VDDD.t1024 VSSD 0.042635f
C2859 VDDD.n2294 VSSD 0.058391f
C2860 VDDD.n2295 VSSD 0.028229f
C2861 VDDD.n2296 VSSD 0.011624f
C2862 VDDD.n2299 VSSD 0.022614f
C2863 VDDD.n2300 VSSD 0.017278f
C2864 VDDD.n2301 VSSD 0.058912f
C2865 VDDD.n2302 VSSD 0.017024f
C2866 VDDD.n2335 VSSD 0.214062f
C2867 VDDD.n2336 VSSD 0.277262f
C2868 VDDD.n2357 VSSD 0.010729f
C2869 VDDD.n2359 VSSD 0.012384f
C2870 VDDD.n2360 VSSD 0.031665f
C2871 VDDD.t443 VSSD 0.029696f
C2872 VDDD.t1411 VSSD 0.019514f
C2873 VDDD.t374 VSSD 0.019514f
C2874 VDDD.t832 VSSD 0.043908f
C2875 VDDD.t882 VSSD 0.043908f
C2876 VDDD.t317 VSSD 0.019514f
C2877 VDDD.t1662 VSSD 0.019514f
C2878 VDDD.t1239 VSSD 0.021211f
C2879 VDDD.t757 VSSD 0.021211f
C2880 VDDD.t1203 VSSD 0.019514f
C2881 VDDD.t31 VSSD 0.018242f
C2882 VDDD.t1460 VSSD 0.017817f
C2883 VDDD.t1928 VSSD 0.019514f
C2884 VDDD.t454 VSSD 0.019727f
C2885 VDDD.t749 VSSD 0.020999f
C2886 VDDD.t602 VSSD 0.041786f
C2887 VDDD.t1672 VSSD 0.041786f
C2888 VDDD.t265 VSSD 0.020575f
C2889 VDDD.t1318 VSSD 0.020575f
C2890 VDDD.t77 VSSD 0.029696f
C2891 VDDD.t1393 VSSD 0.029696f
C2892 VDDD.t453 VSSD 0.020999f
C2893 VDDD.t1204 VSSD 0.020999f
C2894 VDDD.t33 VSSD 0.039029f
C2895 VDDD.t1629 VSSD 0.056634f
C2896 VDDD.t1391 VSSD 0.054937f
C2897 VDDD.t575 VSSD 0.019514f
C2898 VDDD.t1561 VSSD 0.013787f
C2899 VDDD.t363 VSSD 0.01909f
C2900 VDDD.t1744 VSSD 0.064695f
C2901 VDDD.t1127 VSSD 0.032878f
C2902 VDDD.t615 VSSD 0.039029f
C2903 VDDD.t245 VSSD 0.015909f
C2904 VDDD.t1298 VSSD 0.071906f
C2905 VDDD.t1121 VSSD 0.056634f
C2906 VDDD.t108 VSSD 0.01909f
C2907 VDDD.t579 VSSD 0.024393f
C2908 VDDD.t1347 VSSD 0.031605f
C2909 VDDD.t1894 VSSD 0.025666f
C2910 VDDD.t63 VSSD 0.029696f
C2911 VDDD.t571 VSSD 0.017817f
C2912 VDDD.t1433 VSSD 0.019514f
C2913 VDDD.t168 VSSD 0.038605f
C2914 VDDD.t1893 VSSD 0.039029f
C2915 VDDD.t1731 VSSD 0.029696f
C2916 VDDD.t1294 VSSD 0.019514f
C2917 VDDD.t143 VSSD 0.020575f
C2918 VDDD.t1668 VSSD 0.020999f
C2919 VDDD.t380 VSSD 0.037968f
C2920 VDDD.t1363 VSSD 0.033514f
C2921 VDDD.t161 VSSD 0.020575f
C2922 VDDD.t313 VSSD 0.020999f
C2923 VDDD.t405 VSSD 0.022484f
C2924 VDDD.t167 VSSD 0.036059f
C2925 VDDD.t662 VSSD 0.019302f
C2926 VDDD.t1735 VSSD 0.022484f
C2927 VDDD.t1432 VSSD 0.021424f
C2928 VDDD.t1670 VSSD 0.018242f
C2929 VDDD.t895 VSSD 0.035635f
C2930 VDDD.t613 VSSD 0.040726f
C2931 VDDD.t1664 VSSD 0.027787f
C2932 VDDD.t664 VSSD 0.017817f
C2933 VDDD.t1304 VSSD 0.017817f
C2934 VDDD.t803 VSSD 0.036271f
C2935 VDDD.n2361 VSSD 0.04418f
C2936 VDDD.n2362 VSSD 0.012358f
C2937 VDDD.n2368 VSSD 0.011873f
C2938 VDDD.n2377 VSSD 0.277262f
C2939 VDDD.n2414 VSSD 0.012633f
C2940 VDDD.n2417 VSSD 0.01426f
C2941 VDDD.n2418 VSSD 0.015583f
C2942 VDDD.n2419 VSSD 0.012314f
C2943 VDDD.t2020 VSSD 0.081647f
C2944 VDDD.n2441 VSSD 0.038136f
C2945 VDDD.n2456 VSSD 0.011873f
C2946 VDDD.n2475 VSSD 0.011873f
C2947 VDDD.n2491 VSSD 0.013974f
C2948 VDDD.n2492 VSSD 0.024656f
C2949 VDDD.t806 VSSD 0.022696f
C2950 VDDD.t1338 VSSD 0.028211f
C2951 VDDD.t1340 VSSD 0.020575f
C2952 VDDD.t311 VSSD 0.017817f
C2953 VDDD.t706 VSSD 0.041786f
C2954 VDDD.t81 VSSD 0.045604f
C2955 VDDD.t875 VSSD 0.020999f
C2956 VDDD.t805 VSSD 0.017817f
C2957 VDDD.t283 VSSD 0.018242f
C2958 VDDD.t959 VSSD 0.022908f
C2959 VDDD.t1945 VSSD 0.017817f
C2960 VDDD.t1190 VSSD 0.017817f
C2961 VDDD.t1944 VSSD 0.022908f
C2962 VDDD.t291 VSSD 0.018242f
C2963 VDDD.t542 VSSD 0.017817f
C2964 VDDD.t198 VSSD 0.020999f
C2965 VDDD.t19 VSSD 0.045604f
C2966 VDDD.t856 VSSD 0.041786f
C2967 VDDD.t275 VSSD 0.017817f
C2968 VDDD.t0 VSSD 0.020575f
C2969 VDDD.t1446 VSSD 0.034575f
C2970 VDDD.t541 VSSD 0.029272f
C2971 VDDD.t1943 VSSD 0.040514f
C2972 VDDD.t912 VSSD 0.076149f
C2973 VDDD.t825 VSSD 0.074452f
C2974 VDDD.t39 VSSD 0.018242f
C2975 VDDD.t1088 VSSD 0.013787f
C2976 VDDD.t1074 VSSD 0.078482f
C2977 VDDD.t1165 VSSD 0.058543f
C2978 VDDD.t1147 VSSD 0.234173f
C2979 VDDD.t1033 VSSD 0.234173f
C2980 VDDD.n2493 VSSD 0.042127f
C2981 VDDD.t2093 VSSD 0.081647f
C2982 VDDD.t2022 VSSD 0.081647f
C2983 VDDD.n2496 VSSD 0.075101f
C2984 VDDD.n2498 VSSD 0.014343f
C2985 VDDD.t2107 VSSD 0.081647f
C2986 VDDD.t2041 VSSD 0.081647f
C2987 VDDD.n2503 VSSD 0.075101f
C2988 VDDD.n2505 VSSD 0.014343f
C2989 VDDD.t2011 VSSD 0.011988f
C2990 VDDD.n2509 VSSD 0.030737f
C2991 VDDD.n2510 VSSD 0.016743f
C2992 VDDD.t2089 VSSD 0.011988f
C2993 VDDD.n2512 VSSD 0.030737f
C2994 VDDD.n2513 VSSD 0.016743f
C2995 VDDD.n2515 VSSD 0.014115f
C2996 VDDD.n2519 VSSD 0.013875f
C2997 VDDD.n2520 VSSD 0.014343f
C2998 VDDD.n2521 VSSD 0.014343f
C2999 VDDD.n2525 VSSD 0.014343f
C3000 VDDD.n2526 VSSD 0.014343f
C3001 VDDD.n2527 VSSD 0.010523f
C3002 VDDD.n2530 VSSD 0.010991f
C3003 VDDD.n2531 VSSD 0.014343f
C3004 VDDD.n2532 VSSD 0.013875f
C3005 VDDD.n2539 VSSD 0.013875f
C3006 VDDD.n2540 VSSD 0.014343f
C3007 VDDD.n2541 VSSD 0.014343f
C3008 VDDD.n2545 VSSD 0.014343f
C3009 VDDD.n2546 VSSD 0.014343f
C3010 VDDD.n2547 VSSD 0.010523f
C3011 VDDD.n2550 VSSD 0.010991f
C3012 VDDD.n2551 VSSD 0.014343f
C3013 VDDD.n2552 VSSD 0.013875f
C3014 VDDD.n2556 VSSD 0.020887f
C3015 VDDD.n2557 VSSD 0.018467f
C3016 VDDD.n2558 VSSD 0.016441f
C3017 VDDD.n2561 VSSD 0.022614f
C3018 VDDD.n2562 VSSD 0.050519f
C3019 VDDD.n2563 VSSD 0.012867f
C3020 VDDD.n2564 VSSD 0.010064f
C3021 VDDD.n2582 VSSD 0.277262f
C3022 VDDD.n2583 VSSD 0.216356f
C3023 VDDD.n2597 VSSD 0.011873f
C3024 VDDD.t2068 VSSD 0.023382f
C3025 VDDD.n2624 VSSD 0.020582f
C3026 VDDD.n2625 VSSD 0.012766f
C3027 VDDD.t2056 VSSD 0.011988f
C3028 VDDD.n2628 VSSD 0.030737f
C3029 VDDD.n2629 VSSD 0.016743f
C3030 VDDD.t1981 VSSD 0.011988f
C3031 VDDD.n2631 VSSD 0.030737f
C3032 VDDD.n2632 VSSD 0.016743f
C3033 VDDD.n2634 VSSD 0.014113f
C3034 VDDD.n2638 VSSD 0.01681f
C3035 VDDD.n2643 VSSD 0.011723f
C3036 VDDD.n2649 VSSD 0.011427f
C3037 VDDD.n2677 VSSD 0.016331f
C3038 VDDD.n2681 VSSD 0.012371f
C3039 VDDD.t1755 VSSD 0.058331f
C3040 VDDD.t1133 VSSD 0.054513f
C3041 VDDD.t1269 VSSD 0.039453f
C3042 VDDD.t1704 VSSD 0.039029f
C3043 VDDD.t389 VSSD 0.039029f
C3044 VDDD.t408 VSSD 0.024393f
C3045 VDDD.t1872 VSSD 0.024393f
C3046 VDDD.t1658 VSSD 0.039029f
C3047 VDDD.t1862 VSSD 0.022908f
C3048 VDDD.t73 VSSD 0.017817f
C3049 VDDD.t301 VSSD 0.017817f
C3050 VDDD.t1373 VSSD 0.019939f
C3051 VDDD.t1719 VSSD 0.021211f
C3052 VDDD.t387 VSSD 0.020787f
C3053 VDDD.t267 VSSD 0.01803f
C3054 VDDD.t666 VSSD 0.018242f
C3055 VDDD.t1625 VSSD 0.039029f
C3056 VDDD.t945 VSSD 0.023757f
C3057 VDDD.t335 VSSD 0.023333f
C3058 VDDD.t428 VSSD 0.039029f
C3059 VDDD.t281 VSSD 0.029696f
C3060 VDDD.t1881 VSSD 0.020575f
C3061 VDDD.t567 VSSD 0.020999f
C3062 VDDD.t1374 VSSD 0.029696f
C3063 VDDD.t1626 VSSD 0.019514f
C3064 VDDD.t1733 VSSD 0.020999f
C3065 VDDD.t268 VSSD 0.039029f
C3066 VDDD.t1450 VSSD 0.03712f
C3067 VDDD.t1717 VSSD 0.035423f
C3068 VDDD.t1646 VSSD 0.024393f
C3069 VDDD.t1627 VSSD 0.032453f
C3070 VDDD.t902 VSSD 0.020363f
C3071 VDDD.t551 VSSD 0.02312f
C3072 VDDD.n2682 VSSD 0.04418f
C3073 VDDD.t469 VSSD 0.036271f
C3074 VDDD.t1513 VSSD 0.017817f
C3075 VDDD.t1184 VSSD 0.017817f
C3076 VDDD.t319 VSSD 0.027787f
C3077 VDDD.t549 VSSD 0.040726f
C3078 VDDD.t1211 VSSD 0.035635f
C3079 VDDD.t401 VSSD 0.018242f
C3080 VDDD.t1466 VSSD 0.021424f
C3081 VDDD.t163 VSSD 0.022484f
C3082 VDDD.t1182 VSSD 0.019302f
C3083 VDDD.t866 VSSD 0.036059f
C3084 VDDD.t1188 VSSD 0.022484f
C3085 VDDD.t321 VSSD 0.020999f
C3086 VDDD.t1648 VSSD 0.020575f
C3087 VDDD.t772 VSSD 0.033514f
C3088 VDDD.t1463 VSSD 0.037968f
C3089 VDDD.t271 VSSD 0.020999f
C3090 VDDD.t582 VSSD 0.020575f
C3091 VDDD.t1407 VSSD 0.019514f
C3092 VDDD.t941 VSSD 0.029696f
C3093 VDDD.t788 VSSD 0.039029f
C3094 VDDD.t867 VSSD 0.038605f
C3095 VDDD.t1464 VSSD 0.019514f
C3096 VDDD.t910 VSSD 0.017817f
C3097 VDDD.t1223 VSSD 0.022484f
C3098 VDDD.t1186 VSSD 0.032453f
C3099 VDDD.t1633 VSSD 0.024393f
C3100 VDDD.t1775 VSSD 0.071906f
C3101 VDDD.t1060 VSSD 0.084633f
C3102 VDDD.n2683 VSSD 0.042118f
C3103 VDDD.n2692 VSSD 0.022758f
C3104 VDDD.n2695 VSSD 0.024266f
C3105 VDDD.n2696 VSSD 0.018019f
C3106 VDDD.n2697 VSSD 0.029567f
C3107 VDDD.n2698 VSSD 0.045757f
C3108 VDDD.n2699 VSSD 0.02465f
C3109 VDDD.n2707 VSSD 0.216356f
C3110 VDDD.n2708 VSSD 0.138631f
C3111 VDDD.n2709 VSSD 0.509672f
C3112 VDDD.n2710 VSSD 0.957816f
C3113 VDDD.n2711 VSSD 0.33981f
C3114 VDDD.n2712 VSSD 0.199537f
C3115 VDDD.n2733 VSSD 0.011542f
C3116 VDDD.n2734 VSSD 0.013262f
C3117 VDDD.n2735 VSSD 0.010729f
C3118 VDDD.n2738 VSSD 0.012384f
C3119 VDDD.n2739 VSSD 0.031665f
C3120 VDDD.t1929 VSSD 0.029696f
C3121 VDDD.t1292 VSSD 0.019514f
C3122 VDDD.t376 VSSD 0.019514f
C3123 VDDD.t378 VSSD 0.043908f
C3124 VDDD.t341 VSSD 0.043908f
C3125 VDDD.t257 VSSD 0.019514f
C3126 VDDD.t1349 VSSD 0.019514f
C3127 VDDD.t285 VSSD 0.021211f
C3128 VDDD.t1394 VSSD 0.021211f
C3129 VDDD.t205 VSSD 0.019514f
C3130 VDDD.t106 VSSD 0.018242f
C3131 VDDD.t1467 VSSD 0.017817f
C3132 VDDD.t413 VSSD 0.019514f
C3133 VDDD.t916 VSSD 0.019727f
C3134 VDDD.t1209 VSSD 0.020999f
C3135 VDDD.t1419 VSSD 0.041786f
C3136 VDDD.t255 VSSD 0.041786f
C3137 VDDD.t277 VSSD 0.020575f
C3138 VDDD.t591 VSSD 0.020575f
C3139 VDDD.t1517 VSSD 0.029696f
C3140 VDDD.t1915 VSSD 0.029696f
C3141 VDDD.t915 VSSD 0.020999f
C3142 VDDD.t701 VSSD 0.020999f
C3143 VDDD.t412 VSSD 0.039029f
C3144 VDDD.t957 VSSD 0.056634f
C3145 VDDD.t1913 VSSD 0.054937f
C3146 VDDD.t361 VSSD 0.019514f
C3147 VDDD.t917 VSSD 0.013787f
C3148 VDDD.t629 VSSD 0.01909f
C3149 VDDD.t1018 VSSD 0.117087f
C3150 VDDD.t207 VSSD 0.032453f
C3151 VDDD.t1221 VSSD 0.024393f
C3152 VDDD.t1085 VSSD 0.019514f
C3153 VDDD.t53 VSSD 0.058543f
C3154 VDDD.t573 VSSD 0.01909f
C3155 VDDD.t158 VSSD 0.013787f
C3156 VDDD.t1573 VSSD 0.019514f
C3157 VDDD.t5 VSSD 0.054937f
C3158 VDDD.t449 VSSD 0.056634f
C3159 VDDD.t252 VSSD 0.039029f
C3160 VDDD.t868 VSSD 0.020999f
C3161 VDDD.t727 VSSD 0.020999f
C3162 VDDD.t1194 VSSD 0.029696f
C3163 VDDD.t786 VSSD 0.029696f
C3164 VDDD.t599 VSSD 0.020575f
C3165 VDDD.t391 VSSD 0.020575f
C3166 VDDD.t325 VSSD 0.041786f
C3167 VDDD.t1875 VSSD 0.041786f
C3168 VDDD.t1435 VSSD 0.020999f
C3169 VDDD.t160 VSSD 0.019727f
C3170 VDDD.t91 VSSD 0.019514f
C3171 VDDD.t4 VSSD 0.017817f
C3172 VDDD.t1926 VSSD 0.018242f
C3173 VDDD.t597 VSSD 0.019514f
C3174 VDDD.t1231 VSSD 0.021211f
C3175 VDDD.t393 VSSD 0.021211f
C3176 VDDD.t559 VSSD 0.019514f
C3177 VDDD.t289 VSSD 0.019514f
C3178 VDDD.t1931 VSSD 0.043908f
C3179 VDDD.t201 VSSD 0.043908f
C3180 VDDD.t1263 VSSD 0.019514f
C3181 VDDD.t1233 VSSD 0.019514f
C3182 VDDD.t1235 VSSD 0.029696f
C3183 VDDD.n2740 VSSD 0.031241f
C3184 VDDD.n2741 VSSD 0.012205f
C3185 VDDD.n2743 VSSD 0.010729f
C3186 VDDD.n2744 VSSD 0.013262f
C3187 VDDD.n2745 VSSD 0.011542f
C3188 VDDD.n2757 VSSD 0.199537f
C3189 VDDD.n2787 VSSD 0.050066f
C3190 VDDD.n2791 VSSD 0.017188f
C3191 VDDD.n2792 VSSD 0.013558f
C3192 VDDD.n2813 VSSD 0.010232f
C3193 VDDD.n2819 VSSD 0.013718f
C3194 VDDD.n2825 VSSD 0.013224f
C3195 VDDD.n2859 VSSD 0.013413f
C3196 VDDD.n2860 VSSD 0.042685f
C3197 VDDD.t1296 VSSD 0.019514f
C3198 VDDD.t746 VSSD 0.017817f
C3199 VDDD.t225 VSSD 0.020999f
C3200 VDDD.t206 VSSD 0.048786f
C3201 VDDD.t1684 VSSD 0.037544f
C3202 VDDD.t59 VSSD 0.020575f
C3203 VDDD.t1237 VSSD 0.019514f
C3204 VDDD.t110 VSSD 0.027787f
C3205 VDDD.t1425 VSSD 0.034999f
C3206 VDDD.t864 VSSD 0.029696f
C3207 VDDD.t933 VSSD 0.020999f
C3208 VDDD.t1265 VSSD 0.020575f
C3209 VDDD.t333 VSSD 0.018242f
C3210 VDDD.t1291 VSSD 0.020787f
C3211 VDDD.t539 VSSD 0.038817f
C3212 VDDD.t1428 VSSD 0.022908f
C3213 VDDD.t263 VSSD 0.019727f
C3214 VDDD.t921 VSSD 0.01909f
C3215 VDDD.t227 VSSD 0.019514f
C3216 VDDD.t111 VSSD 0.036059f
C3217 VDDD.t694 VSSD 0.02609f
C3218 VDDD.t535 VSSD 0.022908f
C3219 VDDD.t273 VSSD 0.017817f
C3220 VDDD.t537 VSSD 0.017817f
C3221 VDDD.t1715 VSSD 0.054725f
C3222 VDDD.t67 VSSD 0.023333f
C3223 VDDD.t696 VSSD 0.052392f
C3224 VDDD.t481 VSSD 0.045604f
C3225 VDDD.t1168 VSSD 0.052392f
C3226 VDDD.t1644 VSSD 0.015909f
C3227 VDDD.t1144 VSSD 0.058543f
C3228 VDDD.t523 VSSD 0.052392f
C3229 VDDD.t1747 VSSD 0.060665f
C3230 VDDD.t69 VSSD 0.058968f
C3231 VDDD.t71 VSSD 0.039029f
C3232 VDDD.t1969 VSSD 0.039029f
C3233 VDDD.t101 VSSD 0.024393f
C3234 VDDD.t589 VSSD 0.024393f
C3235 VDDD.t261 VSSD 0.039029f
C3236 VDDD.t878 VSSD 0.022908f
C3237 VDDD.t1312 VSSD 0.017817f
C3238 VDDD.t299 VSSD 0.017817f
C3239 VDDD.t908 VSSD 0.019939f
C3240 VDDD.t710 VSSD 0.021211f
C3241 VDDD.t1971 VSSD 0.020787f
C3242 VDDD.t949 VSSD 0.01803f
C3243 VDDD.t381 VSSD 0.018242f
C3244 VDDD.t862 VSSD 0.039029f
C3245 VDDD.t406 VSSD 0.023757f
C3246 VDDD.t1680 VSSD 0.023333f
C3247 VDDD.t1426 VSSD 0.039029f
C3248 VDDD.t339 VSSD 0.029696f
C3249 VDDD.t358 VSSD 0.020575f
C3250 VDDD.t1542 VSSD 0.020999f
C3251 VDDD.t909 VSSD 0.029696f
C3252 VDDD.t863 VSSD 0.019514f
C3253 VDDD.t1421 VSSD 0.020999f
C3254 VDDD.t954 VSSD 0.039029f
C3255 VDDD.t830 VSSD 0.03712f
C3256 VDDD.t708 VSSD 0.035423f
C3257 VDDD.t904 VSSD 0.024393f
C3258 VDDD.t860 VSSD 0.02312f
C3259 VDDD.n2861 VSSD 0.02145f
C3260 VDDD.t2046 VSSD 0.032941f
C3261 VDDD.n2881 VSSD 0.016544f
C3262 VDDD.n2882 VSSD 0.013033f
C3263 VDDD.t2112 VSSD 0.023382f
C3264 VDDD.n2884 VSSD 0.033916f
C3265 VDDD.n2885 VSSD 0.044325f
C3266 VDDD.t2098 VSSD 0.011988f
C3267 VDDD.n2887 VSSD 0.030737f
C3268 VDDD.n2888 VSSD 0.016743f
C3269 VDDD.t2019 VSSD 0.011988f
C3270 VDDD.n2890 VSSD 0.030737f
C3271 VDDD.n2891 VSSD 0.016743f
C3272 VDDD.n2893 VSSD 0.014113f
C3273 VDDD.n2896 VSSD 0.012466f
C3274 VDDD.n2900 VSSD 0.017377f
C3275 VDDD.n2901 VSSD 0.03716f
C3276 VDDD.n2905 VSSD 0.011723f
C3277 VDDD.n2911 VSSD 0.011427f
C3278 VDDD.n2939 VSSD 0.018612f
C3279 VDDD.n2943 VSSD 0.019274f
C3280 VDDD.n2944 VSSD 0.013033f
C3281 VDDD.n2945 VSSD 0.044325f
C3282 VDDD.n2946 VSSD 0.013033f
C3283 VDDD.n2956 VSSD 0.012844f
C3284 VDDD.n2957 VSSD 0.055912f
C3285 VDDD.n2964 VSSD 0.199537f
C3286 VDDD.n2965 VSSD 0.19393f
C3287 VDDD.n2980 VSSD 0.012183f
C3288 VDDD.n2981 VSSD 0.012886f
C3289 VDDD.n2988 VSSD 0.012412f
C3290 VDDD.n2993 VSSD 0.010704f
C3291 VDDD.n3000 VSSD 0.015726f
C3292 VDDD.n3001 VSSD 0.014166f
C3293 VDDD.n3002 VSSD 0.010388f
C3294 VDDD.n3008 VSSD 0.010857f
C3295 VDDD.n3009 VSSD 0.013545f
C3296 VDDD.n3010 VSSD 0.013917f
C3297 VDDD.n3017 VSSD 0.19393f
C3298 VDDD.n3018 VSSD 0.138631f
C3299 VDDD.n3019 VSSD 0.509672f
C3300 VDDD.n3020 VSSD 0.957816f
C3301 VDDD.n3021 VSSD 0.138631f
C3302 VDDD.n3022 VSSD 0.221962f
C3303 VDDD.n3035 VSSD 0.01274f
C3304 VDDD.n3074 VSSD 0.221962f
C3305 VDDD.n3075 VSSD 0.171505f
C3306 VDDD.n3081 VSSD 0.013708f
C3307 VDDD.n3090 VSSD 0.013718f
C3308 VDDD.n3095 VSSD 0.013033f
C3309 VDDD.n3098 VSSD 0.017775f
C3310 VDDD.n3099 VSSD 0.042483f
C3311 VDDD.t1055 VSSD 0.028211f
C3312 VDDD.t1322 VSSD 0.032878f
C3313 VDDD.t1947 VSSD 0.036059f
C3314 VDDD.t323 VSSD 0.045604f
C3315 VDDD.t585 VSSD 0.022484f
C3316 VDDD.t1595 VSSD 0.027787f
C3317 VDDD.t1619 VSSD 0.022908f
C3318 VDDD.t1320 VSSD 0.017817f
C3319 VDDD.t873 VSSD 0.017817f
C3320 VDDD.t763 VSSD 0.024817f
C3321 VDDD.t1362 VSSD 0.039029f
C3322 VDDD.t1207 VSSD 0.020999f
C3323 VDDD.t1201 VSSD 0.017817f
C3324 VDDD.t1490 VSSD 0.040514f
C3325 VDDD.t871 VSSD 0.024181f
C3326 VDDD.t1255 VSSD 0.017817f
C3327 VDDD.t881 VSSD 0.020575f
C3328 VDDD.t329 VSSD 0.018242f
C3329 VDDD.t1962 VSSD 0.029696f
C3330 VDDD.t1361 VSSD 0.020999f
C3331 VDDD.t465 VSSD 0.020999f
C3332 VDDD.t1189 VSSD 0.034999f
C3333 VDDD.t1482 VSSD 0.026302f
C3334 VDDD.t644 VSSD 0.027363f
C3335 VDDD.t1205 VSSD 0.049847f
C3336 VDDD.t185 VSSD 0.029696f
C3337 VDDD.t1961 VSSD 0.017817f
C3338 VDDD.t782 VSSD 0.020999f
C3339 VDDD.t880 VSSD 0.013787f
C3340 VDDD.t1375 VSSD 0.065967f
C3341 VDDD.t1359 VSSD 0.074452f
C3342 VDDD.t1963 VSSD 0.031605f
C3343 VDDD.t1827 VSSD 0.052392f
C3344 VDDD.t1836 VSSD 0.050907f
C3345 VDDD.t1567 VSSD 0.039453f
C3346 VDDD.t1563 VSSD 0.062998f
C3347 VDDD.t438 VSSD 0.018242f
C3348 VDDD.t253 VSSD 0.040726f
C3349 VDDD.t1565 VSSD 0.030757f
C3350 VDDD.t1637 VSSD 0.017817f
C3351 VDDD.t327 VSSD 0.017817f
C3352 VDDD.t1650 VSSD 0.018242f
C3353 VDDD.t228 VSSD 0.017817f
C3354 VDDD.t1635 VSSD 0.020999f
C3355 VDDD.t1330 VSSD 0.017817f
C3356 VDDD.t1546 VSSD 0.02206f
C3357 VDDD.t1550 VSSD 0.035635f
C3358 VDDD.t1544 VSSD 0.019727f
C3359 VDDD.t730 VSSD 0.017817f
C3360 VDDD.t1548 VSSD 0.020575f
C3361 VDDD.t123 VSSD 0.017817f
C3362 VDDD.t1639 VSSD 0.029696f
C3363 VDDD.t1690 VSSD 0.017817f
C3364 VDDD.t209 VSSD 0.01909f
C3365 VDDD.t473 VSSD 0.019727f
C3366 VDDD.t328 VSSD 0.017817f
C3367 VDDD.t211 VSSD 0.019514f
C3368 VDDD.t1691 VSSD 0.051968f
C3369 VDDD.t65 VSSD 0.024393f
C3370 VDDD.t1150 VSSD 0.042847f
C3371 VDDD.n3100 VSSD 0.029119f
C3372 VDDD.n3101 VSSD 0.019479f
C3373 VDDD.n3145 VSSD 0.013783f
C3374 VDDD.n3152 VSSD 0.022728f
C3375 VDDD.n3154 VSSD 0.021263f
C3376 VDDD.t2024 VSSD 0.042585f
C3377 VDDD.n3156 VSSD 0.072669f
C3378 VDDD.n3164 VSSD 0.171505f
C3379 VDDD.n3169 VSSD 0.026093f
C3380 VDDD.n3170 VSSD 0.062257f
C3381 VDDD.t1848 VSSD 0.077846f
C3382 VDDD.t1812 VSSD 0.019514f
C3383 VDDD.t1577 VSSD 0.024393f
C3384 VDDD.t1906 VSSD 0.051968f
C3385 VDDD.t939 VSSD 0.013575f
C3386 VDDD.t721 VSSD 0.019514f
C3387 VDDD.t725 VSSD 0.017817f
C3388 VDDD.t1351 VSSD 0.020999f
C3389 VDDD.t1553 VSSD 0.017817f
C3390 VDDD.t717 VSSD 0.023545f
C3391 VDDD.t1403 VSSD 0.023969f
C3392 VDDD.t1656 VSSD 0.017817f
C3393 VDDD.t1353 VSSD 0.020575f
C3394 VDDD.t728 VSSD 0.017817f
C3395 VDDD.t1405 VSSD 0.026726f
C3396 VDDD.t719 VSSD 0.032878f
C3397 VDDD.t858 VSSD 0.017817f
C3398 VDDD.t723 VSSD 0.020999f
C3399 VDDD.t1552 VSSD 0.036484f
C3400 VDDD.t1560 VSSD 0.036059f
C3401 VDDD.t776 VSSD 0.020575f
C3402 VDDD.t287 VSSD 0.037968f
C3403 VDDD.t604 VSSD 0.063422f
C3404 VDDD.t774 VSSD 0.046029f
C3405 VDDD.t1124 VSSD 0.017817f
C3406 VDDD.t947 VSSD 0.048786f
C3407 VDDD.t505 VSSD 0.058543f
C3408 VDDD.t839 VSSD 0.033302f
C3409 VDDD.t372 VSSD 0.063422f
C3410 VDDD.t426 VSSD 0.063422f
C3411 VDDD.t1227 VSSD 0.032029f
C3412 VDDD.t1859 VSSD 0.022908f
C3413 VDDD.t419 VSSD 0.026514f
C3414 VDDD.t807 VSSD 0.036059f
C3415 VDDD.t700 VSSD 0.039241f
C3416 VDDD.t369 VSSD 0.062786f
C3417 VDDD.t1251 VSSD 0.057483f
C3418 VDDD.t269 VSSD 0.034575f
C3419 VDDD.t847 VSSD 0.050695f
C3420 VDDD.t877 VSSD 0.040514f
C3421 VDDD.t919 VSSD 0.055362f
C3422 VDDD.t1822 VSSD 0.056634f
C3423 VDDD.t698 VSSD 0.038605f
C3424 VDDD.t1967 VSSD 0.024393f
C3425 VDDD.t971 VSSD 0.058543f
C3426 VDDD.n3171 VSSD 0.057967f
C3427 VDDD.n3173 VSSD 0.018356f
C3428 VDDD.t2111 VSSD 0.081647f
C3429 VDDD.t1982 VSSD 0.081647f
C3430 VDDD.n3181 VSSD 0.038136f
C3431 VDDD.n3187 VSSD 0.013211f
C3432 VDDD.t2035 VSSD 0.011988f
C3433 VDDD.n3189 VSSD 0.030737f
C3434 VDDD.n3190 VSSD 0.016743f
C3435 VDDD.t2000 VSSD 0.011988f
C3436 VDDD.n3192 VSSD 0.030737f
C3437 VDDD.n3193 VSSD 0.016743f
C3438 VDDD.n3195 VSSD 0.014123f
C3439 VDDD.n3200 VSSD 0.014872f
C3440 VDDD.n3236 VSSD 0.038045f
C3441 VDDD.n3240 VSSD 0.014405f
C3442 VDDD.n3241 VSSD 0.04001f
C3443 VDDD.t2075 VSSD 0.023828f
C3444 VDDD.n3248 VSSD 0.032397f
C3445 VDDD.n3250 VSSD 0.01711f
C3446 VDDD.n3251 VSSD 0.016338f
C3447 VDDD.n3255 VSSD 0.011994f
C3448 VDDD.n3257 VSSD 0.052607f
C3449 VDDD.n3258 VSSD 0.012655f
C3450 VDDD.n3276 VSSD 0.171505f
C3451 VDDD.n3277 VSSD 0.138631f
C3452 VDDD.n3278 VSSD 0.676845f
C3453 VDDD.n3279 VSSD 0.509672f
C3454 VDDD.n3280 VSSD 0.957816f
C3455 VDDD.n3281 VSSD 0.138631f
C3456 VDDD.n3282 VSSD 0.244388f
C3457 VDDD.n3288 VSSD 0.010913f
C3458 VDDD.n3291 VSSD 0.012787f
C3459 VDDD.n3292 VSSD 0.019574f
C3460 VDDD.t656 VSSD 0.020787f
C3461 VDDD.t950 VSSD 0.038817f
C3462 VDDD.t517 VSSD 0.029696f
C3463 VDDD.t187 VSSD 0.02312f
C3464 VDDD.t178 VSSD 0.028848f
C3465 VDDD.t691 VSSD 0.074876f
C3466 VDDD.t1036 VSSD 0.056634f
C3467 VDDD.t140 VSSD 0.01909f
C3468 VDDD.t891 VSSD 0.031605f
C3469 VDDD.t976 VSSD 0.039029f
C3470 VDDD.t37 VSSD 0.025029f
C3471 VDDD.t21 VSSD 0.036484f
C3472 VDDD.t1247 VSSD 0.036484f
C3473 VDDD.t23 VSSD 0.036484f
C3474 VDDD.t459 VSSD 0.022696f
C3475 VDDD.t1096 VSSD 0.018242f
C3476 VDDD.t125 VSSD 0.032029f
C3477 VDDD.t1601 VSSD 0.036484f
C3478 VDDD.t1597 VSSD 0.036484f
C3479 VDDD.t127 VSSD 0.021636f
C3480 VDDD.t1180 VSSD 0.019514f
C3481 VDDD.t129 VSSD 0.015272f
C3482 VDDD.t75 VSSD 0.018242f
C3483 VDDD.t819 VSSD 0.034575f
C3484 VDDD.t131 VSSD 0.036271f
C3485 VDDD.t461 VSSD 0.034362f
C3486 VDDD.t1761 VSSD 0.018242f
C3487 VDDD.t457 VSSD 0.020363f
C3488 VDDD.t821 VSSD 0.030757f
C3489 VDDD.t1599 VSSD 0.015909f
C3490 VDDD.n3293 VSSD 0.021898f
C3491 VDDD.t2021 VSSD 0.011582f
C3492 VDDD.n3298 VSSD 0.010572f
C3493 VDDD.n3299 VSSD 0.012734f
C3494 VDDD.n3301 VSSD 0.014424f
C3495 VDDD.t2055 VSSD 0.042035f
C3496 VDDD.n3302 VSSD 0.070387f
C3497 VDDD.n3303 VSSD 0.018492f
C3498 VDDD.t2071 VSSD 0.032941f
C3499 VDDD.n3324 VSSD 0.011268f
C3500 VDDD.n3326 VSSD 0.01711f
C3501 VDDD.n3344 VSSD 0.014424f
C3502 VDDD.n3345 VSSD 0.021661f
C3503 VDDD.t1990 VSSD 0.042035f
C3504 VDDD.n3347 VSSD 0.070387f
C3505 VDDD.n3348 VSSD 0.026923f
C3506 VDDD.n3349 VSSD 0.039466f
C3507 VDDD.t2085 VSSD 0.023588f
C3508 VDDD.n3351 VSSD 0.04098f
C3509 VDDD.n3352 VSSD 0.023515f
C3510 VDDD.t2037 VSSD 0.011988f
C3511 VDDD.n3354 VSSD 0.030737f
C3512 VDDD.n3355 VSSD 0.016743f
C3513 VDDD.t1995 VSSD 0.011988f
C3514 VDDD.n3357 VSSD 0.030737f
C3515 VDDD.n3358 VSSD 0.016743f
C3516 VDDD.n3360 VSSD 0.013785f
C3517 VDDD.n3361 VSSD 0.02207f
C3518 VDDD.n3364 VSSD 0.013386f
C3519 VDDD.t133 VSSD 0.026302f
C3520 VDDD.t1178 VSSD 0.030969f
C3521 VDDD.t1784 VSSD 0.018242f
C3522 VDDD.t455 VSSD 0.02312f
C3523 VDDD.t529 VSSD 0.024393f
C3524 VDDD.t1274 VSSD 0.074452f
C3525 VDDD.t1617 VSSD 0.059816f
C3526 VDDD.t1000 VSSD 0.019514f
C3527 VDDD.t418 VSSD 0.037332f
C3528 VDDD.t1229 VSSD 0.050695f
C3529 VDDD.t848 VSSD 0.034575f
C3530 VDDD.t1488 VSSD 0.019514f
C3531 VDDD.t1613 VSSD 0.024817f
C3532 VDDD.t1615 VSSD 0.030969f
C3533 VDDD.t845 VSSD 0.03415f
C3534 VDDD.t1273 VSSD 0.029272f
C3535 VDDD.t815 VSSD 0.018242f
C3536 VDDD.t528 VSSD 0.017817f
C3537 VDDD.t1708 VSSD 0.017817f
C3538 VDDD.t1713 VSSD 0.017817f
C3539 VDDD.t1710 VSSD 0.022908f
C3540 VDDD.t1472 VSSD 0.017817f
C3541 VDDD.t813 VSSD 0.017817f
C3542 VDDD.t619 VSSD 0.015909f
C3543 VDDD.t117 VSSD 0.043483f
C3544 VDDD.t115 VSSD 0.039453f
C3545 VDDD.t1006 VSSD 0.043271f
C3546 VDDD.t250 VSSD 0.039453f
C3547 VDDD.t175 VSSD 0.030757f
C3548 VDDD.t511 VSSD 0.058543f
C3549 VDDD.t1021 VSSD 0.071906f
C3550 VDDD.t1044 VSSD 0.060665f
C3551 VDDD.t1215 VSSD 0.039453f
C3552 VDDD.t1219 VSSD 0.062573f
C3553 VDDD.t1357 VSSD 0.013787f
C3554 VDDD.t531 VSSD 0.017817f
C3555 VDDD.t1587 VSSD 0.017817f
C3556 VDDD.t545 VSSD 0.022908f
C3557 VDDD.t1217 VSSD 0.027787f
C3558 VDDD.t1533 VSSD 0.036059f
C3559 VDDD.t1621 VSSD 0.028848f
C3560 VDDD.t1461 VSSD 0.020999f
C3561 VDDD.t744 VSSD 0.019514f
C3562 VDDD.t960 VSSD 0.03012f
C3563 VDDD.t1099 VSSD 0.032666f
C3564 VDDD.t1398 VSSD 0.029696f
C3565 VDDD.t1271 VSSD 0.020575f
C3566 VDDD.t747 VSSD 0.020575f
C3567 VDDD.t1257 VSSD 0.029696f
C3568 VDDD.t1622 VSSD 0.032666f
C3569 VDDD.t1532 VSSD 0.03012f
C3570 VDDD.t841 VSSD 0.019514f
C3571 VDDD.t686 VSSD 0.020999f
C3572 VDDD.t1100 VSSD 0.028848f
C3573 VDDD.t606 VSSD 0.036059f
C3574 VDDD.t248 VSSD 0.027787f
C3575 VDDD.t680 VSSD 0.022908f
C3576 VDDD.t1492 VSSD 0.017817f
C3577 VDDD.t137 VSSD 0.011454f
C3578 VDDD.t84 VSSD 0.02312f
C3579 VDDD.n3397 VSSD 0.036119f
C3580 VDDD.n3398 VSSD 0.012591f
C3581 VDDD.n3400 VSSD 0.011268f
C3582 VDDD.n3402 VSSD 0.016244f
C3583 VDDD.n3407 VSSD 0.01711f
C3584 VDDD.n3408 VSSD 0.044149f
C3585 VDDD.n3420 VSSD 0.010781f
C3586 VDDD.n3439 VSSD 0.01681f
C3587 VDDD.n3440 VSSD 0.017377f
C3588 VDDD.n3441 VSSD 0.01426f
C3589 VDDD.n3442 VSSD 0.013193f
C3590 VDDD.n3443 VSSD 0.011265f
C3591 VDDD.n3446 VSSD 0.015556f
C3592 VDDD.n3448 VSSD 0.014253f
C3593 VDDD.n3449 VSSD 0.010414f
C3594 VDDD.n3462 VSSD 0.011693f
C3595 VDDD.n3464 VSSD 0.010723f
C3596 VDDD.n3471 VSSD 0.244388f
C3597 VDDD.n3482 VSSD 0.013708f
C3598 VDDD.n3495 VSSD 0.013708f
C3599 VDDD.n3504 VSSD 0.012594f
C3600 VDDD.n3508 VSSD 0.014873f
C3601 VDDD.n3574 VSSD 0.149079f
C3602 VDDD.n3612 VSSD 0.012922f
C3603 VDDD.n3613 VSSD 0.03791f
C3604 VDDD.n3614 VSSD 0.012594f
C3605 VDDD.n3624 VSSD 0.149079f
C3606 VDDD.n3631 VSSD 0.012594f
C3607 VDDD.n3644 VSSD 0.013537f
C3608 VDDD.t1063 VSSD 0.058543f
C3609 VDDD.t496 VSSD 0.071906f
C3610 VDDD.t1793 VSSD 0.04518f
C3611 VDDD.t761 VSSD 0.031605f
C3612 VDDD.t689 VSSD 0.06427f
C3613 VDDD.t587 VSSD 0.02312f
C3614 VDDD.t502 VSSD 0.019514f
C3615 VDDD.t1942 VSSD 0.027575f
C3616 VDDD.t581 VSSD 0.028848f
C3617 VDDD.t889 VSSD 0.021848f
C3618 VDDD.t343 VSSD 0.017817f
C3619 VDDD.t1283 VSSD 0.020575f
C3620 VDDD.t1589 VSSD 0.052604f
C3621 VDDD.t203 VSSD 0.045817f
C3622 VDDD.t1176 VSSD 0.020999f
C3623 VDDD.t688 VSSD 0.019514f
C3624 VDDD.t2 VSSD 0.018242f
C3625 VDDD.t827 VSSD 0.020999f
C3626 VDDD.t1282 VSSD 0.017817f
C3627 VDDD.t791 VSSD 0.029696f
C3628 VDDD.t467 VSSD 0.022908f
C3629 VDDD.t215 VSSD 0.020575f
C3630 VDDD.t1474 VSSD 0.017817f
C3631 VDDD.t937 VSSD 0.041786f
C3632 VDDD.t1285 VSSD 0.045604f
C3633 VDDD.t789 VSSD 0.020999f
C3634 VDDD.t834 VSSD 0.017817f
C3635 VDDD.t793 VSSD 0.018242f
C3636 VDDD.t3 VSSD 0.031393f
C3637 VDDD.n3645 VSSD 0.021474f
C3638 VDDD.t165 VSSD 0.015909f
C3639 VDDD.t1470 VSSD 0.025878f
C3640 VDDD.t471 VSSD 0.063422f
C3641 VDDD.t896 VSSD 0.063422f
C3642 VDDD.t898 VSSD 0.039453f
C3643 VDDD.t493 VSSD 0.043271f
C3644 VDDD.t935 VSSD 0.039453f
C3645 VDDD.t1336 VSSD 0.063422f
C3646 VDDD.t96 VSSD 0.063422f
C3647 VDDD.t1581 VSSD 0.038605f
C3648 VDDD.t1334 VSSD 0.01909f
C3649 VDDD.t584 VSSD 0.013787f
C3650 VDDD.t533 VSSD 0.018242f
C3651 VDDD.t1371 VSSD 0.017817f
C3652 VDDD.t1973 VSSD 0.020999f
C3653 VDDD.t1440 VSSD 0.050271f
C3654 VDDD.t658 VSSD 0.04815f
C3655 VDDD.t1922 VSSD 0.020575f
C3656 VDDD.t156 VSSD 0.019514f
C3657 VDDD.t87 VSSD 0.026302f
C3658 VDDD.t824 VSSD 0.024393f
C3659 VDDD.t1372 VSSD 0.024393f
C3660 VDDD.t88 VSSD 0.026302f
C3661 VDDD.t15 VSSD 0.019514f
C3662 VDDD.t1693 VSSD 0.020575f
C3663 VDDD.t1480 VSSD 0.04815f
C3664 VDDD.t526 VSSD 0.050271f
C3665 VDDD.t1369 VSSD 0.020999f
C3666 VDDD.t823 VSSD 0.017817f
C3667 VDDD.t952 VSSD 0.011878f
C3668 VDDD.t86 VSSD 0.02312f
C3669 VDDD.n3646 VSSD 0.021474f
C3670 VDDD.t869 VSSD 0.016333f
C3671 VDDD.t640 VSSD 0.01909f
C3672 VDDD.t850 VSSD 0.013787f
C3673 VDDD.t887 VSSD 0.025242f
C3674 VDDD.t1300 VSSD 0.038181f
C3675 VDDD.t609 VSSD 0.038181f
C3676 VDDD.t607 VSSD 0.036271f
C3677 VDDD.t92 VSSD 0.027787f
C3678 VDDD.t1367 VSSD 0.013787f
C3679 VDDD.t759 VSSD 0.020999f
C3680 VDDD.t677 VSSD 0.017817f
C3681 VDDD.t1437 VSSD 0.029696f
C3682 VDDD.t1510 VSSD 0.049847f
C3683 VDDD.t674 VSSD 0.027363f
C3684 VDDD.t173 VSSD 0.026302f
C3685 VDDD.t886 VSSD 0.034999f
C3686 VDDD.t403 VSSD 0.020999f
C3687 VDDD.t1905 VSSD 0.020999f
C3688 VDDD.t676 VSSD 0.029696f
C3689 VDDD.t1937 VSSD 0.018242f
C3690 VDDD.t1874 VSSD 0.020575f
C3691 VDDD.t1585 VSSD 0.017817f
C3692 VDDD.t1918 VSSD 0.024181f
C3693 VDDD.t1486 VSSD 0.040514f
C3694 VDDD.t239 VSSD 0.017817f
C3695 VDDD.t1702 VSSD 0.020999f
C3696 VDDD.t1439 VSSD 0.039029f
C3697 VDDD.t885 VSSD 0.024817f
C3698 VDDD.t1920 VSSD 0.017817f
C3699 VDDD.t1444 VSSD 0.017817f
C3700 VDDD.t969 VSSD 0.022908f
C3701 VDDD.t1583 VSSD 0.027787f
C3702 VDDD.t633 VSSD 0.051968f
C3703 VDDD.t961 VSSD 0.063422f
C3704 VDDD.t45 VSSD 0.04921f
C3705 VDDD.n3647 VSSD 0.044604f
C3706 VDDD.n3648 VSSD 0.019479f
C3707 VDDD.n3675 VSSD 0.038136f
C3708 VDDD.n3688 VSSD 0.149079f
C3709 VDDD.n3689 VSSD 0.33981f
C3710 VDDD.n3690 VSSD 0.676845f
C3711 VDDD.n3691 VSSD 0.509672f
C3712 VDDD.n3692 VSSD 0.957816f
C3713 VDDD.n3693 VSSD 0.138631f
C3714 VDDD.n3694 VSSD 0.140415f
C3715 VDDD.n3702 VSSD 0.014638f
C3716 VDDD.n3706 VSSD 0.013942f
C3717 VDDD.n3707 VSSD 0.034813f
C3718 VDDD.t1159 VSSD 0.035247f
C3719 VDDD.t1833 VSSD 0.132808f
C3720 VDDD.t1115 VSSD 0.132808f
C3721 VDDD.t1156 VSSD 0.033201f
C3722 VDDD.t1781 VSSD 0.132808f
C3723 VDDD.t478 VSSD 0.133048f
C3724 VDDD.n3708 VSSD 0.02579f
C3725 VDDD.t893 VSSD 0.017924f
C3726 VDDD.t98 VSSD 0.042224f
C3727 VDDD.t1877 VSSD 0.043187f
C3728 VDDD.t637 VSSD 0.022976f
C3729 VDDD.t100 VSSD 0.028751f
C3730 VDDD.t1623 VSSD 0.02851f
C3731 VDDD.t638 VSSD 0.035367f
C3732 VDDD.t1611 VSSD 0.035607f
C3733 VDDD.t1346 VSSD 0.022255f
C3734 VDDD.t1525 VSSD 0.020451f
C3735 VDDD.t171 VSSD 0.023097f
C3736 VDDD.t1396 VSSD 0.023097f
C3737 VDDD.t1515 VSSD 0.035969f
C3738 VDDD.t711 VSSD 0.035969f
C3739 VDDD.t169 VSSD 0.025864f
C3740 VDDD.t1130 VSSD 0.044509f
C3741 VDDD.n3709 VSSD 0.02555f
C3742 VDDD.n3715 VSSD 0.013984f
C3743 VDDD.n3722 VSSD 0.140415f
C3744 VDDD.n3730 VSSD 0.021149f
C3745 VDDD.n3731 VSSD 0.013033f
C3746 VDDD.n3732 VSSD 0.01681f
C3747 VDDD.n3736 VSSD 0.011152f
C3748 VDDD.n3764 VSSD 0.140415f
C3749 VDDD.n3829 VSSD 0.017816f
C3750 VDDD.n3830 VSSD 0.014638f
C3751 VDDD.n3831 VSSD 0.015255f
.ends

