* NGSPICE file created from all.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_lvt_A33RKA w_n231_n261# a_35_n42# a_n35_n139# a_n93_n42#
X0 a_35_n42# a_n35_n139# a_n93_n42# w_n231_n261# sky130_fd_pr__pfet_01v8_lvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.35
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_BK97Z7 a_n33_n130# a_15_n42# a_n175_n216# a_n73_n42#
X0 a_15_n42# a_n33_n130# a_n73_n42# a_n175_n216# sky130_fd_pr__nfet_01v8_lvt ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
.ends

.subckt epc_delay VSS IN OUT VIN VDD
XXM1 VDD li_225_237# VIN VDD sky130_fd_pr__pfet_01v8_lvt_A33RKA
XXM2 VDD OUT IN li_225_237# sky130_fd_pr__pfet_01v8_lvt_A33RKA
XXM3 IN OUT VSS li_266_n350# sky130_fd_pr__nfet_01v8_lvt_BK97Z7
XXM4 VIN li_266_n350# VSS VSS sky130_fd_pr__nfet_01v8_lvt_BK97Z7
.ends

.subckt epc_delay_line VDD IN VSS OUT VP VN
Xx1 VSS IN x2/IN VP VDD epc_delay
Xx2 VSS x2/IN x3/IN VN VDD epc_delay
Xx3 VSS x3/IN x4/IN VP VDD epc_delay
Xx4 VSS x4/IN x5/IN VN VDD epc_delay
Xx5 VSS x5/IN x6/IN VP VDD epc_delay
Xx6 VSS x6/IN x7/IN VN VDD epc_delay
Xx7 VSS x7/IN x8/IN VP VDD epc_delay
Xx8 VSS x8/IN OUT VN VDD epc_delay
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt all VDDA OUTN VSSA VP VN OUTP
Xx1 VDDA x1/IN VSSA x1/OUT VP VN epc_delay_line
Xx2 VDDA x2/IN VSSA x2/OUT VP VN epc_delay_line
Xx9 x9/A x9/B VSSA VSSA VDDA VDDA x9/Y sky130_fd_sc_hd__nand2_1
Xx10 x10/A x10/B VSSA VSSA VDDA VDDA x10/Y sky130_fd_sc_hd__nand2_1
.ends

