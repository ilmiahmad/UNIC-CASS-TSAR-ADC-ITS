magic
tech sky130A
magscale 1 2
timestamp 1730626724
<< nwell >>
rect -562 89 7 92
rect 13 89 2734 92
rect -562 -473 2734 89
<< pwell >>
rect -562 150 2734 360
rect -562 -742 2734 -532
<< psubdiff >>
rect -562 360 -495 394
rect 2667 360 2734 394
rect -562 -776 -495 -742
rect 2667 -776 2734 -742
<< nsubdiff >>
rect -471 -143 -447 56
rect -295 -143 -271 56
rect 284 32 318 56
rect 284 -438 318 -414
<< psubdiffcont >>
rect -495 360 2667 394
rect -495 -776 2667 -742
<< nsubdiffcont >>
rect -447 -143 -295 56
rect 284 -414 318 32
<< locali >>
rect -524 360 -495 394
rect 2667 360 2696 394
rect -471 -143 -447 56
rect -295 -143 -271 56
rect -471 -174 -271 -143
rect 284 32 318 56
rect 284 -438 318 -414
rect -524 -776 -495 -742
rect 2667 -776 2696 -742
<< viali >>
rect -128 234 -94 268
rect -220 98 -186 132
rect -36 98 -2 132
rect 100 98 134 132
rect 192 98 226 132
rect 376 98 410 132
rect 468 98 502 132
rect 609 98 643 132
rect 701 98 735 132
rect 793 98 827 132
rect 885 98 919 132
rect 977 98 1011 132
rect 1253 98 1287 132
rect 1345 98 1379 132
rect 1437 98 1471 132
rect 1529 98 1563 132
rect 1621 98 1655 132
rect 1713 98 1747 132
rect 1805 98 1839 132
rect 2081 98 2115 132
rect 2173 98 2207 132
rect 2265 98 2299 132
rect 2357 98 2391 132
rect 2449 98 2483 132
rect 2541 98 2575 132
rect 2633 98 2667 132
rect -452 -514 -418 -480
rect -360 -514 -326 -480
rect -220 -514 -186 -480
rect -36 -514 -2 -480
rect 100 -514 134 -480
rect 192 -514 226 -480
rect 376 -514 410 -480
rect 468 -514 502 -480
rect 609 -514 643 -480
rect 701 -514 735 -480
rect 793 -514 827 -480
rect 885 -514 919 -480
rect 977 -514 1011 -480
rect 1253 -514 1287 -480
rect 1345 -514 1379 -480
rect 1437 -514 1471 -480
rect 1529 -514 1563 -480
rect 1621 -514 1655 -480
rect 1713 -514 1747 -480
rect 1805 -514 1839 -480
rect 2081 -514 2115 -480
rect 2173 -514 2207 -480
rect 2265 -514 2299 -480
rect 2357 -514 2391 -480
rect 2449 -514 2483 -480
rect 2541 -514 2575 -480
rect 2633 -514 2667 -480
rect -128 -650 -94 -616
<< metal1 >>
rect -524 395 -248 401
rect -524 305 -255 395
rect -140 268 143 277
rect -140 234 -128 268
rect -94 234 143 268
rect -140 225 143 234
rect -229 132 -177 144
rect -229 98 -220 132
rect -186 98 -177 132
rect -229 58 -177 98
rect -117 89 -111 141
rect -59 132 10 141
rect -59 98 -36 132
rect -2 98 10 132
rect -59 89 10 98
rect 91 132 143 225
rect 568 169 574 221
rect 626 169 2676 221
rect 91 98 100 132
rect 134 98 143 132
rect 91 86 143 98
rect 180 132 422 141
rect 180 98 192 132
rect 226 98 376 132
rect 410 98 422 132
rect 180 89 422 98
rect 453 89 459 141
rect 511 132 931 141
rect 511 98 609 132
rect 643 98 701 132
rect 735 98 793 132
rect 827 98 885 132
rect 919 98 931 132
rect 511 89 931 98
rect 965 132 1759 141
rect 965 98 977 132
rect 1011 98 1253 132
rect 1287 98 1345 132
rect 1379 98 1437 132
rect 1471 98 1529 132
rect 1563 98 1621 132
rect 1655 98 1713 132
rect 1747 98 1759 132
rect 965 89 1759 98
rect 1793 132 2587 141
rect 1793 98 1805 132
rect 1839 98 2081 132
rect 2115 98 2173 132
rect 2207 98 2265 132
rect 2299 98 2357 132
rect 2391 98 2449 132
rect 2483 98 2541 132
rect 2575 98 2587 132
rect 1793 89 2587 98
rect 2624 132 2676 169
rect 2624 98 2633 132
rect 2667 98 2676 132
rect -229 6 543 58
rect 595 6 601 58
rect 1793 -22 1845 89
rect 2624 85 2676 98
rect -467 -74 -461 -22
rect -409 -74 -111 -22
rect -59 -74 -53 -22
rect 76 -74 82 -22
rect 134 -74 1845 -22
rect -45 -440 459 -388
rect 511 -440 517 -388
rect 1446 -440 1452 -388
rect 1504 -440 1845 -388
rect 1938 -440 1944 -388
rect 1996 -440 2676 -388
rect -467 -523 -461 -471
rect -409 -523 -403 -471
rect -372 -480 -174 -471
rect -372 -514 -360 -480
rect -326 -514 -220 -480
rect -186 -514 -174 -480
rect -372 -523 -174 -514
rect -45 -480 7 -440
rect -45 -514 -36 -480
rect -2 -514 7 -480
rect -45 -526 7 -514
rect 91 -480 143 -468
rect 1793 -471 1845 -440
rect 91 -514 100 -480
rect 134 -514 143 -480
rect 91 -607 143 -514
rect 180 -480 422 -471
rect 180 -514 192 -480
rect 226 -514 376 -480
rect 410 -514 422 -480
rect 180 -523 422 -514
rect 456 -480 543 -471
rect 456 -514 468 -480
rect 502 -514 543 -480
rect 456 -523 543 -514
rect 595 -480 931 -471
rect 595 -514 609 -480
rect 643 -514 701 -480
rect 735 -514 793 -480
rect 827 -514 885 -480
rect 919 -514 931 -480
rect 595 -523 931 -514
rect 965 -480 1759 -471
rect 965 -514 977 -480
rect 1011 -514 1253 -480
rect 1287 -514 1345 -480
rect 1379 -514 1437 -480
rect 1471 -514 1529 -480
rect 1563 -514 1621 -480
rect 1655 -514 1713 -480
rect 1747 -514 1759 -480
rect 965 -523 1759 -514
rect 1793 -480 2587 -471
rect 1793 -514 1805 -480
rect 1839 -514 2081 -480
rect 2115 -514 2173 -480
rect 2207 -514 2265 -480
rect 2299 -514 2357 -480
rect 2391 -514 2449 -480
rect 2483 -514 2541 -480
rect 2575 -514 2587 -480
rect 1793 -523 2587 -514
rect 2624 -480 2676 -440
rect 2624 -514 2633 -480
rect 2667 -514 2676 -480
rect 2624 -526 2676 -514
rect -140 -616 143 -607
rect -140 -650 -128 -616
rect -94 -650 143 -616
rect -140 -659 143 -650
<< via1 >>
rect -255 305 -159 395
rect -111 89 -59 141
rect 574 169 626 221
rect 459 132 511 141
rect 459 98 468 132
rect 468 98 502 132
rect 502 98 511 132
rect 459 89 511 98
rect 543 6 595 58
rect -461 -74 -409 -22
rect -111 -74 -59 -22
rect 82 -74 134 -22
rect 182 -233 278 -143
rect 459 -440 511 -388
rect 1452 -440 1504 -388
rect 1944 -440 1996 -388
rect -461 -480 -409 -471
rect -461 -514 -452 -480
rect -452 -514 -418 -480
rect -418 -514 -409 -480
rect -461 -523 -409 -514
rect 543 -523 595 -471
rect -255 -777 -159 -687
<< metal2 >>
rect -255 395 -159 401
rect -463 -22 -407 -16
rect -463 -74 -461 -22
rect -409 -74 -407 -22
rect -463 -471 -407 -74
rect -463 -523 -461 -471
rect -409 -523 -407 -471
rect -463 -529 -407 -523
rect -255 -687 -159 305
rect -113 141 -57 401
rect -113 89 -111 141
rect -59 89 -57 141
rect -113 -22 -57 89
rect -113 -74 -111 -22
rect -59 -74 -57 -22
rect -113 -80 -57 -74
rect 80 -22 136 401
rect 80 -74 82 -22
rect 134 -74 136 -22
rect 80 -80 136 -74
rect 182 -143 278 401
rect 572 221 628 401
rect 572 169 574 221
rect 626 169 628 221
rect 572 163 628 169
rect 182 -239 278 -233
rect 457 141 513 147
rect 457 89 459 141
rect 511 89 513 141
rect 457 -388 513 89
rect 457 -440 459 -388
rect 511 -440 513 -388
rect 457 -446 513 -440
rect 541 58 597 64
rect 541 6 543 58
rect 595 6 597 58
rect 541 -471 597 6
rect 1450 -388 1506 401
rect 1450 -440 1452 -388
rect 1504 -440 1506 -388
rect 1450 -446 1506 -440
rect 1942 -388 1998 401
rect 1942 -440 1944 -388
rect 1996 -440 1998 -388
rect 1942 -446 1998 -440
rect 541 -523 543 -471
rect 595 -523 597 -471
rect 541 -529 597 -523
rect -255 -783 -159 -777
use sky130_fd_sc_hd__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1720120574
transform 1 0 -248 0 -1 353
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1720120574
transform 1 0 -248 0 1 -735
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1720120574
transform 1 0 -524 0 1 -735
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x4
timestamp 1720120574
transform 1 0 28 0 -1 353
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1720120574
transform 1 0 28 0 1 -735
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1720120574
transform 1 0 304 0 -1 353
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1720120574
transform 1 0 304 0 1 -735
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1720120574
transform 1 0 580 0 -1 353
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  x9
timestamp 1720120574
transform 1 0 580 0 1 -735
box -38 -48 498 592
use sky130_fd_sc_hd__inv_8  x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1720120574
transform 1 0 1040 0 -1 353
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x11
timestamp 1720120574
transform 1 0 1040 0 1 -735
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x12
timestamp 1720120574
transform 1 0 1868 0 -1 353
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x13
timestamp 1720120574
transform 1 0 1868 0 1 -735
box -38 -48 866 592
<< labels >>
flabel metal2 -113 345 -57 401 0 FreeSans 320 0 0 0 in
port 2 nsew
flabel metal2 80 345 136 401 0 FreeSans 320 0 0 0 clkb0
port 5 nsew
flabel metal2 572 345 628 401 0 FreeSans 320 0 0 0 clk0
port 4 nsew
flabel metal2 1450 345 1506 401 0 FreeSans 320 0 0 0 clkb1
port 7 nsew
flabel metal2 1942 345 1998 401 0 FreeSans 320 0 0 0 clk1
port 6 nsew
flabel metal2 -255 305 -159 401 0 FreeSans 320 0 0 0 vssa
port 3 nsew
flabel metal2 182 305 278 401 0 FreeSans 320 0 0 0 vdda
port 1 nsew
<< end >>
