magic
tech sky130A
magscale 1 2
timestamp 1730783553
<< nwell >>
rect 9948 -18 9980 114
rect 10032 -16 10064 112
rect 10295 26 10521 161
rect 10294 0 10521 26
rect 10295 -65 10521 0
<< pwell >>
rect 176 388 10468 572
rect 176 -476 10468 -292
<< psubdiff >>
rect 10348 548 10468 572
rect 10348 404 10468 428
rect 10348 -332 10468 -308
rect 10348 -476 10468 -452
<< nsubdiff >>
rect 10331 91 10391 125
rect 10425 91 10485 125
rect 10331 65 10365 91
rect 10331 5 10365 31
rect 10451 65 10485 91
rect 10451 5 10485 31
rect 10331 -29 10391 5
rect 10425 -29 10485 5
<< psubdiffcont >>
rect 10348 428 10468 548
rect 10348 -452 10468 -332
<< nsubdiffcont >>
rect 10391 91 10425 125
rect 10331 31 10365 65
rect 10451 31 10485 65
rect 10391 -29 10425 5
<< locali >>
rect 10348 548 10468 564
rect 10348 412 10468 428
rect 10331 91 10391 125
rect 10425 91 10485 125
rect 10331 65 10365 91
rect 10331 5 10365 31
rect 10451 65 10485 91
rect 10451 5 10485 31
rect 10331 -29 10391 5
rect 10425 -29 10485 5
rect 10348 -332 10468 -316
rect 10348 -468 10468 -452
<< viali >>
rect 10348 428 10468 548
rect 10046 334 10086 374
rect 10228 256 10268 296
rect 9856 166 9896 236
rect 10331 31 10365 65
rect 10451 31 10485 65
rect 9856 -140 9896 -70
rect 10228 -200 10268 -160
rect 10046 -276 10086 -236
rect 10348 -452 10468 -332
<< metal1 >>
rect -66 544 178 640
rect 10294 548 10574 640
rect 10294 544 10348 548
rect 10336 428 10348 544
rect 10468 428 10480 548
rect 10336 422 10480 428
rect 10030 328 10040 380
rect 10092 328 10102 380
rect 10212 250 10222 302
rect 10274 250 10284 302
rect 9850 236 9902 248
rect 9840 166 9850 236
rect 9902 166 9912 236
rect 9850 154 9902 166
rect -66 0 178 96
rect 10294 65 10504 96
rect 10294 31 10331 65
rect 10365 31 10451 65
rect 10485 31 10504 65
rect 10294 0 10504 31
rect 9850 -70 9902 -58
rect 9840 -140 9850 -70
rect 9902 -140 9912 -70
rect 9850 -152 9902 -140
rect 10212 -206 10222 -154
rect 10274 -206 10284 -154
rect 10030 -282 10040 -230
rect 10092 -282 10102 -230
rect 10336 -332 10480 -326
rect 10336 -448 10348 -332
rect -66 -544 178 -448
rect 10294 -452 10348 -448
rect 10468 -452 10480 -332
rect 10294 -544 10574 -452
<< via1 >>
rect 10040 374 10092 380
rect 10040 334 10046 374
rect 10046 334 10086 374
rect 10086 334 10092 374
rect 10040 328 10092 334
rect 10222 296 10274 302
rect 10222 256 10228 296
rect 10228 256 10268 296
rect 10268 256 10274 296
rect 10222 250 10274 256
rect 9850 166 9856 236
rect 9856 166 9896 236
rect 9896 166 9902 236
rect 9850 -140 9856 -70
rect 9856 -140 9896 -70
rect 9896 -140 9902 -70
rect 10222 -160 10274 -154
rect 10222 -200 10228 -160
rect 10228 -200 10268 -160
rect 10268 -200 10274 -160
rect 10222 -206 10274 -200
rect 10040 -236 10092 -230
rect 10040 -276 10046 -236
rect 10046 -276 10086 -236
rect 10086 -276 10092 -236
rect 10040 -282 10092 -276
<< metal2 >>
rect -182 399 216 451
rect 5297 400 5306 456
rect 5362 400 5371 456
rect 10040 380 10092 390
rect -179 277 449 327
rect 1936 231 1996 240
rect 1936 162 1996 171
rect 3874 231 3934 240
rect 3874 162 3934 171
rect 452 129 512 138
rect 452 60 512 69
rect 2386 129 2446 138
rect 2386 60 2446 69
rect 4316 129 4376 138
rect 4316 60 4376 69
rect 281 24 341 33
rect 281 -45 341 -36
rect 2213 24 2273 33
rect 2213 -45 2273 -36
rect 4145 27 4205 36
rect 4145 -42 4205 -33
rect 1770 -76 1830 -67
rect 1770 -145 1830 -136
rect 3702 -75 3762 -66
rect 3702 -144 3762 -135
rect 4829 -231 4879 325
rect 5806 231 5866 240
rect 5806 162 5866 171
rect 7738 231 7798 240
rect 7738 162 7798 171
rect 9670 231 9730 240
rect 9670 162 9730 171
rect 9850 236 9902 246
rect 9850 156 9902 166
rect 6248 129 6308 138
rect 6248 60 6308 69
rect 8180 129 8240 138
rect 8180 60 8240 69
rect 6076 27 6136 36
rect 6076 -42 6136 -33
rect 8014 27 8074 36
rect 8014 -42 8074 -33
rect 9851 -60 9901 156
rect 5634 -75 5694 -66
rect 5634 -144 5694 -135
rect 7564 -75 7624 -66
rect 7564 -144 7624 -135
rect 9498 -75 9558 -66
rect 9498 -144 9558 -135
rect 9850 -70 9902 -60
rect 9850 -150 9902 -140
rect 9851 -181 9901 -150
rect 9699 -231 9901 -181
rect 10040 -230 10092 328
rect 5304 -299 5364 -290
rect 5304 -368 5364 -359
rect 10040 -872 10092 -282
rect 10222 302 10274 312
rect 10222 -154 10274 250
rect 10222 -864 10274 -206
<< via2 >>
rect 5306 400 5362 456
rect 1936 171 1996 231
rect 3874 171 3934 231
rect 452 69 512 129
rect 2386 69 2446 129
rect 4316 69 4376 129
rect 281 -36 341 24
rect 2213 -36 2273 24
rect 4145 -33 4205 27
rect 1770 -136 1830 -76
rect 3702 -135 3762 -75
rect 5806 171 5866 231
rect 7738 171 7798 231
rect 9670 171 9730 231
rect 6248 69 6308 129
rect 8180 69 8240 129
rect 6076 -33 6136 27
rect 8014 -33 8074 27
rect 5634 -135 5694 -75
rect 7564 -135 7624 -75
rect 9498 -135 9558 -75
rect 5304 -359 5364 -299
<< metal3 >>
rect 281 29 341 956
rect 1936 236 1996 956
rect 1931 231 2001 236
rect 1931 171 1936 231
rect 1996 171 2001 231
rect 1931 166 2001 171
rect 447 129 517 134
rect 447 69 452 129
rect 512 69 517 129
rect 447 64 517 69
rect 276 24 346 29
rect 276 -36 281 24
rect 341 -36 346 24
rect 276 -41 346 -36
rect 452 -873 512 64
rect 2213 29 2273 956
rect 3874 236 3934 956
rect 3869 231 3939 236
rect 3869 171 3874 231
rect 3934 171 3939 231
rect 3869 166 3939 171
rect 2381 129 2451 134
rect 2381 69 2386 129
rect 2446 69 2451 129
rect 2381 64 2451 69
rect 2208 24 2278 29
rect 2208 -36 2213 24
rect 2273 -36 2278 24
rect 2208 -41 2278 -36
rect 1765 -76 1835 -71
rect 1765 -136 1770 -76
rect 1830 -136 1835 -76
rect 1765 -141 1835 -136
rect 1770 -873 1830 -141
rect 2386 -873 2446 64
rect 4145 32 4205 956
rect 5301 456 5367 461
rect 5301 400 5306 456
rect 5362 400 5367 456
rect 5301 395 5367 400
rect 4311 129 4381 134
rect 4311 69 4316 129
rect 4376 69 4381 129
rect 4311 64 4381 69
rect 4140 27 4210 32
rect 4140 -33 4145 27
rect 4205 -33 4210 27
rect 4140 -38 4210 -33
rect 3697 -75 3767 -70
rect 3697 -135 3702 -75
rect 3762 -135 3767 -75
rect 3697 -140 3767 -135
rect 3702 -873 3762 -140
rect 4316 -873 4376 64
rect 5304 -294 5364 395
rect 5806 236 5866 956
rect 5801 231 5871 236
rect 5801 171 5806 231
rect 5866 171 5871 231
rect 5801 166 5871 171
rect 6076 32 6136 956
rect 7738 236 7798 956
rect 7733 231 7803 236
rect 7733 171 7738 231
rect 7798 171 7803 231
rect 7733 166 7803 171
rect 6243 129 6313 134
rect 6243 69 6248 129
rect 6308 69 6313 129
rect 6243 64 6313 69
rect 6071 27 6141 32
rect 6071 -33 6076 27
rect 6136 -33 6141 27
rect 6071 -38 6141 -33
rect 5629 -75 5699 -70
rect 5629 -135 5634 -75
rect 5694 -135 5699 -75
rect 5629 -140 5699 -135
rect 5299 -299 5369 -294
rect 5299 -359 5304 -299
rect 5364 -359 5369 -299
rect 5299 -364 5369 -359
rect 5634 -873 5694 -140
rect 6248 -873 6308 64
rect 8014 32 8074 956
rect 9670 236 9730 956
rect 9665 231 9735 236
rect 9665 171 9670 231
rect 9730 171 9735 231
rect 9665 166 9735 171
rect 8175 129 8245 134
rect 8175 69 8180 129
rect 8240 69 8245 129
rect 8175 64 8245 69
rect 8009 27 8079 32
rect 8009 -33 8014 27
rect 8074 -33 8079 27
rect 8009 -38 8079 -33
rect 7559 -75 7629 -70
rect 7559 -135 7564 -75
rect 7624 -135 7629 -75
rect 7559 -140 7629 -135
rect 7564 -873 7624 -140
rect 8180 -873 8240 64
rect 9493 -75 9563 -70
rect 9493 -135 9498 -75
rect 9558 -135 9563 -75
rect 9493 -140 9563 -135
rect 9498 -872 9558 -140
use and_latch  and_latch_0
timestamp 1730774538
transform -1 0 29994 0 1 -16
box 19662 -528 20198 112
use and_latch  and_latch_1
timestamp 1730774538
transform -1 0 29994 0 -1 112
box 19662 -528 20198 112
use flip_flop_5_latch  flip_flop_5_latch_0
timestamp 1730776770
transform 1 0 342 0 -1 -974
box -205 -1614 9531 -974
use flip_flop_5_latch  flip_flop_5_latch_1
timestamp 1730776770
transform -1 0 9668 0 1 1070
box -205 -1614 9531 -974
<< labels >>
flabel metal2 10250 -850 10250 -850 0 FreeSans 800 0 0 0 FINAL
port 0 nsew
flabel metal2 10066 -754 10066 -754 0 FreeSans 800 0 0 0 CLKS
port 1 nsew
flabel metal1 -54 -504 -54 -504 0 FreeSans 800 0 0 0 VSSD
port 2 nsew
flabel metal1 -54 48 -54 48 0 FreeSans 800 0 0 0 VDDD
port 3 nsew
flabel metal2 -164 424 -164 424 0 FreeSans 800 0 0 0 EN
port 4 nsew
flabel metal2 -170 290 -170 290 0 FreeSans 800 0 0 0 CK
port 5 nsew
flabel metal3 1962 930 1968 930 0 FreeSans 800 0 0 0 DOUT[1]
port 8 nsew
flabel metal3 2248 718 2254 718 0 FreeSans 800 0 0 0 DOUT[2]
port 9 nsew
flabel metal3 3904 936 3910 936 0 FreeSans 800 0 0 0 DOUT[3]
port 10 nsew
flabel metal3 4176 714 4182 714 0 FreeSans 800 0 0 0 DOUT[4]
port 11 nsew
flabel metal3 5834 930 5840 930 0 FreeSans 800 0 0 0 DOUT[5]
port 12 nsew
flabel metal3 6110 712 6116 712 0 FreeSans 800 0 0 0 DOUT[6]
port 13 nsew
flabel metal3 7758 918 7764 918 0 FreeSans 800 0 0 0 DOUT[7]
port 14 nsew
flabel metal3 8044 714 8050 714 0 FreeSans 800 0 0 0 DOUT[8]
port 15 nsew
flabel metal3 9696 922 9702 922 0 FreeSans 800 0 0 0 DOUT[9]
port 16 nsew
flabel metal3 1802 -828 1802 -828 0 FreeSans 800 0 0 0 SWP[0]
port 17 nsew
flabel metal3 474 -846 474 -846 0 FreeSans 800 0 0 0 SWP[1]
port 18 nsew
flabel metal3 3736 -832 3736 -832 0 FreeSans 800 0 0 0 SWP[2]
port 19 nsew
flabel metal3 2412 -836 2412 -836 0 FreeSans 800 0 0 0 SWP[3]
port 20 nsew
flabel metal3 5666 -848 5666 -848 0 FreeSans 800 0 0 0 SWP[4]
port 21 nsew
flabel metal3 4342 -834 4342 -834 0 FreeSans 800 0 0 0 SWP[5]
port 22 nsew
flabel metal3 7598 -848 7598 -848 0 FreeSans 800 0 0 0 SWP[6]
port 23 nsew
flabel metal3 6278 -838 6278 -838 0 FreeSans 800 0 0 0 SWP[7]
port 24 nsew
flabel metal3 9528 -846 9528 -846 0 FreeSans 800 0 0 0 SWP[8]
port 25 nsew
flabel metal3 8212 -852 8212 -838 0 FreeSans 800 0 0 0 SWP[9]
port 26 nsew
flabel metal3 314 924 314 938 0 FreeSans 800 0 0 0 DOUT[0]
port 27 nsew
flabel metal1 -28 598 -28 598 0 FreeSans 800 0 0 0 VSSD
port 28 nsew
<< end >>
