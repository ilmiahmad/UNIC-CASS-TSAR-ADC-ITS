magic
tech sky130A
magscale 1 2
timestamp 1727318435
<< nwell >>
rect 234 2695 699 3216
rect 7422 2695 7867 3216
rect 235 2088 700 2089
rect 235 1879 710 2088
rect 235 1568 700 1879
rect 7424 1566 7866 2088
<< pwell >>
rect 234 2118 699 2639
rect 7414 2116 7867 2636
rect 7422 2115 7867 2116
rect 234 991 843 1511
rect 235 988 843 991
rect 7421 988 7866 1510
rect 331 987 843 988
<< viali >>
rect 7498 2648 7534 2684
rect 7664 2646 7702 2684
rect 7536 2528 7572 2562
rect 404 1528 438 1562
rect 584 1528 618 1562
rect 532 1396 570 1434
<< metal1 >>
rect 233 3140 7866 3216
rect 7460 2929 7736 3140
rect 7312 2688 7548 2708
rect 7658 2698 7722 2704
rect 7658 2696 7664 2698
rect 7312 2632 7330 2688
rect 7396 2684 7548 2688
rect 7396 2648 7498 2684
rect 7534 2648 7548 2684
rect 7396 2632 7548 2648
rect 7656 2646 7664 2696
rect 7716 2696 7722 2698
rect 7716 2646 7742 2696
rect 7656 2634 7742 2646
rect 7312 2608 7548 2632
rect 234 2439 639 2518
rect 719 2439 729 2518
rect 7513 2513 7523 2573
rect 7583 2513 7593 2573
rect 7460 2192 7736 2413
rect 234 2116 685 2192
rect 7415 2116 7773 2192
rect 234 1064 294 2116
rect 7806 2088 7866 3140
rect 331 2012 931 2088
rect 7410 2012 7866 2088
rect 369 1802 645 2012
rect 390 1570 452 1576
rect 388 1518 394 1570
rect 446 1518 452 1570
rect 388 1510 452 1518
rect 557 1562 786 1580
rect 557 1528 584 1562
rect 618 1560 786 1562
rect 618 1528 648 1560
rect 557 1502 648 1528
rect 700 1502 786 1560
rect 557 1480 786 1502
rect 511 1386 521 1446
rect 581 1386 591 1446
rect 369 1064 645 1275
rect 234 986 7867 1064
<< via1 >>
rect 7330 2632 7396 2688
rect 7664 2684 7716 2698
rect 7664 2646 7702 2684
rect 7702 2646 7716 2684
rect 639 2439 719 2518
rect 7523 2562 7583 2573
rect 7523 2528 7536 2562
rect 7536 2528 7572 2562
rect 7572 2528 7583 2562
rect 7523 2513 7583 2528
rect 394 1562 446 1570
rect 394 1528 404 1562
rect 404 1528 438 1562
rect 438 1528 446 1562
rect 394 1518 446 1528
rect 648 1502 700 1560
rect 521 1434 581 1446
rect 521 1396 532 1434
rect 532 1396 570 1434
rect 570 1396 581 1434
rect 521 1386 581 1396
<< metal2 >>
rect 5702 2876 5782 2886
rect 234 2797 783 2876
rect 5702 2786 5782 2796
rect 7322 2698 7402 2708
rect 521 2598 686 2648
rect 7656 2698 7786 2704
rect 7656 2646 7664 2698
rect 7716 2646 7786 2698
rect 7656 2634 7786 2646
rect 7322 2608 7402 2618
rect 390 1572 452 1576
rect 378 1570 452 1572
rect 378 1518 394 1570
rect 446 1518 452 1570
rect 378 1510 452 1518
rect 378 1260 430 1510
rect 521 1446 581 2598
rect 7523 2573 7583 2583
rect 639 2518 719 2528
rect 639 2429 719 2439
rect 1435 2518 1515 2528
rect 1435 2429 1515 2439
rect 5704 1748 5784 1758
rect 5704 1658 5784 1668
rect 632 1570 712 1580
rect 7523 1520 7583 2513
rect 632 1480 712 1490
rect 7423 1470 7583 1520
rect 521 1376 581 1386
rect 1434 1390 1514 1400
rect 1434 1300 1514 1310
rect 7734 1260 7786 2634
rect 216 1208 7786 1260
<< via2 >>
rect 5702 2796 5782 2876
rect 7322 2688 7402 2698
rect 7322 2632 7330 2688
rect 7330 2632 7396 2688
rect 7396 2632 7402 2688
rect 7322 2618 7402 2632
rect 1435 2439 1515 2518
rect 5704 1668 5784 1748
rect 632 1560 712 1570
rect 632 1502 648 1560
rect 648 1502 700 1560
rect 700 1502 712 1560
rect 632 1490 712 1502
rect 1434 1310 1514 1390
<< metal3 >>
rect 5692 2876 5794 2884
rect 5692 2796 5702 2876
rect 5782 2796 5794 2876
rect 1424 2518 1526 2523
rect 1424 2439 1435 2518
rect 1515 2439 1526 2518
rect 208 1570 722 1576
rect 208 1490 632 1570
rect 712 1490 722 1570
rect 208 1486 722 1490
rect 622 1485 722 1486
rect 1424 1390 1526 2439
rect 5692 1748 5794 2796
rect 7312 2702 7412 2703
rect 7312 2698 7867 2702
rect 7312 2618 7322 2698
rect 7402 2618 7867 2698
rect 7312 2612 7867 2618
rect 5692 1668 5704 1748
rect 5784 1668 5794 1748
rect 5692 1661 5794 1668
rect 1424 1310 1434 1390
rect 1514 1310 1526 1390
rect 1424 1300 1526 1310
use epc_delay_line  x1
timestamp 1727241376
transform 1 0 628 0 1 1904
box 53 212 6795 1312
use epc_delay_line  x2
timestamp 1727241376
transform -1 0 7477 0 1 776
box 53 212 6795 1312
use sky130_fd_sc_hd__nand2_1  x9 /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 369 0 1 1306
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x10
timestamp 1710522493
transform -1 0 7736 0 1 2433
box -38 -48 314 592
<< labels >>
flabel metal1 268 3164 300 3194 0 FreeSans 320 0 0 0 VDDA
port 0 nsew
flabel metal3 312 1524 344 1554 0 FreeSans 320 0 0 0 OUTN
port 1 nsew
flabel metal1 278 1010 310 1040 0 FreeSans 320 0 0 0 VSSA
port 3 nsew
flabel metal3 7815 2646 7840 2673 0 FreeSans 320 0 0 0 OUTP
port 7 nsew
flabel metal2 s 218 1234 218 1234 0 FreeSans 320 0 0 0 START
port 9 nsew
flabel metal1 256 2466 281 2493 0 FreeSans 320 0 0 0 VN
port 5 nsew
flabel metal2 259 2826 284 2853 0 FreeSans 320 0 0 0 VP
port 4 nsew
<< end >>
