magic
tech sky130A
magscale 1 2
timestamp 1731182005
<< nwell >>
rect -1174 918 1367 1956
rect 199 905 372 918
<< pwell >>
rect -872 200 1164 864
<< viali >>
rect -1042 1902 -268 1936
rect 806 1902 1580 1936
rect 483 1027 517 1061
rect -62 859 -28 893
rect 106 859 140 893
rect 396 859 430 893
rect 564 859 598 893
rect 109 737 143 771
rect 525 737 559 771
rect -1042 216 -686 250
rect 1224 216 1580 250
<< metal1 >>
rect -1174 1936 1712 1972
rect -1174 1902 -1042 1936
rect -268 1902 806 1936
rect 1580 1902 1712 1936
rect -1174 1875 1712 1902
rect -1062 1728 -1052 1794
rect -996 1728 -986 1794
rect -405 1782 -355 1875
rect -1184 1412 -1174 1478
rect -1118 1412 -1108 1478
rect -1062 1412 -1052 1478
rect -996 1412 -986 1478
rect -955 1466 -905 1740
rect -324 1728 -314 1794
rect -258 1728 -248 1794
rect -314 1656 -258 1728
rect -324 1590 -314 1656
rect -258 1590 -248 1656
rect -1174 424 -1122 1412
rect -407 1322 -355 1425
rect -324 1412 -314 1478
rect -258 1412 -248 1478
rect -417 1270 -407 1322
rect -355 1270 -345 1322
rect -208 1270 -198 1322
rect -146 1270 -136 1322
rect -1052 882 -996 1162
rect -417 1150 -407 1202
rect -355 1150 -345 1202
rect -814 1006 -764 1108
rect -314 1096 -258 1162
rect -198 1006 -146 1270
rect 573 1236 636 1875
rect 786 1728 796 1794
rect 852 1728 862 1794
rect 893 1782 943 1875
rect 674 1656 730 1666
rect 674 1590 687 1656
rect 744 1590 754 1656
rect 674 1478 730 1590
rect 664 1412 674 1478
rect 730 1412 740 1478
rect 786 1412 796 1478
rect 852 1412 862 1478
rect 1443 1466 1493 1740
rect 1534 1728 1590 1794
rect 893 1322 945 1424
rect 1524 1412 1534 1478
rect 1590 1412 1600 1478
rect 1646 1412 1656 1478
rect 1712 1412 1722 1478
rect 674 1270 684 1322
rect 736 1270 746 1322
rect 883 1270 893 1322
rect 945 1270 955 1322
rect -98 1184 -72 1236
rect -20 1184 113 1236
rect 165 1184 389 1236
rect 441 1184 573 1236
rect 625 1184 636 1236
rect -98 1140 636 1184
rect 461 1077 471 1100
rect 90 1044 471 1077
rect 529 1044 539 1100
rect 90 1027 483 1044
rect 517 1027 529 1044
rect 90 1010 529 1027
rect -824 954 -814 1006
rect -758 954 -748 1006
rect -208 954 -198 1006
rect -146 954 -136 1006
rect -1062 830 -1052 882
rect -996 830 -986 882
rect -1052 674 -996 830
rect -814 728 -764 954
rect -91 922 -81 976
rect -14 922 -4 976
rect -81 893 -14 922
rect -81 859 -62 893
rect -28 859 -14 893
rect -81 853 -14 859
rect 90 893 157 1010
rect 90 859 106 893
rect 140 859 157 893
rect 90 843 157 859
rect 238 893 446 904
rect 238 859 396 893
rect 430 859 446 893
rect 238 848 446 859
rect 238 787 294 848
rect 538 843 548 909
rect 615 843 625 909
rect 684 882 736 1270
rect 796 1096 852 1162
rect 883 1150 893 1202
rect 945 1150 955 1202
rect 1302 882 1352 1108
rect 1534 1006 1590 1162
rect 1524 954 1534 1006
rect 1590 954 1600 1006
rect 674 830 684 882
rect 736 830 746 882
rect 1286 830 1296 882
rect 1352 830 1362 882
rect -1184 358 -1174 424
rect -1118 358 -1108 424
rect -1072 358 -1062 424
rect -1006 358 -996 424
rect -814 412 -764 686
rect -732 674 -676 740
rect 87 731 97 787
rect 155 731 294 787
rect 503 726 513 782
rect 571 726 581 782
rect -98 596 637 692
rect 1214 674 1270 740
rect 1302 728 1352 830
rect -814 277 -764 370
rect -732 358 -676 424
rect 573 277 636 596
rect 1214 358 1270 424
rect 1302 412 1352 686
rect 1534 674 1590 954
rect 1660 424 1712 1412
rect 1302 277 1352 368
rect 1534 358 1544 424
rect 1600 358 1610 424
rect 1646 358 1656 424
rect 1712 358 1722 424
rect -1174 250 1712 277
rect -1174 216 -1042 250
rect -686 216 1224 250
rect 1580 216 1712 250
rect -1174 180 1712 216
<< via1 >>
rect -1052 1728 -996 1794
rect -1174 1412 -1118 1478
rect -1052 1412 -996 1478
rect -314 1728 -258 1794
rect -314 1590 -258 1656
rect -314 1412 -258 1478
rect -407 1270 -355 1322
rect -198 1270 -146 1322
rect -407 1150 -355 1202
rect 796 1728 852 1794
rect 687 1590 744 1656
rect 674 1412 730 1478
rect 796 1412 852 1478
rect 1534 1412 1590 1478
rect 1656 1412 1712 1478
rect 684 1270 736 1322
rect 893 1270 945 1322
rect -72 1184 -20 1236
rect 113 1184 165 1236
rect 389 1184 441 1236
rect 573 1184 625 1236
rect 471 1061 529 1100
rect 471 1044 483 1061
rect 483 1044 517 1061
rect 517 1044 529 1061
rect -814 954 -758 1006
rect -198 954 -146 1006
rect -1052 830 -996 882
rect -81 922 -14 976
rect 548 893 615 909
rect 548 859 564 893
rect 564 859 598 893
rect 598 859 615 893
rect 548 843 615 859
rect 893 1150 945 1202
rect 1534 954 1590 1006
rect 684 830 736 882
rect 1296 830 1352 882
rect -1174 358 -1118 424
rect -1062 358 -1006 424
rect 97 771 155 787
rect 97 737 109 771
rect 109 737 143 771
rect 143 737 155 771
rect 97 731 155 737
rect 513 771 571 782
rect 513 737 525 771
rect 525 737 559 771
rect 559 737 571 771
rect 513 726 571 737
rect 1544 358 1600 424
rect 1656 358 1712 424
<< metal2 >>
rect -1052 1794 -996 1804
rect -1174 1728 -1052 1794
rect -1052 1718 -996 1728
rect -314 1794 -258 1804
rect -314 1718 -258 1728
rect 796 1794 852 1804
rect 796 1718 852 1728
rect -314 1656 -258 1666
rect 687 1656 744 1666
rect -258 1590 687 1656
rect -314 1580 -258 1590
rect 687 1580 744 1590
rect -1174 1478 -1118 1488
rect -1052 1478 -996 1488
rect -1118 1412 -1052 1478
rect -1174 1402 -1118 1412
rect -1052 1402 -996 1412
rect -314 1478 -258 1488
rect -192 1478 -136 1488
rect -258 1412 -192 1478
rect -314 1402 -258 1412
rect -192 1402 -136 1412
rect 674 1478 730 1488
rect 796 1478 852 1488
rect 730 1412 796 1478
rect 674 1402 730 1412
rect 796 1402 852 1412
rect 1534 1478 1590 1488
rect 1656 1478 1712 1488
rect 1590 1412 1656 1478
rect 1534 1402 1590 1412
rect 1656 1402 1712 1412
rect -407 1322 -355 1332
rect -198 1322 -146 1332
rect -355 1270 -198 1322
rect -407 1260 -355 1270
rect -198 1260 -146 1270
rect 684 1322 736 1332
rect 893 1322 945 1332
rect 736 1270 893 1322
rect 684 1260 736 1270
rect 893 1260 945 1270
rect -72 1236 -20 1246
rect -407 1202 -355 1212
rect -355 1184 -72 1202
rect 113 1236 165 1246
rect -20 1184 113 1202
rect 389 1236 441 1246
rect 165 1184 389 1202
rect 573 1236 625 1246
rect 441 1184 573 1202
rect 893 1202 945 1212
rect 625 1184 893 1202
rect -355 1150 893 1184
rect -407 1140 -355 1150
rect 893 1140 945 1150
rect 471 1100 529 1110
rect 471 1034 529 1044
rect -814 1006 -758 1016
rect -198 1006 -146 1016
rect 1534 1006 1590 1016
rect -758 954 -198 1006
rect -146 976 1534 1006
rect -146 954 -81 976
rect -814 944 -758 954
rect -198 944 -146 954
rect -14 954 1534 976
rect 1534 944 1590 954
rect -81 912 -14 922
rect 548 909 615 919
rect -1052 882 -996 892
rect -996 843 548 882
rect 684 882 736 892
rect 1296 882 1352 892
rect 615 843 684 882
rect -996 830 684 843
rect 736 830 1296 882
rect -1052 820 -996 830
rect 684 820 736 830
rect 1296 820 1352 830
rect 97 787 155 797
rect -268 735 97 787
rect 97 721 155 731
rect 513 782 571 792
rect 571 726 806 782
rect 513 716 571 726
rect -1174 424 -1118 434
rect -1062 424 -1006 434
rect -1118 358 -1062 424
rect -1174 348 -1118 358
rect -1062 348 -1006 358
rect 1544 424 1600 434
rect 1656 424 1712 434
rect 1600 358 1656 424
rect 1544 348 1600 358
rect 1656 348 1712 358
<< via2 >>
rect 796 1728 852 1794
rect -192 1412 -136 1478
<< metal3 >>
rect 776 1804 872 1815
rect -212 1718 -202 1804
rect -126 1718 -116 1804
rect 776 1718 786 1804
rect 862 1718 872 1804
rect -202 1478 -126 1718
rect 776 1708 872 1718
rect -202 1412 -192 1478
rect -136 1412 -126 1478
rect -202 1407 -126 1412
<< via3 >>
rect -202 1718 -126 1804
rect 786 1794 862 1804
rect 786 1728 796 1794
rect 796 1728 852 1794
rect 852 1728 862 1794
rect 786 1718 862 1728
<< metal4 >>
rect -203 1804 863 1805
rect -203 1718 -202 1804
rect -126 1718 786 1804
rect 862 1718 863 1804
rect -203 1717 863 1718
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -98 0 1 644
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1704896540
transform 1 0 360 0 1 644
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_R8XU9D  XM1
timestamp 1730240227
transform 0 1 -655 -1 0 1761
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM2
timestamp 1730240227
transform 0 -1 -655 1 0 1445
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM3
timestamp 1730240227
transform 0 1 1193 -1 0 1761
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM4
timestamp 1730240227
transform 0 1 1193 -1 0 1445
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM5
timestamp 1730240227
transform 0 1 -655 -1 0 1129
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_TGNW9T  XM6
timestamp 1730240227
transform 0 -1 -864 1 0 707
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM7
timestamp 1730240227
transform 0 1 -864 -1 0 391
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_R8XU9D  XM8
timestamp 1730240227
transform 0 1 1193 -1 0 1129
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_TGNW9T  XM9
timestamp 1730240227
transform 0 1 1402 -1 0 707
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM10
timestamp 1730240227
transform 0 1 1402 -1 0 391
box -211 -310 211 310
<< labels >>
flabel metal2 -262 735 -210 787 0 FreeSans 800 0 0 0 OUT
port 0 nsew
flabel metal2 750 726 806 782 0 FreeSans 800 0 0 0 OUTN
port 1 nsew
flabel metal2 -1118 1728 -1052 1794 0 FreeSans 800 0 0 0 INN
port 2 nsew
flabel metal2 -1118 1412 -1052 1478 0 FreeSans 800 0 0 0 INP
port 3 nsew
flabel metal1 237 1875 336 1972 0 FreeSans 800 0 0 0 VDD
port 4 nsew
flabel metal1 252 180 351 277 0 FreeSans 800 0 0 0 VSS
port 5 nsew
<< end >>
