magic
tech sky130A
magscale 1 2
timestamp 1731351601
<< dnwell >>
rect -12808 30642 -12778 30984
rect -12808 30000 -12778 30342
rect 68477 27523 71679 33313
<< nwell >>
rect -12808 30699 -12778 30984
rect -12917 30133 -11985 30699
rect -12808 30000 -12778 30133
<< metal1 >>
rect -10804 61777 -1450 61961
rect -1266 61777 67606 61961
rect 67790 61777 67800 61961
rect -10804 61552 68087 61604
rect 68139 61552 68149 61604
rect -10804 61410 67915 61462
rect 67967 61410 67977 61462
rect -10804 61095 68277 61227
rect 68406 61095 68416 61227
rect -10804 60553 133 60554
rect -10804 60369 -26 60553
rect 158 60369 168 60553
rect -10804 60036 186 60220
rect 370 60036 380 60220
rect -10804 59715 398 59899
rect 582 59715 592 59899
rect 67002 33591 67012 33791
rect 67212 33591 71819 33791
rect 72019 33591 72029 33791
rect -11892 33279 -398 33391
rect -510 27548 -398 33279
rect 71809 31715 71819 31915
rect 72019 31715 72029 31915
rect 68267 30832 68277 30961
rect 68406 30832 68708 30961
rect 71819 30775 72019 31715
rect 71356 30575 72019 30775
rect 67906 30492 67916 30544
rect 67968 30492 68679 30544
rect 68076 30392 68086 30444
rect 68138 30392 68678 30444
rect 71053 30061 72019 30261
rect 71819 29121 72019 30061
rect 71809 28921 71819 29121
rect 72019 28921 72029 29121
rect -12139 27436 -398 27548
rect 67676 27523 67686 27627
rect 67790 27523 68701 27627
rect -1412 27298 -1300 27436
rect -1418 27186 -1412 27298
rect -1300 27186 -1294 27298
rect 71819 27244 72019 27245
rect 67002 27044 67012 27244
rect 67212 27044 71819 27244
rect 72019 27044 72029 27244
rect -1460 -944 -1450 -760
rect -1266 -944 68222 -760
rect 68406 -944 68416 -760
<< via1 >>
rect -1450 61777 -1266 61961
rect 67606 61777 67790 61961
rect 68087 61552 68139 61604
rect 67915 61410 67967 61462
rect 68277 61095 68406 61227
rect -26 60369 158 60553
rect 186 60036 370 60220
rect 398 59715 582 59899
rect 67012 33591 67212 33791
rect 71819 33591 72019 33791
rect 71819 31715 72019 31915
rect 68277 30832 68406 30961
rect 67916 30492 67968 30544
rect 68086 30392 68138 30444
rect 71819 28921 72019 29121
rect 67686 27523 67790 27627
rect -1412 27186 -1300 27298
rect 67012 27044 67212 27244
rect 71819 27044 72019 27244
rect -1450 -944 -1266 -760
rect 68222 -944 68406 -760
<< metal2 >>
rect -1450 61961 -1266 61971
rect -9150 35052 -8966 60807
rect -9150 34859 -8966 34868
rect -8650 35052 -8466 60807
rect -8650 34859 -8466 34868
rect -8150 35052 -7966 60807
rect -8150 34859 -7966 34868
rect -7650 35052 -7466 60807
rect -7650 34859 -7466 34868
rect -7150 35052 -6966 60807
rect -7150 34859 -6966 34868
rect -6450 35394 -6266 60807
rect -6450 35308 -6396 35394
rect -6310 35308 -6266 35394
rect -6450 33915 -6266 35308
rect -5950 35550 -5766 60807
rect -5950 35464 -5898 35550
rect -5812 35464 -5766 35550
rect -5950 33915 -5766 35464
rect -5450 35706 -5266 60807
rect -5450 35620 -5402 35706
rect -5316 35620 -5266 35706
rect -5450 33915 -5266 35620
rect -4950 35862 -4766 60807
rect -4950 35776 -4903 35862
rect -4817 35776 -4766 35862
rect -4950 33915 -4766 35776
rect -4450 36018 -4266 60807
rect -4450 35932 -4405 36018
rect -4319 35932 -4266 36018
rect -4450 33915 -4266 35932
rect -3950 36174 -3766 60807
rect -3950 36088 -3903 36174
rect -3817 36088 -3766 36174
rect -3950 33915 -3766 36088
rect -3450 36330 -3266 60807
rect -3450 36244 -3404 36330
rect -3318 36244 -3266 36330
rect -3450 33915 -3266 36244
rect -2950 36486 -2766 60807
rect -2950 36400 -2905 36486
rect -2819 36400 -2766 36486
rect -2950 33915 -2766 36400
rect -2450 36642 -2266 60807
rect -2450 36556 -2402 36642
rect -2316 36556 -2266 36642
rect -2450 33915 -2266 36556
rect -1950 36798 -1766 60807
rect -1950 36712 -1905 36798
rect -1819 36712 -1766 36798
rect -1950 33915 -1766 36712
rect -1450 33915 -1266 61777
rect 67606 61961 67790 61971
rect 67606 61767 67790 61777
rect -956 33972 -772 60810
rect -238 60807 -54 60817
rect -922 33911 -802 33972
rect -926 33801 -917 33911
rect -807 33801 -798 33911
rect -922 33796 -802 33801
rect -1450 33722 -1266 33731
rect -238 33266 -54 60703
rect -26 60585 158 61101
rect -26 60553 158 60563
rect 186 60521 370 61099
rect 398 60511 582 61098
rect 67012 60807 67196 60817
rect -26 60359 158 60369
rect 186 60220 370 60230
rect 186 60026 370 60036
rect 398 59899 582 59909
rect 398 59705 582 59715
rect 67012 33801 67196 60703
rect 67012 33791 67212 33801
rect 67012 33581 67212 33591
rect -1391 33082 -54 33266
rect -1267 32355 -922 32475
rect -802 32355 -793 32475
rect -580 31739 -317 31835
rect -580 31644 -494 31739
rect -399 31644 -317 31739
rect -580 31559 -317 31644
rect -15790 30981 -15088 31054
rect -15790 30929 -14742 30981
rect -15790 30870 -15088 30929
rect -494 30461 -399 31559
rect -800 30366 -398 30461
rect -15788 29904 -15084 29972
rect -15788 29848 -14674 29904
rect -15788 29788 -15084 29848
rect -1267 28352 -923 28472
rect -803 28352 -794 28472
rect -1592 27563 -54 27747
rect -1412 27298 -1300 27318
rect -1412 27100 -1300 27186
rect -9079 25945 -8895 25954
rect -9079 6 -8895 25761
rect -8579 25945 -8395 25954
rect -8579 6 -8395 25761
rect -8079 25945 -7895 25954
rect -8079 6 -7895 25761
rect -7579 25945 -7395 25954
rect -7579 6 -7395 25761
rect -7079 25945 -6895 25954
rect -7079 6 -6895 25761
rect -6350 25528 -6166 27100
rect -6350 25442 -6304 25528
rect -6218 25442 -6166 25528
rect -6350 29 -6166 25442
rect -5850 25372 -5666 27100
rect -5850 25286 -5800 25372
rect -5714 25286 -5666 25372
rect -5850 29 -5666 25286
rect -5350 25216 -5166 27100
rect -5350 25130 -5299 25216
rect -5213 25130 -5166 25216
rect -5350 29 -5166 25130
rect -4850 25060 -4666 27100
rect -4850 24974 -4796 25060
rect -4710 24974 -4666 25060
rect -4850 29 -4666 24974
rect -4450 24904 -4266 27100
rect -4450 24818 -4400 24904
rect -4314 24818 -4266 24904
rect -4450 29 -4266 24818
rect -3950 24748 -3766 27100
rect -3950 24662 -3899 24748
rect -3813 24662 -3766 24748
rect -3950 29 -3766 24662
rect -3450 24592 -3266 27100
rect -3450 24506 -3402 24592
rect -3316 24506 -3266 24592
rect -3450 29 -3266 24506
rect -2950 24436 -2766 27100
rect -2950 24350 -2902 24436
rect -2816 24350 -2766 24436
rect -2950 29 -2766 24350
rect -2450 24280 -2266 27100
rect -2450 24194 -2399 24280
rect -2313 24194 -2266 24280
rect -2450 29 -2266 24194
rect -1950 24124 -1766 27100
rect -1950 24038 -1902 24124
rect -1816 24038 -1766 24124
rect -1950 29 -1766 24038
rect -1450 -760 -1266 27100
rect -922 27038 -802 27043
rect -926 26928 -917 27038
rect -807 26928 -798 27038
rect -922 26886 -802 26928
rect -952 30 -768 26886
rect -238 134 -54 27563
rect 67686 27627 67790 61767
rect -238 19 -54 29
rect 67012 27244 67212 27254
rect 67012 27034 67212 27044
rect 67012 133 67196 27034
rect 67012 19 67196 29
rect 67686 -750 67790 27523
rect 67915 61462 67967 61901
rect 67915 30554 67967 61410
rect 68087 61604 68139 61907
rect 67915 30544 67968 30554
rect 67915 30492 67916 30544
rect 67915 30482 67968 30492
rect 67915 -750 67967 30482
rect 68087 30454 68139 61552
rect 68086 30444 68139 30454
rect 68138 30392 68139 30444
rect 68086 30382 68139 30392
rect 68087 -750 68139 30382
rect 68277 61227 68406 61905
rect 68277 30961 68406 61095
rect 71819 33791 72019 33801
rect 71819 33581 72019 33591
rect 71819 31915 72019 31925
rect 71819 31705 72019 31715
rect 68277 -750 68406 30832
rect 71341 30831 74799 31031
rect 71356 29805 74799 30005
rect 71819 29121 72019 29131
rect 71819 28911 72019 28921
rect 71819 27244 72019 27254
rect 71819 27034 72019 27044
rect -1450 -954 -1266 -944
rect 68222 -760 68406 -750
rect 68222 -954 68406 -944
<< via2 >>
rect -9150 34868 -8966 35052
rect -8650 34868 -8466 35052
rect -8150 34868 -7966 35052
rect -7650 34868 -7466 35052
rect -7150 34868 -6966 35052
rect -6396 35308 -6310 35394
rect -5898 35464 -5812 35550
rect -5402 35620 -5316 35706
rect -4903 35776 -4817 35862
rect -4405 35932 -4319 36018
rect -3903 36088 -3817 36174
rect -3404 36244 -3318 36330
rect -2905 36400 -2819 36486
rect -2402 36556 -2316 36642
rect -1905 36712 -1819 36798
rect -238 60703 -54 60807
rect -1450 33731 -1266 33915
rect -917 33801 -807 33911
rect 67012 60703 67196 60807
rect -922 32355 -802 32475
rect -494 31644 -399 31739
rect -923 28352 -803 28472
rect -9079 25761 -8895 25945
rect -8579 25761 -8395 25945
rect -8079 25761 -7895 25945
rect -7579 25761 -7395 25945
rect -7079 25761 -6895 25945
rect -6304 25442 -6218 25528
rect -5800 25286 -5714 25372
rect -5299 25130 -5213 25216
rect -4796 24974 -4710 25060
rect -4400 24818 -4314 24904
rect -3899 24662 -3813 24748
rect -3402 24506 -3316 24592
rect -2902 24350 -2816 24436
rect -2399 24194 -2313 24280
rect -1902 24038 -1816 24124
rect -917 26928 -807 27038
rect -238 29 -54 134
rect 67012 29 67196 133
rect 71819 33591 72019 33791
rect 71819 31715 72019 31915
rect 71819 28921 72019 29121
rect 71819 27044 72019 27244
<< metal3 >>
rect -248 60807 -44 60812
rect -248 60703 -238 60807
rect -54 60703 -44 60807
rect -248 60698 -44 60703
rect 67002 60807 67207 60812
rect 67002 60703 67012 60807
rect 67197 60703 67207 60807
rect 67002 60698 67207 60703
rect -2098 36798 215 36803
rect -2098 36712 -1905 36798
rect -1819 36712 215 36798
rect -2098 36707 215 36712
rect -2451 36642 230 36647
rect -2451 36556 -2402 36642
rect -2316 36556 230 36642
rect -2451 36551 230 36556
rect -2950 36486 250 36491
rect -2950 36400 -2905 36486
rect -2819 36400 250 36486
rect -2950 36395 250 36400
rect -3456 36330 255 36335
rect -3456 36244 -3404 36330
rect -3318 36244 255 36330
rect -3456 36239 255 36244
rect -3996 36174 265 36179
rect -3996 36088 -3903 36174
rect -3817 36088 265 36174
rect -3996 36083 265 36088
rect -4448 36018 250 36023
rect -4448 35932 -4405 36018
rect -4319 35932 250 36018
rect -4448 35927 250 35932
rect -4950 35862 196 35867
rect -4950 35776 -4903 35862
rect -4817 35776 196 35862
rect -4950 35771 196 35776
rect -5452 35706 235 35711
rect -5452 35620 -5402 35706
rect -5316 35620 235 35706
rect -5452 35615 235 35620
rect -5948 35550 206 35555
rect -5948 35464 -5898 35550
rect -5812 35464 206 35550
rect -5948 35459 206 35464
rect -6447 35394 206 35399
rect -6447 35308 -6396 35394
rect -6310 35308 206 35394
rect -6447 35303 206 35308
rect -9155 35052 -8961 35057
rect -9155 34868 -9150 35052
rect -8966 34868 -8961 35052
rect -9155 34863 -8961 34868
rect -8655 35052 -8461 35057
rect -8655 34868 -8650 35052
rect -8466 34868 -8461 35052
rect -8655 34863 -8461 34868
rect -8155 35052 -7961 35057
rect -8155 34868 -8150 35052
rect -7966 34868 -7961 35052
rect -8155 34863 -7961 34868
rect -7655 35052 -7461 35057
rect -7655 34868 -7650 35052
rect -7466 34868 -7461 35052
rect -7655 34863 -7461 34868
rect -7155 35052 -6961 35057
rect -7155 34868 -7150 35052
rect -6966 34868 -6961 35052
rect -7155 34863 -6961 34868
rect -9106 30544 -9010 34863
rect -8606 30700 -8510 34863
rect -8100 30856 -8004 34863
rect -7604 31012 -7508 34863
rect -7109 34231 -7013 34863
rect -7110 31168 -7014 34231
rect -1455 33915 -1261 33920
rect -1455 33731 -1450 33915
rect -1266 33731 -1261 33915
rect -1455 33726 -1261 33731
rect -922 33911 -802 33916
rect -922 33801 -917 33911
rect -807 33801 -802 33911
rect -1450 31784 -1266 33726
rect -922 32480 -802 33801
rect 71809 33791 72029 33796
rect 71809 33591 71819 33791
rect 72019 33591 72029 33791
rect 71809 33586 72029 33591
rect -927 32475 -797 32480
rect -927 32355 -922 32475
rect -802 32355 -797 32475
rect -927 32350 -797 32355
rect 71819 31920 72019 33586
rect 71809 31915 72029 31920
rect -1450 31739 -317 31784
rect -1450 31644 -494 31739
rect -399 31644 -317 31739
rect 71809 31715 71819 31915
rect 72019 31715 72029 31915
rect 71809 31710 72029 31715
rect -1450 31600 -317 31644
rect -7110 31072 372 31168
rect -7604 30916 387 31012
rect -8100 30760 446 30856
rect -8606 30604 475 30700
rect -9106 30448 437 30544
rect -9036 30292 331 30388
rect -9036 25950 -8940 30292
rect -8535 30136 380 30232
rect -8535 25950 -8439 30136
rect -8029 29980 224 30076
rect -8029 25950 -7933 29980
rect -7532 29824 434 29920
rect -7532 26041 -7436 29824
rect -7533 25950 -7436 26041
rect -7040 29668 451 29764
rect -7040 25950 -6944 29668
rect 71809 29121 72029 29126
rect 71809 28921 71819 29121
rect 72019 28921 72029 29121
rect 71809 28916 72029 28921
rect -928 28472 -798 28477
rect -928 28352 -923 28472
rect -803 28352 -798 28472
rect -928 28347 -798 28352
rect -923 28251 -802 28347
rect -922 27038 -802 28251
rect 71819 27249 72019 28916
rect 71809 27244 72029 27249
rect 71809 27044 71819 27244
rect 72019 27044 72029 27244
rect 71809 27039 72029 27044
rect -922 26928 -917 27038
rect -807 26928 -802 27038
rect -922 26923 -802 26928
rect -9084 25945 -8890 25950
rect -9084 25761 -9079 25945
rect -8895 25761 -8890 25945
rect -9084 25756 -8890 25761
rect -8584 25945 -8390 25950
rect -8584 25761 -8579 25945
rect -8395 25761 -8390 25945
rect -8584 25756 -8390 25761
rect -8084 25945 -7890 25950
rect -8084 25761 -8079 25945
rect -7895 25761 -7890 25945
rect -8084 25756 -7890 25761
rect -7584 25945 -7390 25950
rect -7584 25761 -7579 25945
rect -7395 25761 -7390 25945
rect -7584 25756 -7390 25761
rect -7084 25945 -6890 25950
rect -7084 25761 -7079 25945
rect -6895 25761 -6890 25945
rect -7084 25756 -6890 25761
rect -7040 25747 -6944 25756
rect -6348 25528 78 25533
rect -6348 25442 -6304 25528
rect -6218 25442 78 25528
rect -6348 25437 78 25442
rect -5848 25372 208 25377
rect -5848 25286 -5800 25372
rect -5714 25286 208 25372
rect -5848 25281 208 25286
rect -5348 25216 188 25221
rect -5348 25130 -5299 25216
rect -5213 25130 188 25216
rect -5348 25125 188 25130
rect -4848 25060 128 25065
rect -4848 24974 -4796 25060
rect -4710 24974 128 25060
rect -4848 24969 128 24974
rect -4448 24904 153 24909
rect -4448 24818 -4400 24904
rect -4314 24818 153 24904
rect -4448 24813 153 24818
rect -3948 24748 148 24753
rect -3948 24662 -3899 24748
rect -3813 24662 148 24748
rect -3948 24657 148 24662
rect -3448 24592 128 24597
rect -3448 24506 -3402 24592
rect -3316 24506 128 24592
rect -3448 24501 128 24506
rect -2951 24436 163 24441
rect -2951 24350 -2902 24436
rect -2816 24350 163 24436
rect -2951 24345 163 24350
rect -2451 24280 173 24285
rect -2451 24194 -2399 24280
rect -2313 24194 173 24280
rect -2451 24189 173 24194
rect -2100 24124 198 24129
rect -2100 24038 -1902 24124
rect -1816 24038 198 24124
rect -2100 24033 198 24038
rect -248 134 -44 139
rect -248 29 -238 134
rect -54 29 -44 134
rect -248 24 -44 29
rect 67002 133 67206 138
rect 67002 29 67012 133
rect 67196 29 67206 133
rect 67002 24 67206 29
<< via3 >>
rect -238 60703 -54 60807
rect 67012 60703 67196 60807
rect 67196 60703 67197 60807
rect -238 29 -54 134
rect 67012 29 67196 133
<< metal4 >>
rect -239 60807 -53 60808
rect 67011 60807 67198 60808
rect -239 60703 -238 60807
rect -54 60703 933 60807
rect 65782 60703 67012 60807
rect 67197 60703 67198 60807
rect -239 60702 -53 60703
rect 67011 60702 67198 60703
rect -239 134 -53 135
rect -239 29 -238 134
rect -54 133 -53 134
rect 67011 133 67197 134
rect -54 29 1187 133
rect 66025 29 67012 133
rect 67196 29 67197 133
rect -239 28 -53 29
rect 67011 28 67197 29
use bsw_diff  bsw_diff_0
timestamp 1731002366
transform 1 0 67704 0 1 34294
box 773 -6771 7052 -981
use cdac_10b  cdac_10b_0
timestamp 1731349849
transform 1 0 -18 0 1 30
box -246 -63 67002 60828
use tdc  tdc_0
timestamp 1731351586
transform -1 0 -5541 0 1 31145
box -4836 -3709 9311 2246
<< labels >>
flabel metal2 -15790 30870 -15606 31054 0 FreeSans 800 0 0 0 COMP_P
port 0 nsew
flabel metal2 -15788 29788 -15604 29972 0 FreeSans 800 0 0 0 COMP_N
port 1 nsew
flabel metal2 -1950 60623 -1766 60807 0 FreeSans 800 270 0 0 SWP[0]
port 2 nsew
flabel metal2 -2450 60623 -2266 60807 0 FreeSans 800 270 0 0 SWP[1]
port 3 nsew
flabel metal2 -2950 60623 -2766 60807 0 FreeSans 800 270 0 0 SWP[2]
port 4 nsew
flabel metal2 -3450 60623 -3266 60807 0 FreeSans 800 270 0 0 SWP[3]
port 5 nsew
flabel metal2 -3950 60623 -3766 60807 0 FreeSans 800 270 0 0 SWP[4]
port 6 nsew
flabel metal2 -4450 60623 -4266 60807 0 FreeSans 800 270 0 0 SWP[5]
port 7 nsew
flabel metal2 -4950 60623 -4766 60807 0 FreeSans 800 270 0 0 SWP[6]
port 8 nsew
flabel metal2 -5450 60623 -5266 60807 0 FreeSans 800 270 0 0 SWP[7]
port 9 nsew
flabel metal2 -5950 60623 -5766 60807 0 FreeSans 800 270 0 0 SWP[8]
port 10 nsew
flabel metal2 -6450 60623 -6266 60807 0 FreeSans 800 270 0 0 SWP[9]
port 11 nsew
flabel metal2 -1950 29 -1766 213 0 FreeSans 800 270 0 0 SWN[0]
port 12 nsew
flabel metal2 -2450 29 -2266 213 0 FreeSans 800 270 0 0 SWN[1]
port 13 nsew
flabel metal2 -2950 29 -2766 213 0 FreeSans 800 270 0 0 SWN[2]
port 14 nsew
flabel metal2 -3450 32 -3266 216 0 FreeSans 800 270 0 0 SWN[3]
port 15 nsew
flabel metal2 -3950 29 -3766 213 0 FreeSans 800 270 0 0 SWN[4]
port 16 nsew
flabel metal2 -4450 29 -4266 213 0 FreeSans 800 270 0 0 SWN[5]
port 17 nsew
flabel metal2 -4850 29 -4666 213 0 FreeSans 800 270 0 0 SWN[6]
port 18 nsew
flabel metal2 -5350 32 -5166 216 0 FreeSans 800 270 0 0 SWN[7]
port 19 nsew
flabel metal2 -5850 29 -5666 213 0 FreeSans 800 270 0 0 SWN[8]
port 20 nsew
flabel metal2 -6350 41 -6166 225 0 FreeSans 800 270 0 0 SWN[9]
port 21 nsew
flabel metal2 -7079 6 -6895 190 0 FreeSans 800 270 0 0 CF[0]
port 22 nsew
flabel metal2 -7579 6 -7395 190 0 FreeSans 800 270 0 0 CF[1]
port 23 nsew
flabel metal2 -8079 6 -7895 190 0 FreeSans 800 270 0 0 CF[2]
port 24 nsew
flabel metal2 -8579 6 -8395 190 0 FreeSans 800 270 0 0 CF[3]
port 25 nsew
flabel metal2 -9079 6 -8895 190 0 FreeSans 800 270 0 0 CF[4]
port 26 nsew
flabel metal2 -9150 60623 -8966 60807 0 FreeSans 800 270 0 0 CF[5]
port 27 nsew
flabel metal2 -8650 60623 -8466 60807 0 FreeSans 800 270 0 0 CF[6]
port 28 nsew
flabel metal2 -8150 60623 -7966 60807 0 FreeSans 800 270 0 0 CF[7]
port 29 nsew
flabel metal2 -7650 60623 -7466 60807 0 FreeSans 800 270 0 0 CF[8]
port 30 nsew
flabel metal2 -7150 60623 -6966 60807 0 FreeSans 800 270 0 0 CF[9]
port 31 nsew
flabel metal2 -952 30 -768 214 0 FreeSans 800 270 0 0 CLK
port 32 nsew
flabel metal2 -956 60626 -772 60810 0 FreeSans 800 270 0 0 CLK
port 33 nsew
flabel metal2 -1450 60623 -1266 60807 0 FreeSans 800 270 0 0 VDDA
port 34 nsew
flabel metal2 -1450 29 -1266 213 0 FreeSans 800 270 0 0 VSSA
port 35 nsew
flabel metal2 -26 60917 158 61101 0 FreeSans 800 270 0 0 VCM
port 36 nsew
flabel metal2 398 60914 582 61098 0 FreeSans 800 270 0 0 VDDR
port 37 nsew
flabel metal2 186 60915 370 61099 0 FreeSans 800 270 0 0 VSSR
port 38 nsew
flabel metal2 72601 30885 72665 30965 0 FreeSans 1600 0 0 0 VIP
port 39 nsew
flabel metal2 72599 29870 72663 29950 0 FreeSans 1600 0 0 0 VIN
port 40 nsew
flabel metal1 -10784 61566 -10764 61590 0 FreeSans 400 0 0 0 CLKS
port 42 nsew
flabel metal1 -10778 61426 -10758 61450 0 FreeSans 400 0 0 0 CLKSB
port 43 nsew
<< end >>
