magic
tech sky130A
magscale 1 2
timestamp 1730796434
<< error_s >>
rect 3259 3932 3659 4100
rect 2118 3549 2142 3804
rect 2146 3521 2170 3776
rect 3519 3700 3659 3932
rect 3827 4060 4227 4100
rect 3827 3932 4187 4060
rect 4188 4019 4227 4060
rect 3827 3700 3967 3932
rect 2706 3580 2758 3632
rect 2700 3574 2764 3580
rect 2706 3568 2712 3574
rect 2752 3568 2758 3574
rect 2783 3570 2786 3628
rect 1621 3091 1633 3143
rect 1649 3081 1661 3133
rect 3259 3100 3659 3268
rect 2138 2989 2190 3012
rect 2110 2961 2218 2984
rect 1071 2802 1093 2910
rect 1099 2830 1121 2882
rect 3259 2879 3427 3100
rect 3519 2868 3659 3100
rect 3827 3100 4227 3268
rect 3827 2868 3967 3100
rect 2201 2729 2212 2781
rect 2229 2701 2240 2809
rect 2002 1786 2013 1894
rect 2030 1814 2041 1866
rect 275 1495 415 1727
rect 15 1327 415 1495
rect 583 1495 723 1727
rect 815 1495 983 1716
rect 3121 1713 3143 1765
rect 3149 1685 3171 1793
rect 2024 1611 2132 1634
rect 2052 1583 2104 1606
rect 583 1327 983 1495
rect 2581 1462 2593 1514
rect 2609 1452 2621 1504
rect 1456 967 1459 1025
rect 1484 1021 1490 1027
rect 1530 1021 1536 1027
rect 1478 1015 1542 1021
rect 1484 963 1536 1015
rect 275 663 415 895
rect 15 535 54 576
rect 55 535 415 663
rect 15 495 415 535
rect 583 663 723 895
rect 2072 819 2096 1074
rect 2100 791 2124 1046
rect 583 495 983 663
<< metal1 >>
rect 987 4973 993 5025
rect 1045 4973 4599 5025
rect 4651 4973 4657 5025
rect 352 4767 360 4923
rect 516 4768 4341 4923
rect 4496 4768 4502 4923
rect 516 4767 4267 4768
rect -343 4719 -291 4725
rect -291 4667 3097 4719
rect 3149 4667 3159 4719
rect -343 4661 -291 4667
rect 360 3191 516 3197
rect 516 3035 950 3191
rect 360 3029 516 3035
rect -193 2916 -37 2922
rect -37 2760 924 2916
rect -193 2754 -37 2760
rect 3318 1679 3694 1835
rect 3849 1679 3855 1835
rect 3319 1404 4342 1560
rect 4497 1404 4503 1560
rect 4599 -21 4651 -15
rect -349 -73 -343 -21
rect -291 -73 1093 -21
rect 1145 -73 1151 -21
rect 3190 -73 3196 -21
rect 3248 -73 4599 -21
rect 4599 -79 4651 -73
rect -199 -419 -193 -263
rect -37 -264 3855 -263
rect -37 -419 3694 -264
rect 3849 -419 3855 -264
<< via1 >>
rect 993 4973 1045 5025
rect 4599 4973 4651 5025
rect 360 4767 516 4923
rect 4341 4768 4496 4923
rect -343 4667 -291 4719
rect 3097 4667 3149 4719
rect 360 3035 516 3191
rect -193 2760 -37 2916
rect 3694 1679 3849 1835
rect 4342 1404 4497 1560
rect -343 -73 -291 -21
rect 1093 -73 1145 -21
rect 3196 -73 3248 -21
rect 4599 -73 4651 -21
rect -193 -419 -37 -263
rect 3694 -419 3849 -264
<< metal2 >>
rect 993 5025 1045 5031
rect 360 4923 516 4929
rect -349 4667 -343 4719
rect -291 4667 -285 4719
rect -343 -21 -291 4667
rect 360 3191 516 4767
rect 993 4652 1045 4973
rect 4599 5025 4651 5031
rect 4341 4923 4496 4929
rect 3097 4719 3149 4725
rect 3097 4661 3149 4667
rect 354 3035 360 3191
rect 516 3035 522 3191
rect -199 2760 -193 2916
rect -37 2760 -31 2916
rect -343 -79 -291 -73
rect -193 -263 -37 2760
rect 3694 1835 3849 1841
rect 1093 -21 1145 119
rect 1093 -79 1145 -73
rect 3196 -21 3248 80
rect 3196 -79 3248 -73
rect -193 -425 -37 -419
rect 3694 -264 3849 1679
rect 4341 1566 4496 4768
rect 4341 1560 4497 1566
rect 4341 1407 4342 1560
rect 4342 1398 4497 1404
rect 4599 -21 4651 4973
rect 4593 -73 4599 -21
rect 4651 -73 4657 -21
rect 3694 -425 3849 -419
use sh_bsw  sh_bsw_0
timestamp 1730796434
transform -1 0 4869 0 -1 2183
box 602 -2485 4228 -5
use sh_bsw  sh_bsw_1
timestamp 1730796434
transform 1 0 -627 0 1 2412
box 602 -2485 4228 -5
<< labels >>
flabel metal1 s 2535 4844 2535 4844 0 FreeSans 3200 0 0 0 VDDA
port 1 nsew
flabel metal1 s 3949 4996 3949 4996 0 FreeSans 1600 0 0 0 CLKS
port 2 nsew
flabel metal1 s -39 4690 -39 4690 0 FreeSans 1600 0 0 0 CLKSB
port 3 nsew
flabel metal2 s 2582 4568 2582 4568 0 FreeSans 1600 0 0 0 VIP
port 4 nsew
flabel metal2 s 1663 -6 1663 -6 0 FreeSans 1600 0 0 0 VIN
port 5 nsew
flabel metal1 s 1662 -349 1662 -349 0 FreeSans 1600 0 0 0 VSSA
port 6 nsew
flabel metal2 s 2466 4359 2466 4359 0 FreeSans 1600 0 0 0 VCP
port 7 nsew
flabel metal2 s 1777 231 1777 231 0 FreeSans 1600 0 0 0 VCN
port 8 nsew
<< end >>
