magic
tech sky130A
magscale 1 2
timestamp 1727241376
<< nwell >>
rect 53 790 6794 1312
<< pwell >>
rect 54 212 6795 734
<< metal1 >>
rect 53 1236 6794 1312
rect 244 902 254 962
rect 314 902 324 962
rect 1937 902 1947 962
rect 2007 902 2017 962
rect 3629 902 3639 962
rect 3699 902 3709 962
rect 5321 902 5331 962
rect 5391 902 5401 962
rect 792 724 802 784
rect 862 724 872 784
rect 1639 723 1649 783
rect 1709 723 1719 783
rect 2486 724 2496 784
rect 2556 724 2566 784
rect 3332 724 3342 784
rect 3402 724 3412 784
rect 4177 724 4187 784
rect 4247 724 4257 784
rect 5023 724 5033 784
rect 5093 724 5103 784
rect 5869 724 5879 784
rect 5939 724 5949 784
rect 6691 704 6790 804
rect 1152 544 1162 604
rect 1222 544 1232 604
rect 2844 544 2854 604
rect 2914 544 2924 604
rect 4536 544 4546 604
rect 4606 544 4616 604
rect 6228 544 6238 604
rect 6298 544 6308 604
rect 54 212 6795 288
<< via1 >>
rect 254 902 314 962
rect 1947 902 2007 962
rect 3639 902 3699 962
rect 5331 902 5391 962
rect 802 724 862 784
rect 1649 723 1709 783
rect 2496 724 2556 784
rect 3342 724 3402 784
rect 4187 724 4247 784
rect 5033 724 5093 784
rect 5879 724 5939 784
rect 1162 544 1222 604
rect 2854 544 2914 604
rect 4546 544 4606 604
rect 6238 544 6298 604
<< metal2 >>
rect 53 962 5391 972
rect 53 902 254 962
rect 314 902 1947 962
rect 2007 902 3639 962
rect 3699 902 5331 962
rect 53 892 5391 902
rect 802 784 862 794
rect 53 694 111 744
rect 1649 783 1709 793
rect 862 724 964 744
rect 802 694 964 724
rect 2496 784 2556 794
rect 1709 723 1802 744
rect 1649 694 1802 723
rect 3342 784 3402 794
rect 2556 724 2652 744
rect 2496 694 2652 724
rect 4187 784 4247 794
rect 3402 724 3498 744
rect 3342 694 3498 724
rect 5033 784 5093 794
rect 4247 724 4343 744
rect 4187 694 4343 724
rect 5879 784 5939 794
rect 5093 724 5189 744
rect 5033 694 5189 724
rect 5939 724 6035 744
rect 5879 694 6035 724
rect 54 604 6298 614
rect 54 544 1162 604
rect 1222 544 2854 604
rect 2914 544 4546 604
rect 4606 544 6238 604
rect 54 535 6298 544
rect 1162 534 6298 535
use epc_delay  x1
timestamp 1727241002
transform 1 0 106 0 1 784
box -53 -572 766 528
use epc_delay  x2
timestamp 1727241002
transform 1 0 953 0 1 784
box -53 -572 766 528
use epc_delay  x3
timestamp 1727241002
transform 1 0 1799 0 1 784
box -53 -572 766 528
use epc_delay  x4
timestamp 1727241002
transform 1 0 2645 0 1 784
box -53 -572 766 528
use epc_delay  x5
timestamp 1727241002
transform 1 0 3491 0 1 784
box -53 -572 766 528
use epc_delay  x6
timestamp 1727241002
transform 1 0 4337 0 1 784
box -53 -572 766 528
use epc_delay  x7
timestamp 1727241002
transform 1 0 5183 0 1 784
box -53 -572 766 528
use epc_delay  x8
timestamp 1727241002
transform 1 0 6029 0 1 784
box -53 -572 766 528
<< labels >>
flabel metal1 86 1274 94 1278 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal2 86 928 94 932 0 FreeSans 320 0 0 0 VP
port 1 nsew
flabel metal2 76 716 84 720 0 FreeSans 320 0 0 0 IN
port 2 nsew
flabel metal2 80 572 88 576 0 FreeSans 320 0 0 0 VN
port 3 nsew
flabel metal1 84 244 92 248 0 FreeSans 320 0 0 0 VSS
port 4 nsew
flabel metal1 6750 756 6758 760 0 FreeSans 320 0 0 0 OUT
port 6 nsew
<< end >>
