magic
tech sky130A
magscale 1 2
timestamp 1730796434
<< error_s >>
rect 2629 -626 2640 -518
rect 2657 -598 2668 -546
rect 902 -917 1042 -685
rect 642 -1085 1042 -917
rect 1210 -917 1350 -685
rect 1442 -917 1610 -696
rect 3748 -699 3770 -647
rect 3776 -727 3798 -619
rect 2651 -801 2759 -778
rect 2679 -829 2731 -806
rect 1210 -1085 1610 -917
rect 3208 -950 3220 -898
rect 3236 -960 3248 -908
rect 2083 -1445 2086 -1387
rect 2111 -1391 2117 -1385
rect 2157 -1391 2163 -1385
rect 2105 -1397 2169 -1391
rect 2111 -1449 2163 -1397
rect 902 -1749 1042 -1517
rect 642 -1877 681 -1836
rect 682 -1877 1042 -1749
rect 642 -1917 1042 -1877
rect 1210 -1749 1350 -1517
rect 2699 -1593 2723 -1338
rect 2727 -1621 2751 -1366
rect 1210 -1917 1610 -1749
<< nwell >>
rect 2591 -842 2637 -679
rect 3846 -1344 4198 -1232
rect 3894 -1578 3930 -1522
rect 3894 -1612 3952 -1578
<< pwell >>
rect 1727 -989 1795 -981
rect 2679 -989 2731 -981
rect 1727 -1041 2083 -989
rect 2679 -1041 2737 -989
rect 1727 -1049 1795 -1041
rect 1922 -1074 2000 -1041
rect 2679 -1047 2731 -1041
rect 1720 -1095 1772 -1089
rect 1714 -1147 1778 -1095
rect 1917 -1147 1981 -1095
rect 1720 -1153 1772 -1147
rect 1923 -1153 1975 -1147
rect 1837 -1223 1988 -1177
rect 2031 -1221 2083 -1142
rect 3162 -1470 3214 -1468
rect 3130 -1481 3220 -1470
rect 3130 -1482 3499 -1481
rect 3130 -1522 3526 -1482
rect 3130 -1568 3499 -1522
rect 3846 -1957 4112 -1706
<< nsubdiff >>
rect 3928 -1302 3952 -1268
rect 4086 -1302 4110 -1268
<< nsubdiffcont >>
rect 3952 -1302 4086 -1268
<< locali >>
rect 3928 -1302 3952 -1268
rect 4086 -1302 4110 -1268
<< viali >>
rect 3788 -727 3822 -583
rect 3952 -1302 4086 -1268
rect 3956 -1688 3990 -1654
rect 4059 -1688 4093 -1654
<< metal1 >>
rect 2061 -481 2284 -429
rect 2336 -481 2342 -429
rect 3776 -583 4101 -577
rect 2591 -808 2637 -679
rect 3776 -727 3788 -583
rect 3822 -727 4101 -583
rect 3776 -733 4101 -727
rect 2140 -842 2637 -808
rect 2679 -812 2731 -806
rect 2679 -870 2731 -864
rect 2278 -950 2284 -898
rect 2336 -950 3125 -898
rect 3214 -950 3220 -898
rect 3817 -909 4102 -852
rect 3480 -956 4102 -909
rect 1729 -1041 1735 -989
rect 1787 -1041 2679 -989
rect 2731 -1041 3350 -989
rect 3480 -996 3823 -956
rect 3817 -1008 3823 -996
rect 3875 -1008 4102 -956
rect 1714 -1147 1720 -1095
rect 1772 -1101 1778 -1095
rect 1917 -1101 1923 -1095
rect 1772 -1147 1923 -1101
rect 1975 -1147 1981 -1095
rect 1094 -1221 1100 -1169
rect 1152 -1175 1158 -1169
rect 2031 -1175 2083 -1142
rect 1152 -1221 2083 -1175
rect 3823 -1268 4160 -1254
rect 3823 -1302 3952 -1268
rect 4086 -1302 4160 -1268
rect 3823 -1352 4160 -1302
rect 3875 -1404 4160 -1352
rect 3823 -1413 4160 -1404
rect 2111 -1449 2163 -1443
rect 3130 -1556 3136 -1470
rect 3214 -1481 3220 -1470
rect 3214 -1556 3526 -1481
rect 3130 -1568 3526 -1556
rect 3817 -1698 3823 -1646
rect 3875 -1654 4014 -1646
rect 3875 -1688 3956 -1654
rect 3990 -1688 4014 -1654
rect 3875 -1698 4014 -1688
rect 4047 -1654 4170 -1646
rect 4047 -1688 4059 -1654
rect 4093 -1688 4170 -1654
rect 4047 -1698 4170 -1688
rect 4222 -1698 4228 -1646
rect 942 -2005 948 -1953
rect 1000 -2005 3242 -1953
rect 3294 -2005 3300 -1953
rect 1509 -2085 1515 -2033
rect 1567 -2085 3712 -2033
rect 3764 -2085 3770 -2033
rect 679 -2165 685 -2113
rect 737 -2165 1720 -2113
rect 1772 -2165 2958 -2113
rect 3010 -2165 3016 -2113
rect 1247 -2245 1253 -2193
rect 1305 -2245 3823 -2193
rect 3875 -2245 3881 -2193
rect 3032 -2325 3038 -2273
rect 3090 -2325 4170 -2273
rect 4222 -2325 4228 -2273
rect 2721 -2405 2727 -2353
rect 2779 -2405 3903 -2353
rect 3955 -2405 3961 -2353
<< via1 >>
rect 2284 -481 2336 -429
rect 2679 -864 2731 -812
rect 2284 -950 2336 -898
rect 3125 -950 3214 -898
rect 1735 -1041 1787 -989
rect 2679 -1041 2731 -989
rect 3823 -1008 3875 -956
rect 1720 -1147 1772 -1095
rect 1923 -1147 1975 -1095
rect 1100 -1221 1152 -1169
rect 2111 -1443 2163 -1391
rect 3823 -1404 3875 -1352
rect 3136 -1556 3214 -1470
rect 3823 -1698 3875 -1646
rect 4170 -1698 4222 -1646
rect 3903 -1935 3955 -1883
rect 948 -2005 1000 -1953
rect 3242 -2005 3294 -1953
rect 1515 -2085 1567 -2033
rect 3712 -2085 3764 -2033
rect 685 -2165 737 -2113
rect 1720 -2165 1772 -2113
rect 2958 -2165 3010 -2113
rect 1253 -2245 1305 -2193
rect 3823 -2245 3875 -2193
rect 3038 -2325 3090 -2273
rect 4170 -2325 4222 -2273
rect 2727 -2405 2779 -2353
rect 3903 -2405 3955 -2353
<< metal2 >>
rect 2284 -429 2336 -423
rect 1733 -987 1789 -977
rect 1967 -1022 2019 -665
rect 1098 -1058 1154 -1049
rect 1733 -1052 1789 -1043
rect 1923 -1074 2019 -1022
rect 1098 -1123 1154 -1114
rect 1720 -1095 1772 -1089
rect 1100 -1169 1152 -1123
rect 1100 -1227 1152 -1221
rect 948 -1953 1000 -1947
rect 948 -2026 1000 -2005
rect 945 -2035 1001 -2026
rect 945 -2100 1001 -2091
rect 1513 -2033 1569 -2027
rect 1513 -2037 1515 -2033
rect 1567 -2037 1569 -2033
rect 683 -2109 739 -2100
rect 1513 -2102 1569 -2093
rect 683 -2174 739 -2165
rect 1720 -2113 1772 -1147
rect 1923 -1095 1975 -1074
rect 2198 -1147 2250 -751
rect 2284 -898 2336 -481
rect 2657 -598 3090 -546
rect 2284 -956 2336 -950
rect 2679 -812 2731 -806
rect 2679 -989 2731 -864
rect 2679 -1047 2731 -1041
rect 1923 -1153 1975 -1147
rect 2111 -1199 2250 -1147
rect 2111 -1391 2163 -1199
rect 2111 -1449 2163 -1443
rect 1251 -2191 1307 -2182
rect 1251 -2256 1307 -2247
rect 1720 -2485 1772 -2165
rect 2261 -2485 2313 -1473
rect 2379 -2485 2431 -1448
rect 2727 -2353 2779 -1366
rect 3038 -1574 3090 -598
rect 3125 -898 3214 -892
rect 3125 -1470 3214 -950
rect 3823 -956 3875 -950
rect 3823 -1352 3875 -1008
rect 3823 -1413 3875 -1404
rect 3125 -1556 3136 -1470
rect 3125 -1568 3214 -1556
rect 2958 -2113 3010 -1583
rect 3823 -1646 3875 -1640
rect 2958 -2171 3010 -2165
rect 3038 -2273 3090 -1703
rect 3242 -1953 3294 -1707
rect 3242 -2011 3294 -2005
rect 3712 -2033 3764 -1720
rect 3712 -2091 3764 -2085
rect 3038 -2331 3090 -2325
rect 3823 -2193 3875 -1698
rect 4170 -1646 4222 -1640
rect 2727 -2411 2779 -2405
rect 3823 -2485 3875 -2245
rect 3903 -1883 3955 -1877
rect 3903 -2353 3955 -1935
rect 4170 -2273 4222 -1698
rect 4170 -2331 4222 -2325
rect 3903 -2411 3955 -2405
<< via2 >>
rect 1733 -989 1789 -987
rect 1733 -1041 1735 -989
rect 1735 -1041 1787 -989
rect 1787 -1041 1789 -989
rect 1733 -1043 1789 -1041
rect 1098 -1114 1154 -1058
rect 945 -2091 1001 -2035
rect 1513 -2085 1515 -2037
rect 1515 -2085 1567 -2037
rect 1567 -2085 1569 -2037
rect 1513 -2093 1569 -2085
rect 683 -2113 739 -2109
rect 683 -2165 685 -2113
rect 685 -2165 737 -2113
rect 737 -2165 739 -2113
rect 1251 -2193 1307 -2191
rect 1251 -2245 1253 -2193
rect 1253 -2245 1305 -2193
rect 1305 -2245 1307 -2193
rect 1251 -2247 1307 -2245
<< metal3 >>
rect 1710 -983 1810 -964
rect 1710 -1047 1729 -983
rect 1793 -1047 1810 -983
rect 1082 -1058 1170 -1049
rect 1082 -1114 1098 -1058
rect 1154 -1114 1170 -1058
rect 1710 -1064 1810 -1047
rect 1082 -1125 1170 -1114
rect 681 -2104 741 -1956
rect 923 -2031 1023 -2017
rect 923 -2095 941 -2031
rect 1005 -2095 1023 -2031
rect 678 -2109 744 -2104
rect 678 -2165 683 -2109
rect 739 -2165 744 -2109
rect 923 -2117 1023 -2095
rect 678 -2174 744 -2165
rect 1249 -2174 1309 -1945
rect 1490 -2033 1590 -2017
rect 1490 -2097 1509 -2033
rect 1573 -2097 1590 -2033
rect 1490 -2117 1590 -2097
rect 1246 -2191 1312 -2174
rect 1246 -2247 1251 -2191
rect 1307 -2247 1312 -2191
rect 1246 -2256 1312 -2247
<< via3 >>
rect 1729 -987 1793 -983
rect 1729 -1043 1733 -987
rect 1733 -1043 1789 -987
rect 1789 -1043 1793 -987
rect 1729 -1047 1793 -1043
rect 941 -2035 1005 -2031
rect 941 -2091 945 -2035
rect 945 -2091 1001 -2035
rect 1001 -2091 1005 -2035
rect 941 -2095 1005 -2091
rect 1509 -2037 1573 -2033
rect 1509 -2093 1513 -2037
rect 1513 -2093 1569 -2037
rect 1569 -2093 1573 -2037
rect 1509 -2097 1573 -2093
<< metal4 >>
rect 1727 -983 1795 -981
rect 1727 -985 1729 -983
rect 1256 -1045 1729 -985
rect 1727 -1047 1729 -1045
rect 1793 -1047 1795 -983
rect 1727 -1049 1795 -1047
rect 943 -1994 1003 -1861
rect 941 -2030 1005 -1994
rect 940 -2031 1006 -2030
rect 940 -2095 941 -2031
rect 1005 -2095 1006 -2031
rect 1511 -2032 1571 -1870
rect 940 -2096 1006 -2095
rect 1508 -2033 1574 -2032
rect 1508 -2097 1509 -2033
rect 1573 -2097 1574 -2033
rect 1508 -2098 1574 -2097
use cap_bsw  cap_bsw_1
timestamp 1730796434
transform 0 -1 516 1 0 -3419
box 1462 -1134 3066 -86
use ncell_bsw  ncell_bsw_1
timestamp 1730778869
transform 1 0 -1493 0 1 -281
box 4653 -1676 5339 -261
use ncell_bsw_dischrg  ncell_bsw_dischrg_1
timestamp 1730741927
transform -1 0 2198 0 -1 -1730
box -138 -1725 548 -824
use ncell_bsw_sw  ncell_bsw_sw_1
timestamp 1730741762
transform -1 0 2593 0 -1 -4705
box -503 -3662 879 -2886
use pcell_bsw_dischrg  pcell_bsw_dischrg_1
timestamp 1730722715
transform 1 0 1748 0 1 -420
box 611 -449 1297 145
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform 1 0 3884 0 1 -1909
box -38 -48 314 592
<< labels >>
flabel metal1 s 4102 -926 4102 -926 0 FreeSans 480 0 0 0 VDDA
port 1 nsew
flabel metal2 s 3850 -2485 3850 -2485 0 FreeSans 480 0 0 0 CLKS
port 2 nsew
flabel metal2 s 1746 -2485 1746 -2485 0 FreeSans 480 0 0 0 CLKSB
port 3 nsew
flabel metal2 s 2287 -2485 2287 -2485 0 FreeSans 480 0 0 0 VI
port 4 nsew
flabel metal1 s 4101 -656 4101 -656 0 FreeSans 480 0 0 0 VSSA
port 5 nsew
flabel metal2 s 2405 -2485 2405 -2485 0 FreeSans 480 0 0 0 VO
port 6 nsew
<< end >>
