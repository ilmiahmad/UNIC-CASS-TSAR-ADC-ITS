* PEX produced on Sel 12 Nov 2024 06:37:25  CST using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from nooverlap_clk.ext - technology: sky130A

.subckt nooverlap_clk vdda in vssa clk0 clkb0 clk1 clkb1
X0 x2.B.t0 in.t0 vdda.t40 vdda.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1 clkb1.t15 x9.Y.t8 vssa.t33 vssa.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 clkb1.t7 x9.Y.t9 vdda.t17 vdda.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 vdda.t30 x2.A.t2 x8.Y.t3 vdda.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 clk0.t7 clkb0.t16 vdda.t52 vdda.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 clk0.t6 clkb0.t17 vdda.t47 vdda.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 vssa.t45 x8.Y.t8 clkb0.t15 vssa.t44 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 clkb1.t14 x9.Y.t10 vssa.t31 vssa.t30 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 clkb1.t6 x9.Y.t11 vdda.t16 vdda.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 vdda.t56 x2.A.t3 x8.Y.t2 vdda.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 vssa.t67 clkb0.t18 clk0.t15 vssa.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 clkb0.t7 x8.Y.t9 vdda.t50 vdda.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 x2.Y.t0 x2.A.t4 a_n135_n688.t0 vssa.t63 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 clk0.t5 clkb0.t19 vdda.t9 vdda.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 clkb0.t14 x8.Y.t10 vssa.t39 vssa.t38 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 vdda.t37 x2.A.t5 x2.Y.t1 vdda.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 x9.Y.t1 x1.B.t2 vssa.t13 vssa.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 x9.Y.t3 x1.B.t3 vdda.t49 vdda.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 vssa.t58 clkb1.t16 clk1.t15 vssa.t57 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 x1.B.t0 x5.Y.t2 vssa.t15 vssa.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X20 clkb0.t6 x8.Y.t11 vdda.t32 vdda.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 vdda.t43 clkb1.t17 clk1.t7 vdda.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X22 x1.B.t1 x5.Y.t3 vdda.t68 vdda.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X23 clk0.t14 clkb0.t20 vssa.t71 vssa.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 x9.Y.t7 x1.B.t4 vssa.t85 vssa.t84 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X25 x9.Y.t2 x1.B.t5 vdda.t33 vdda.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 vssa.t41 x8.Y.t12 clkb0.t13 vssa.t40 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 vssa.t73 clkb1.t18 clk1.t14 vssa.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 vdda.t58 clkb1.t19 clk1.t6 vdda.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 clkb0.t5 x8.Y.t13 vdda.t3 vdda.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 vssa.t47 clkb0.t21 clk0.t13 vssa.t46 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 x1.Y.t1 in.t1 a_n135_176.t0 vssa.t50 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 x5.Y.t1 x2.Y.t3 vssa.t62 vssa.t61 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X33 x5.Y.t0 x2.Y.t4 vdda.t62 vdda.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X34 clkb0.t12 x8.Y.t14 vssa.t65 vssa.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X35 vssa.t29 x9.Y.t12 clkb1.t13 vssa.t28 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 vssa.t87 clkb1.t20 clk1.t13 vssa.t86 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 vdda.t14 x9.Y.t13 clkb1.t5 vdda.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 vdda.t42 clkb1.t21 clk1.t5 vdda.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 clkb0.t4 x8.Y.t15 vdda.t73 vdda.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X40 a_n135_176.t1 x1.B.t6 vssa.t69 vssa.t68 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X41 vdda.t38 in.t2 x1.Y.t0 vdda.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 clk0.t12 clkb0.t22 vssa.t37 vssa.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X43 vssa.t27 x9.Y.t14 clkb1.t12 vssa.t26 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X44 vssa.t79 clkb1.t22 clk1.t12 vssa.t78 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X45 vdda.t60 x9.Y.t15 clkb1.t4 vdda.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X46 x8.Y.t1 x2.A.t6 vdda.t64 vdda.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X47 vssa.t43 x8.Y.t16 clkb0.t11 vssa.t42 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X48 vssa.t75 x2.A.t7 x8.Y.t7 vssa.t74 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 vssa.t25 x9.Y.t16 clkb1.t11 vssa.t24 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X50 vdda.t24 clkb1.t23 clk1.t4 vdda.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X51 vdda.t35 x9.Y.t17 clkb1.t3 vdda.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X52 x2.A.t0 x4.Y.t2 vssa.t17 vssa.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X53 vdda.t13 clkb0.t23 clk0.t4 vdda.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X54 x2.A.t1 x4.Y.t3 vdda.t70 vdda.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X55 vssa.t9 clkb0.t24 clk0.t11 vssa.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X56 x8.Y.t0 x2.A.t8 vdda.t1 vdda.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X57 vssa.t23 x9.Y.t18 clkb1.t10 vssa.t22 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X58 vdda.t20 x9.Y.t19 clkb1.t2 vdda.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 clkb0.t10 x8.Y.t17 vssa.t91 vssa.t90 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X60 x8.Y.t6 x2.A.t9 vssa.t5 vssa.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X61 vdda.t45 clkb0.t25 clk0.t3 vdda.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X62 x4.Y.t1 x1.Y.t3 vssa.t93 vssa.t92 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X63 x4.Y.t0 x1.Y.t4 vdda.t69 vdda.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X64 vdda.t7 x8.Y.t18 clkb0.t3 vdda.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X65 vssa.t7 x8.Y.t19 clkb0.t9 vssa.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X66 vssa.t3 x2.A.t10 x8.Y.t5 vssa.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X67 vdda.t55 clkb0.t26 clk0.t2 vdda.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X68 a_n135_n688.t1 x2.B.t2 vssa.t77 vssa.t76 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X69 x2.Y.t2 x2.B.t3 vdda.t22 vdda.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X70 clk1.t11 clkb1.t24 vssa.t56 vssa.t55 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X71 vdda.t71 x8.Y.t20 clkb0.t2 vdda.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X72 clk1.t3 clkb1.t25 vdda.t66 vdda.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X73 vdda.t51 clkb0.t27 clk0.t1 vdda.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X74 vssa.t11 clkb0.t28 clk0.t10 vssa.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X75 vdda.t72 x8.Y.t21 clkb0.t1 vdda.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X76 clkb0.t8 x8.Y.t22 vssa.t89 vssa.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X77 x8.Y.t4 x2.A.t11 vssa.t95 vssa.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X78 vssa.t83 x1.B.t7 x9.Y.t6 vssa.t82 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X79 clk1.t10 clkb1.t26 vssa.t1 vssa.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X80 clk1.t9 clkb1.t27 vssa.t52 vssa.t51 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X81 clk1.t2 clkb1.t28 vdda.t57 vdda.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X82 vdda.t53 x1.B.t8 x9.Y.t4 vdda.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X83 clk1.t1 clkb1.t29 vdda.t26 vdda.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X84 clk0.t9 clkb0.t29 vssa.t35 vssa.t34 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X85 vdda.t5 x8.Y.t23 clkb0.t0 vdda.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X86 clk0.t8 clkb0.t30 vssa.t60 vssa.t59 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X87 vssa.t81 x1.B.t9 x9.Y.t5 vssa.t80 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X88 clkb1.t9 x9.Y.t20 vssa.t21 vssa.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X89 vdda.t11 x1.B.t10 x9.Y.t0 vdda.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X90 clk1.t8 clkb1.t30 vssa.t54 vssa.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X91 clkb1.t1 x9.Y.t21 vdda.t19 vdda.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X92 clk1.t0 clkb1.t31 vdda.t65 vdda.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X93 x1.Y.t2 x1.B.t11 vdda.t54 vdda.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X94 clkb1.t8 x9.Y.t22 vssa.t19 vssa.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X95 clkb1.t0 x9.Y.t23 vdda.t63 vdda.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X96 clk0.t0 clkb0.t31 vdda.t28 vdda.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X97 x2.B.t1 in.t3 vssa.t49 vssa.t48 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 in.n0 in.t0 230.576
R1 in.n1 in.t2 230.155
R2 in.n0 in.t3 158.275
R3 in.n1 in.t1 157.856
R4 in.n4 in.n0 154.133
R5 in.n2 in.n1 153.147
R6 in.n4 in.n3 25.0079
R7 in.n3 in.n2 13.9592
R8 in in.n4 4.53383
R9 in.n2 in 3.24826
R10 in.n3 in 0.513893
R11 vdda.n20 vdda.t30 877.144
R12 vdda.n20 vdda.t53 877.144
R13 vdda.n12 vdda.n11 402
R14 vdda.n52 vdda.t57 342.377
R15 vdda.n70 vdda.t16 342.377
R16 vdda.n52 vdda.t47 342.375
R17 vdda.n70 vdda.t73 342.375
R18 vdda.n37 vdda.t43 338.892
R19 vdda.n57 vdda.t35 338.892
R20 vdda.n37 vdda.t13 338.892
R21 vdda.n57 vdda.t72 338.892
R22 vdda.n76 vdda.n18 320.976
R23 vdda.n41 vdda.n40 320.976
R24 vdda.n44 vdda.n43 320.976
R25 vdda.n50 vdda.n35 320.976
R26 vdda.n30 vdda.n29 320.976
R27 vdda.n63 vdda.n27 320.976
R28 vdda.n24 vdda.n23 320.976
R29 vdda.n76 vdda.n19 320.976
R30 vdda.n41 vdda.n39 320.976
R31 vdda.n44 vdda.n42 320.976
R32 vdda.n50 vdda.n34 320.976
R33 vdda.n30 vdda.n28 320.976
R34 vdda.n63 vdda.n26 320.976
R35 vdda.n24 vdda.n22 320.976
R36 vdda.t67 vdda 285.337
R37 vdda vdda.t39 283.658
R38 vdda.n2 vdda.t62 255.905
R39 vdda.n83 vdda.t68 255.905
R40 vdda.n2 vdda.t69 255.904
R41 vdda.n83 vdda.t70 255.904
R42 vdda.n11 vdda.t40 254.475
R43 vdda.n92 vdda.t37 249.363
R44 vdda.n92 vdda.t38 249.362
R45 vdda.n16 vdda.t33 248.843
R46 vdda.n16 vdda.t1 248.843
R47 vdda.n6 vdda.t22 247.394
R48 vdda.n6 vdda.t54 247.394
R49 vdda.t34 vdda 238.339
R50 vdda.n13 vdda.t61 231.625
R51 vdda.t29 vdda 223.233
R52 vdda vdda.t36 206.45
R53 vdda vdda.t67 177.916
R54 vdda.t61 vdda 177.916
R55 vdda vdda.t46 164.488
R56 vdda vdda.t15 164.488
R57 vdda.t8 vdda.t12 140.989
R58 vdda.t44 vdda.t8 140.989
R59 vdda.t27 vdda.t44 140.989
R60 vdda.t41 vdda.t27 140.989
R61 vdda.t25 vdda.t41 140.989
R62 vdda.t23 vdda.t25 140.989
R63 vdda.t46 vdda.t23 140.989
R64 vdda.t18 vdda.t34 140.989
R65 vdda.t4 vdda.t18 140.989
R66 vdda.t31 vdda.t4 140.989
R67 vdda.t6 vdda.t31 140.989
R68 vdda.t2 vdda.t6 140.989
R69 vdda.t59 vdda.t2 140.989
R70 vdda.t15 vdda.t59 140.989
R71 vdda.t48 vdda.t29 140.989
R72 vdda.t10 vdda.t48 140.989
R73 vdda.t0 vdda.t10 140.989
R74 vdda.t36 vdda.t21 140.989
R75 vdda vdda.t0 125.883
R76 vdda.t21 vdda 117.492
R77 vdda.n12 vdda 105.743
R78 vdda.t39 vdda.n12 72.1736
R79 vdda.n13 vdda 53.7107
R80 vdda.n14 vdda.n13 52.8576
R81 vdda.n10 vdda.n5 34.6358
R82 vdda.n49 vdda.n36 34.6358
R83 vdda.n53 vdda.n51 34.6358
R84 vdda.n59 vdda.n58 34.6358
R85 vdda.n65 vdda.n64 34.6358
R86 vdda.n69 vdda.n68 34.6358
R87 vdda.n76 vdda.n75 34.6358
R88 vdda.n77 vdda.n76 34.6358
R89 vdda.n82 vdda.n81 34.6358
R90 vdda.n88 vdda.n87 34.6358
R91 vdda.n45 vdda.n44 32.0005
R92 vdda.n63 vdda.n62 32.0005
R93 vdda.n45 vdda.n41 31.2476
R94 vdda.n62 vdda.n30 31.2476
R95 vdda.n71 vdda.n20 31.2476
R96 vdda.n57 vdda.n32 27.8593
R97 vdda.n81 vdda.n16 27.1064
R98 vdda.n19 vdda.t64 26.5955
R99 vdda.n19 vdda.t56 26.5955
R100 vdda.n18 vdda.t49 26.5955
R101 vdda.n18 vdda.t11 26.5955
R102 vdda.n40 vdda.t65 26.5955
R103 vdda.n40 vdda.t58 26.5955
R104 vdda.n39 vdda.t9 26.5955
R105 vdda.n39 vdda.t45 26.5955
R106 vdda.n43 vdda.t66 26.5955
R107 vdda.n43 vdda.t42 26.5955
R108 vdda.n42 vdda.t28 26.5955
R109 vdda.n42 vdda.t55 26.5955
R110 vdda.n35 vdda.t26 26.5955
R111 vdda.n35 vdda.t24 26.5955
R112 vdda.n34 vdda.t52 26.5955
R113 vdda.n34 vdda.t51 26.5955
R114 vdda.n29 vdda.t19 26.5955
R115 vdda.n29 vdda.t20 26.5955
R116 vdda.n28 vdda.t50 26.5955
R117 vdda.n28 vdda.t5 26.5955
R118 vdda.n27 vdda.t63 26.5955
R119 vdda.n27 vdda.t14 26.5955
R120 vdda.n26 vdda.t32 26.5955
R121 vdda.n26 vdda.t7 26.5955
R122 vdda.n23 vdda.t17 26.5955
R123 vdda.n23 vdda.t60 26.5955
R124 vdda.n22 vdda.t3 26.5955
R125 vdda.n22 vdda.t71 26.5955
R126 vdda.n92 vdda.n1 25.977
R127 vdda.n50 vdda.n49 25.977
R128 vdda.n65 vdda.n24 25.977
R129 vdda.n6 vdda.n1 24.4711
R130 vdda.n6 vdda.n5 23.7181
R131 vdda.n92 vdda.n91 23.7181
R132 vdda.n75 vdda.n20 22.2123
R133 vdda.n77 vdda.n16 22.2123
R134 vdda.n58 vdda.n57 18.824
R135 vdda.n84 vdda.n14 18.4476
R136 vdda.n87 vdda.n14 16.1887
R137 vdda.n11 vdda.n4 15.7005
R138 vdda.n53 vdda.n52 13.5534
R139 vdda.n70 vdda.n69 13.5534
R140 vdda.n41 vdda.n38 10.5481
R141 vdda.n83 vdda.n82 10.5417
R142 vdda.n88 vdda.n2 10.5417
R143 vdda.n85 vdda.n84 9.3005
R144 vdda.n46 vdda.n45 9.3005
R145 vdda.n47 vdda.n36 9.3005
R146 vdda.n49 vdda.n48 9.3005
R147 vdda.n51 vdda.n33 9.3005
R148 vdda.n54 vdda.n53 9.3005
R149 vdda.n55 vdda.n32 9.3005
R150 vdda.n57 vdda.n56 9.3005
R151 vdda.n58 vdda.n31 9.3005
R152 vdda.n60 vdda.n59 9.3005
R153 vdda.n62 vdda.n61 9.3005
R154 vdda.n64 vdda.n25 9.3005
R155 vdda.n66 vdda.n65 9.3005
R156 vdda.n68 vdda.n67 9.3005
R157 vdda.n69 vdda.n21 9.3005
R158 vdda.n72 vdda.n71 9.3005
R159 vdda.n73 vdda.n20 9.3005
R160 vdda.n75 vdda.n74 9.3005
R161 vdda.n76 vdda.n17 9.3005
R162 vdda.n78 vdda.n77 9.3005
R163 vdda.n79 vdda.n16 9.3005
R164 vdda.n81 vdda.n80 9.3005
R165 vdda.n82 vdda.n15 9.3005
R166 vdda.n10 vdda.n9 9.3005
R167 vdda.n8 vdda.n5 9.3005
R168 vdda.n7 vdda.n6 9.3005
R169 vdda.n87 vdda.n86 9.3005
R170 vdda.n89 vdda.n88 9.3005
R171 vdda.n91 vdda.n90 9.3005
R172 vdda.n93 vdda.n92 9.3005
R173 vdda.n1 vdda.n0 9.3005
R174 vdda.n51 vdda.n50 8.65932
R175 vdda.n68 vdda.n24 8.65932
R176 vdda.n91 vdda.n2 8.28285
R177 vdda.n84 vdda.n83 8.28285
R178 vdda.n38 vdda.n37 6.6132
R179 vdda.n11 vdda.n10 6.4005
R180 vdda.n3 vdda 5.14243
R181 vdda.n59 vdda.n30 3.38874
R182 vdda.n44 vdda.n36 2.63579
R183 vdda.n64 vdda.n63 2.63579
R184 vdda.n52 vdda.n32 1.88285
R185 vdda.n71 vdda.n70 1.88285
R186 vdda.n46 vdda.n38 0.567773
R187 vdda.n47 vdda.n46 0.120292
R188 vdda.n48 vdda.n47 0.120292
R189 vdda.n48 vdda.n33 0.120292
R190 vdda.n54 vdda.n33 0.120292
R191 vdda.n55 vdda.n54 0.120292
R192 vdda.n56 vdda.n31 0.120292
R193 vdda.n60 vdda.n31 0.120292
R194 vdda.n61 vdda.n60 0.120292
R195 vdda.n61 vdda.n25 0.120292
R196 vdda.n66 vdda.n25 0.120292
R197 vdda.n67 vdda.n66 0.120292
R198 vdda.n67 vdda.n21 0.120292
R199 vdda.n72 vdda.n21 0.120292
R200 vdda.n74 vdda.n73 0.120292
R201 vdda.n74 vdda.n17 0.120292
R202 vdda.n78 vdda.n17 0.120292
R203 vdda.n79 vdda.n78 0.120292
R204 vdda.n80 vdda.n15 0.120292
R205 vdda.n85 vdda.n15 0.120292
R206 vdda.n90 vdda.n89 0.120292
R207 vdda.n93 vdda.n0 0.120292
R208 vdda.n7 vdda.n0 0.120292
R209 vdda.n9 vdda.n8 0.120292
R210 vdda.n9 vdda.n4 0.120292
R211 vdda.n89 vdda.n3 0.0838333
R212 vdda.n56 vdda 0.0603958
R213 vdda.n73 vdda 0.0603958
R214 vdda.n80 vdda 0.0603958
R215 vdda.n86 vdda 0.0603958
R216 vdda vdda.n93 0.0603958
R217 vdda.n8 vdda 0.0603958
R218 vdda.n86 vdda.n3 0.0369583
R219 vdda vdda.n7 0.0239375
R220 vdda vdda.n55 0.0226354
R221 vdda vdda.n72 0.0226354
R222 vdda vdda.n79 0.0226354
R223 vdda vdda.n85 0.0226354
R224 vdda.n90 vdda 0.0226354
R225 vdda.n4 vdda 0.0226354
R226 x2.B.n3 x2.B.t0 235.56
R227 x2.B.n0 x2.B.t3 229.369
R228 x2.B.n0 x2.B.t2 157.07
R229 x2.B.n1 x2.B.n0 153.897
R230 x2.B x2.B.t1 152.889
R231 x2.B.n2 x2.B.n1 18.937
R232 x2.B x2.B.n2 14.1918
R233 x2.B.n2 x2.B 4.73093
R234 x2.B.n1 x2.B 4.03013
R235 x2.B.n3 x2.B 2.22659
R236 x2.B x2.B.n3 1.55202
R237 x9.Y.n8 x9.Y.n7 244.069
R238 x9.Y.n5 x9.Y.n3 236.589
R239 x9.Y.n13 x9.Y.t17 212.081
R240 x9.Y.n12 x9.Y.t21 212.081
R241 x9.Y.n17 x9.Y.t19 212.081
R242 x9.Y.n19 x9.Y.t23 212.081
R243 x9.Y.n10 x9.Y.t13 212.081
R244 x9.Y.n25 x9.Y.t9 212.081
R245 x9.Y.n27 x9.Y.t15 212.081
R246 x9.Y.n28 x9.Y.t11 212.081
R247 x9.Y.n8 x9.Y.n6 204.893
R248 x9.Y.n5 x9.Y.n4 200.321
R249 x9.Y x9.Y.n29 163.264
R250 x9.Y.n26 x9.Y.n9 152
R251 x9.Y.n24 x9.Y.n23 152
R252 x9.Y.n18 x9.Y.n11 152
R253 x9.Y.n2 x9.Y.n20 152
R254 x9.Y.n16 x9.Y.n15 152
R255 x9.Y x9.Y.n14 152
R256 x9.Y.n13 x9.Y.t16 139.78
R257 x9.Y.n12 x9.Y.t20 139.78
R258 x9.Y.n17 x9.Y.t18 139.78
R259 x9.Y.n19 x9.Y.t22 139.78
R260 x9.Y.n10 x9.Y.t12 139.78
R261 x9.Y.n25 x9.Y.t8 139.78
R262 x9.Y.n27 x9.Y.t14 139.78
R263 x9.Y.n28 x9.Y.t10 139.78
R264 x9.Y.n14 x9.Y.n13 30.6732
R265 x9.Y.n14 x9.Y.n12 30.6732
R266 x9.Y.n16 x9.Y.n12 30.6732
R267 x9.Y.n17 x9.Y.n16 30.6732
R268 x9.Y.n20 x9.Y.n17 30.6732
R269 x9.Y.n20 x9.Y.n19 30.6732
R270 x9.Y.n19 x9.Y.n18 30.6732
R271 x9.Y.n18 x9.Y.n10 30.6732
R272 x9.Y.n24 x9.Y.n10 30.6732
R273 x9.Y.n25 x9.Y.n24 30.6732
R274 x9.Y.n26 x9.Y.n25 30.6732
R275 x9.Y.n27 x9.Y.n26 30.6732
R276 x9.Y.n29 x9.Y.n27 30.6732
R277 x9.Y.n29 x9.Y.n28 30.6732
R278 x9.Y.n6 x9.Y.t4 26.5955
R279 x9.Y.n6 x9.Y.t3 26.5955
R280 x9.Y.n7 x9.Y.t0 26.5955
R281 x9.Y.n7 x9.Y.t2 26.5955
R282 x9.Y.n3 x9.Y.t5 24.9236
R283 x9.Y.n3 x9.Y.t7 24.9236
R284 x9.Y.n4 x9.Y.t6 24.9236
R285 x9.Y.n4 x9.Y.t1 24.9236
R286 x9.Y.n15 x9.Y.n1 6.51899
R287 x9.Y.n2 x9.Y 19.2005
R288 x9.Y x9.Y.n8 18.4569
R289 x9.Y x9.Y.n11 17.4085
R290 x9.Y.n23 x9.Y 15.3605
R291 x9.Y.n32 x9.Y 14.008
R292 x9.Y x9.Y.n1 6.28716
R293 x9.Y x9.Y.n9 13.3125
R294 x9.Y.n31 x9.Y 12.3175
R295 x9.Y.n32 x9.Y.n5 12.0894
R296 x9.Y.n31 x9.Y.n0 9.96396
R297 x9.Y.n0 x9.Y.n30 9.3005
R298 x9.Y.n22 x9.Y.n0 9.3005
R299 x9.Y.n21 x9.Y.n0 9.3005
R300 x9.Y.n0 x9.Y.n2 9.3005
R301 x9.Y.n30 x9.Y.n9 5.8885
R302 x9.Y x9.Y.n21 4.3525
R303 x9.Y.n22 x9.Y 4.3525
R304 x9.Y.n30 x9.Y 4.3525
R305 x9.Y.n2 x9.Y 4.3525
R306 x9.Y x9.Y.n31 4.10616
R307 x9.Y.n1 x9.Y.n0 3.93048
R308 x9.Y.n23 x9.Y.n22 3.8405
R309 x9.Y x9.Y.n32 2.41559
R310 x9.Y.n15 x9.Y 2.0485
R311 x9.Y.n21 x9.Y.n11 1.7925
R312 vssa vssa.t16 2420.71
R313 vssa vssa.t92 2420.71
R314 vssa vssa.t14 2420.71
R315 vssa vssa.t61 2420.71
R316 vssa vssa.t48 2406.47
R317 vssa.t42 vssa 2022.01
R318 vssa.t24 vssa 2022.01
R319 vssa vssa.t74 1893.85
R320 vssa vssa.t82 1893.85
R321 vssa vssa.t50 1751.46
R322 vssa vssa.t63 1751.46
R323 vssa.t16 vssa 1509.39
R324 vssa.t92 vssa 1509.39
R325 vssa.t14 vssa 1509.39
R326 vssa.t61 vssa 1509.39
R327 vssa.t48 vssa 1509.39
R328 vssa vssa.t59 1395.47
R329 vssa vssa.t51 1395.47
R330 vssa.t34 vssa.t10 1196.12
R331 vssa.t66 vssa.t34 1196.12
R332 vssa.t70 vssa.t66 1196.12
R333 vssa.t46 vssa.t70 1196.12
R334 vssa.t36 vssa.t46 1196.12
R335 vssa.t8 vssa.t36 1196.12
R336 vssa.t59 vssa.t8 1196.12
R337 vssa.t90 vssa.t42 1196.12
R338 vssa.t6 vssa.t90 1196.12
R339 vssa.t88 vssa.t6 1196.12
R340 vssa.t44 vssa.t88 1196.12
R341 vssa.t38 vssa.t44 1196.12
R342 vssa.t40 vssa.t38 1196.12
R343 vssa.t64 vssa.t40 1196.12
R344 vssa.t74 vssa.t4 1196.12
R345 vssa.t4 vssa.t2 1196.12
R346 vssa.t2 vssa.t94 1196.12
R347 vssa.t50 vssa.t68 1196.12
R348 vssa.t53 vssa.t57 1196.12
R349 vssa.t72 vssa.t53 1196.12
R350 vssa.t55 vssa.t72 1196.12
R351 vssa.t86 vssa.t55 1196.12
R352 vssa.t0 vssa.t86 1196.12
R353 vssa.t78 vssa.t0 1196.12
R354 vssa.t51 vssa.t78 1196.12
R355 vssa.t20 vssa.t24 1196.12
R356 vssa.t22 vssa.t20 1196.12
R357 vssa.t18 vssa.t22 1196.12
R358 vssa.t28 vssa.t18 1196.12
R359 vssa.t32 vssa.t28 1196.12
R360 vssa.t26 vssa.t32 1196.12
R361 vssa.t30 vssa.t26 1196.12
R362 vssa.t82 vssa.t12 1196.12
R363 vssa.t12 vssa.t80 1196.12
R364 vssa.t80 vssa.t84 1196.12
R365 vssa.t63 vssa.t76 1196.12
R366 vssa.n10 vssa.t64 1153.4
R367 vssa.n93 vssa.t30 1153.4
R368 vssa.t94 vssa 1067.96
R369 vssa.t84 vssa 1067.96
R370 vssa.t68 vssa 996.764
R371 vssa.t76 vssa 996.764
R372 vssa.n24 vssa.t11 289.87
R373 vssa.n107 vssa.t58 289.87
R374 vssa.n37 vssa.t43 284.024
R375 vssa.n120 vssa.t25 284.024
R376 vssa.n9 vssa.t65 282.885
R377 vssa.n34 vssa.t60 282.885
R378 vssa.n117 vssa.t52 282.885
R379 vssa.n92 vssa.t31 282.885
R380 vssa.n5 vssa.t95 282.327
R381 vssa.n88 vssa.t85 282.327
R382 vssa.n8 vssa.t75 281.13
R383 vssa.n91 vssa.t83 281.13
R384 vssa.n10 vssa 242.071
R385 vssa.n93 vssa 242.071
R386 vssa.n60 vssa.n7 207.213
R387 vssa.n50 vssa.n12 207.213
R388 vssa.n44 vssa.n43 207.213
R389 vssa.n42 vssa.n15 207.213
R390 vssa.n19 vssa.n18 207.213
R391 vssa.n27 vssa.n21 207.213
R392 vssa.n23 vssa.n22 207.213
R393 vssa.n143 vssa.n90 207.213
R394 vssa.n106 vssa.n105 207.213
R395 vssa.n110 vssa.n104 207.213
R396 vssa.n102 vssa.n101 207.213
R397 vssa.n125 vssa.n98 207.213
R398 vssa.n127 vssa.n126 207.213
R399 vssa.n133 vssa.n95 207.213
R400 vssa.n71 vssa.t93 153.631
R401 vssa.n3 vssa.t17 153.631
R402 vssa.n86 vssa.t15 153.631
R403 vssa.n84 vssa.t62 153.631
R404 vssa.n165 vssa.t49 153.631
R405 vssa.n78 vssa.t69 150.922
R406 vssa.n162 vssa.t77 150.922
R407 vssa.n7 vssa.t5 24.9236
R408 vssa.n7 vssa.t3 24.9236
R409 vssa.n12 vssa.t39 24.9236
R410 vssa.n12 vssa.t41 24.9236
R411 vssa.n43 vssa.t89 24.9236
R412 vssa.n43 vssa.t45 24.9236
R413 vssa.n15 vssa.t91 24.9236
R414 vssa.n15 vssa.t7 24.9236
R415 vssa.n18 vssa.t37 24.9236
R416 vssa.n18 vssa.t9 24.9236
R417 vssa.n21 vssa.t71 24.9236
R418 vssa.n21 vssa.t47 24.9236
R419 vssa.n22 vssa.t35 24.9236
R420 vssa.n22 vssa.t67 24.9236
R421 vssa.n90 vssa.t13 24.9236
R422 vssa.n90 vssa.t81 24.9236
R423 vssa.n105 vssa.t54 24.9236
R424 vssa.n105 vssa.t73 24.9236
R425 vssa.n104 vssa.t56 24.9236
R426 vssa.n104 vssa.t87 24.9236
R427 vssa.n101 vssa.t1 24.9236
R428 vssa.n101 vssa.t79 24.9236
R429 vssa.n98 vssa.t21 24.9236
R430 vssa.n98 vssa.t23 24.9236
R431 vssa.n126 vssa.t19 24.9236
R432 vssa.n126 vssa.t29 24.9236
R433 vssa.n95 vssa.t33 24.9236
R434 vssa.n95 vssa.t27 24.9236
R435 vssa.n55 vssa.n10 24.8941
R436 vssa.n138 vssa.n93 24.8941
R437 vssa.n41 vssa.n40 20.3039
R438 vssa.n49 vssa.n13 20.3039
R439 vssa.n52 vssa.n51 20.3039
R440 vssa.n56 vssa.n55 20.3039
R441 vssa.n60 vssa.n59 20.3039
R442 vssa.n61 vssa.n60 20.3039
R443 vssa.n65 vssa.n64 20.3039
R444 vssa.n66 vssa.n65 20.3039
R445 vssa.n70 vssa.n69 20.3039
R446 vssa.n72 vssa.n70 20.3039
R447 vssa.n76 vssa.n1 20.3039
R448 vssa.n77 vssa.n76 20.3039
R449 vssa.n29 vssa.n28 20.3039
R450 vssa.n33 vssa.n32 20.3039
R451 vssa.n112 vssa.n111 20.3039
R452 vssa.n116 vssa.n115 20.3039
R453 vssa.n124 vssa.n123 20.3039
R454 vssa.n132 vssa.n96 20.3039
R455 vssa.n135 vssa.n134 20.3039
R456 vssa.n139 vssa.n138 20.3039
R457 vssa.n143 vssa.n142 20.3039
R458 vssa.n144 vssa.n143 20.3039
R459 vssa.n148 vssa.n147 20.3039
R460 vssa.n149 vssa.n148 20.3039
R461 vssa.n153 vssa.n152 20.3039
R462 vssa.n154 vssa.n153 20.3039
R463 vssa.n158 vssa.n157 20.3039
R464 vssa.n158 vssa.n83 20.3039
R465 vssa.n167 vssa.n166 20.3039
R466 vssa.n61 vssa.n5 18.9798
R467 vssa.n144 vssa.n88 18.9798
R468 vssa.n45 vssa.n44 18.7591
R469 vssa.n27 vssa.n26 18.7591
R470 vssa.n110 vssa.n109 18.7591
R471 vssa.n128 vssa.n127 18.7591
R472 vssa.n59 vssa.n8 18.5384
R473 vssa.n142 vssa.n91 18.5384
R474 vssa.n165 vssa.n164 18.3488
R475 vssa.n45 vssa.n42 18.3177
R476 vssa.n26 vssa.n23 18.3177
R477 vssa.n109 vssa.n106 18.3177
R478 vssa.n128 vssa.n125 18.3177
R479 vssa.n35 vssa.n16 16.1108
R480 vssa.n118 vssa.n99 16.1108
R481 vssa.n78 vssa.n77 15.4986
R482 vssa.n50 vssa.n49 15.2281
R483 vssa.n29 vssa.n19 15.2281
R484 vssa.n112 vssa.n102 15.2281
R485 vssa.n133 vssa.n132 15.2281
R486 vssa.n167 vssa.n163 13.9039
R487 vssa.n52 vssa.n9 13.6833
R488 vssa.n34 vssa.n33 13.6833
R489 vssa.n117 vssa.n116 13.6833
R490 vssa.n135 vssa.n92 13.6833
R491 vssa.n163 vssa.n83 13.0212
R492 vssa.n66 vssa.n3 11.2557
R493 vssa.n72 vssa.n71 11.2557
R494 vssa.n149 vssa.n86 11.2557
R495 vssa.n154 vssa.n84 11.2557
R496 vssa.n166 vssa.n165 11.2557
R497 vssa.n40 vssa.n16 11.035
R498 vssa.n123 vssa.n99 11.035
R499 vssa.n26 vssa.n25 9.3005
R500 vssa.n28 vssa.n20 9.3005
R501 vssa.n30 vssa.n29 9.3005
R502 vssa.n32 vssa.n31 9.3005
R503 vssa.n33 vssa.n17 9.3005
R504 vssa.n36 vssa.n35 9.3005
R505 vssa.n38 vssa.n37 9.3005
R506 vssa.n40 vssa.n39 9.3005
R507 vssa.n41 vssa.n14 9.3005
R508 vssa.n46 vssa.n45 9.3005
R509 vssa.n47 vssa.n13 9.3005
R510 vssa.n49 vssa.n48 9.3005
R511 vssa.n51 vssa.n11 9.3005
R512 vssa.n53 vssa.n52 9.3005
R513 vssa.n55 vssa.n54 9.3005
R514 vssa.n57 vssa.n56 9.3005
R515 vssa.n59 vssa.n58 9.3005
R516 vssa.n60 vssa.n6 9.3005
R517 vssa.n62 vssa.n61 9.3005
R518 vssa.n64 vssa.n63 9.3005
R519 vssa.n65 vssa.n4 9.3005
R520 vssa.n67 vssa.n66 9.3005
R521 vssa.n69 vssa.n68 9.3005
R522 vssa.n70 vssa.n2 9.3005
R523 vssa.n73 vssa.n72 9.3005
R524 vssa.n74 vssa.n1 9.3005
R525 vssa.n76 vssa.n75 9.3005
R526 vssa.n77 vssa.n0 9.3005
R527 vssa.n79 vssa.n78 9.3005
R528 vssa.n109 vssa.n108 9.3005
R529 vssa.n111 vssa.n103 9.3005
R530 vssa.n113 vssa.n112 9.3005
R531 vssa.n115 vssa.n114 9.3005
R532 vssa.n116 vssa.n100 9.3005
R533 vssa.n119 vssa.n118 9.3005
R534 vssa.n121 vssa.n120 9.3005
R535 vssa.n123 vssa.n122 9.3005
R536 vssa.n124 vssa.n97 9.3005
R537 vssa.n129 vssa.n128 9.3005
R538 vssa.n130 vssa.n96 9.3005
R539 vssa.n132 vssa.n131 9.3005
R540 vssa.n134 vssa.n94 9.3005
R541 vssa.n136 vssa.n135 9.3005
R542 vssa.n138 vssa.n137 9.3005
R543 vssa.n140 vssa.n139 9.3005
R544 vssa.n142 vssa.n141 9.3005
R545 vssa.n143 vssa.n89 9.3005
R546 vssa.n145 vssa.n144 9.3005
R547 vssa.n147 vssa.n146 9.3005
R548 vssa.n148 vssa.n87 9.3005
R549 vssa.n150 vssa.n149 9.3005
R550 vssa.n152 vssa.n151 9.3005
R551 vssa.n153 vssa.n85 9.3005
R552 vssa.n155 vssa.n154 9.3005
R553 vssa.n157 vssa.n156 9.3005
R554 vssa.n159 vssa.n158 9.3005
R555 vssa.n160 vssa.n83 9.3005
R556 vssa.n162 vssa.n161 9.3005
R557 vssa.n168 vssa.n167 9.3005
R558 vssa.n166 vssa.n82 9.3005
R559 vssa.n69 vssa.n3 9.04877
R560 vssa.n71 vssa.n1 9.04877
R561 vssa.n152 vssa.n86 9.04877
R562 vssa.n157 vssa.n84 9.04877
R563 vssa.n24 vssa.n23 8.18207
R564 vssa.n107 vssa.n106 8.18207
R565 vssa.n55 vssa.n9 6.62119
R566 vssa.n35 vssa.n34 6.62119
R567 vssa.n118 vssa.n117 6.62119
R568 vssa.n138 vssa.n92 6.62119
R569 vssa.n81 vssa 5.85076
R570 vssa.n51 vssa.n50 5.07636
R571 vssa.n32 vssa.n19 5.07636
R572 vssa.n115 vssa.n102 5.07636
R573 vssa.n134 vssa.n133 5.07636
R574 vssa vssa.n80 4.55909
R575 vssa.n37 vssa.n16 2.51853
R576 vssa.n120 vssa.n99 2.51853
R577 vssa.n163 vssa.n162 2.47792
R578 vssa.n42 vssa.n41 1.98671
R579 vssa.n125 vssa.n124 1.98671
R580 vssa.n56 vssa.n8 1.76602
R581 vssa.n139 vssa.n91 1.76602
R582 vssa.n44 vssa.n13 1.54533
R583 vssa.n28 vssa.n27 1.54533
R584 vssa.n111 vssa.n110 1.54533
R585 vssa.n127 vssa.n96 1.54533
R586 vssa.n64 vssa.n5 1.32464
R587 vssa.n147 vssa.n88 1.32464
R588 vssa.n25 vssa.n24 0.846184
R589 vssa.n108 vssa.n107 0.846184
R590 vssa.n25 vssa.n20 0.120292
R591 vssa.n30 vssa.n20 0.120292
R592 vssa.n31 vssa.n30 0.120292
R593 vssa.n31 vssa.n17 0.120292
R594 vssa.n36 vssa.n17 0.120292
R595 vssa.n39 vssa.n38 0.120292
R596 vssa.n39 vssa.n14 0.120292
R597 vssa.n46 vssa.n14 0.120292
R598 vssa.n47 vssa.n46 0.120292
R599 vssa.n48 vssa.n47 0.120292
R600 vssa.n48 vssa.n11 0.120292
R601 vssa.n53 vssa.n11 0.120292
R602 vssa.n54 vssa.n53 0.120292
R603 vssa.n58 vssa.n57 0.120292
R604 vssa.n58 vssa.n6 0.120292
R605 vssa.n62 vssa.n6 0.120292
R606 vssa.n63 vssa.n62 0.120292
R607 vssa.n67 vssa.n4 0.120292
R608 vssa.n68 vssa.n67 0.120292
R609 vssa.n73 vssa.n2 0.120292
R610 vssa.n74 vssa.n73 0.120292
R611 vssa.n75 vssa.n0 0.120292
R612 vssa.n79 vssa.n0 0.120292
R613 vssa.n108 vssa.n103 0.120292
R614 vssa.n113 vssa.n103 0.120292
R615 vssa.n114 vssa.n113 0.120292
R616 vssa.n114 vssa.n100 0.120292
R617 vssa.n119 vssa.n100 0.120292
R618 vssa.n122 vssa.n121 0.120292
R619 vssa.n122 vssa.n97 0.120292
R620 vssa.n129 vssa.n97 0.120292
R621 vssa.n130 vssa.n129 0.120292
R622 vssa.n131 vssa.n130 0.120292
R623 vssa.n131 vssa.n94 0.120292
R624 vssa.n136 vssa.n94 0.120292
R625 vssa.n137 vssa.n136 0.120292
R626 vssa.n141 vssa.n140 0.120292
R627 vssa.n141 vssa.n89 0.120292
R628 vssa.n145 vssa.n89 0.120292
R629 vssa.n146 vssa.n145 0.120292
R630 vssa.n150 vssa.n87 0.120292
R631 vssa.n151 vssa.n150 0.120292
R632 vssa.n155 vssa.n85 0.120292
R633 vssa.n156 vssa.n155 0.120292
R634 vssa.n160 vssa.n159 0.120292
R635 vssa.n161 vssa.n160 0.120292
R636 vssa.n168 vssa.n82 0.120292
R637 vssa.n164 vssa.n82 0.120292
R638 vssa.n38 vssa 0.0603958
R639 vssa.n57 vssa 0.0603958
R640 vssa vssa.n4 0.0603958
R641 vssa vssa.n2 0.0603958
R642 vssa.n75 vssa 0.0603958
R643 vssa.n121 vssa 0.0603958
R644 vssa.n140 vssa 0.0603958
R645 vssa vssa.n87 0.0603958
R646 vssa vssa.n85 0.0603958
R647 vssa.n159 vssa 0.0603958
R648 vssa vssa.n168 0.0603958
R649 vssa vssa.n36 0.0226354
R650 vssa.n54 vssa 0.0226354
R651 vssa.n63 vssa 0.0226354
R652 vssa.n68 vssa 0.0226354
R653 vssa vssa.n74 0.0226354
R654 vssa vssa.n119 0.0226354
R655 vssa.n137 vssa 0.0226354
R656 vssa.n146 vssa 0.0226354
R657 vssa.n151 vssa 0.0226354
R658 vssa.n156 vssa 0.0226354
R659 vssa.n164 vssa 0.0226354
R660 vssa.n80 vssa 0.0174271
R661 vssa vssa.n81 0.0174271
R662 vssa.n80 vssa.n79 0.00701042
R663 vssa.n161 vssa.n81 0.00701042
R664 clkb1.n2 clkb1.t17 212.081
R665 clkb1.n46 clkb1.t31 212.081
R666 clkb1.n3 clkb1.t19 212.081
R667 clkb1.n9 clkb1.t25 212.081
R668 clkb1.n11 clkb1.t21 212.081
R669 clkb1.n37 clkb1.t29 212.081
R670 clkb1.n12 clkb1.t23 212.081
R671 clkb1.n13 clkb1.t28 212.081
R672 clkb1.n26 clkb1.n21 205.28
R673 clkb1.n25 clkb1.n22 205.28
R674 clkb1.n24 clkb1.n23 205.28
R675 clkb1.n16 clkb1.n15 205.28
R676 clkb1 clkb1.n14 163.264
R677 clkb1.n36 clkb1.n35 152
R678 clkb1.n39 clkb1.n38 152
R679 clkb1.n10 clkb1.n6 152
R680 clkb1.n8 clkb1.n4 152
R681 clkb1.n45 clkb1.n44 152
R682 clkb1 clkb1.n47 152
R683 clkb1.n2 clkb1.t16 139.78
R684 clkb1.n46 clkb1.t30 139.78
R685 clkb1.n3 clkb1.t18 139.78
R686 clkb1.n9 clkb1.t24 139.78
R687 clkb1.n11 clkb1.t20 139.78
R688 clkb1.n37 clkb1.t26 139.78
R689 clkb1.n12 clkb1.t22 139.78
R690 clkb1.n13 clkb1.t27 139.78
R691 clkb1.n30 clkb1.n17 99.1759
R692 clkb1.n29 clkb1.n18 99.1759
R693 clkb1.n28 clkb1.n19 99.1759
R694 clkb1.n27 clkb1.n20 99.1759
R695 clkb1.n26 clkb1.n25 38.4005
R696 clkb1.n25 clkb1.n24 38.4005
R697 clkb1.n24 clkb1.n16 38.4005
R698 clkb1 clkb1.n26 36.4472
R699 clkb1.n30 clkb1.n29 34.3584
R700 clkb1.n29 clkb1.n28 34.3584
R701 clkb1.n28 clkb1.n27 34.3584
R702 clkb1.n31 clkb1.n16 31.0358
R703 clkb1.n47 clkb1.n2 30.6732
R704 clkb1.n47 clkb1.n46 30.6732
R705 clkb1.n46 clkb1.n45 30.6732
R706 clkb1.n45 clkb1.n3 30.6732
R707 clkb1.n8 clkb1.n3 30.6732
R708 clkb1.n9 clkb1.n8 30.6732
R709 clkb1.n10 clkb1.n9 30.6732
R710 clkb1.n11 clkb1.n10 30.6732
R711 clkb1.n38 clkb1.n11 30.6732
R712 clkb1.n38 clkb1.n37 30.6732
R713 clkb1.n37 clkb1.n36 30.6732
R714 clkb1.n36 clkb1.n12 30.6732
R715 clkb1.n14 clkb1.n12 30.6732
R716 clkb1.n14 clkb1.n13 30.6732
R717 clkb1.n27 clkb1 27.7875
R718 clkb1.n21 clkb1.t4 26.5955
R719 clkb1.n21 clkb1.t6 26.5955
R720 clkb1.n22 clkb1.t5 26.5955
R721 clkb1.n22 clkb1.t7 26.5955
R722 clkb1.n23 clkb1.t2 26.5955
R723 clkb1.n23 clkb1.t0 26.5955
R724 clkb1.n15 clkb1.t3 26.5955
R725 clkb1.n15 clkb1.t1 26.5955
R726 clkb1 clkb1.n30 25.611
R727 clkb1.n17 clkb1.t11 24.9236
R728 clkb1.n17 clkb1.t9 24.9236
R729 clkb1.n18 clkb1.t10 24.9236
R730 clkb1.n18 clkb1.t8 24.9236
R731 clkb1.n19 clkb1.t13 24.9236
R732 clkb1.n19 clkb1.t15 24.9236
R733 clkb1.n20 clkb1.t12 24.9236
R734 clkb1.n20 clkb1.t14 24.9236
R735 clkb1 clkb1.n1 19.2005
R736 clkb1 clkb1.n43 19.2005
R737 clkb1.n6 clkb1 17.4085
R738 clkb1 clkb1.n39 15.3605
R739 clkb1 clkb1.n0 13.8737
R740 clkb1.n35 clkb1 13.3125
R741 clkb1.n34 clkb1.n33 9.3005
R742 clkb1.n7 clkb1.n5 9.3005
R743 clkb1.n41 clkb1.n40 9.3005
R744 clkb1.n43 clkb1.n42 9.3005
R745 clkb1.n1 clkb1.n0 9.3005
R746 clkb1.n32 clkb1.n31 9.3005
R747 clkb1.n32 clkb1 7.09614
R748 clkb1.n35 clkb1.n34 5.8885
R749 clkb1.n40 clkb1 4.3525
R750 clkb1 clkb1.n7 4.3525
R751 clkb1.n34 clkb1 4.3525
R752 clkb1 clkb1.n4 4.0965
R753 clkb1.n39 clkb1.n7 3.8405
R754 clkb1.n31 clkb1 3.4005
R755 clkb1.n44 clkb1.n1 2.3045
R756 clkb1.n44 clkb1 2.0485
R757 clkb1.n40 clkb1.n6 1.7925
R758 clkb1.n33 clkb1.n32 0.663962
R759 clkb1.n43 clkb1.n4 0.2565
R760 clkb1.n42 clkb1.n0 0.221654
R761 clkb1.n42 clkb1.n41 0.221654
R762 clkb1.n41 clkb1.n5 0.221654
R763 clkb1.n33 clkb1.n5 0.221654
R764 x2.A x2.A.t1 230.518
R765 x2.A.n14 x2.A.t5 230.155
R766 x2.A.n3 x2.A.t2 212.081
R767 x2.A.n4 x2.A.t6 212.081
R768 x2.A.n1 x2.A.t3 212.081
R769 x2.A.n11 x2.A.t8 212.081
R770 x2.A.n12 x2.A.n11 188.516
R771 x2.A.n14 x2.A.t4 157.856
R772 x2.A.n16 x2.A.t0 157.62
R773 x2.A.n10 x2.A.n9 152
R774 x2.A.n7 x2.A.n2 152
R775 x2.A.n6 x2.A.n5 152
R776 x2.A.n15 x2.A.n14 152
R777 x2.A.n3 x2.A.t7 139.78
R778 x2.A.n4 x2.A.t9 139.78
R779 x2.A.n1 x2.A.t10 139.78
R780 x2.A.n11 x2.A.t11 139.78
R781 x2.A.n5 x2.A.n3 30.6732
R782 x2.A.n5 x2.A.n4 30.6732
R783 x2.A.n4 x2.A.n2 30.6732
R784 x2.A.n2 x2.A.n1 30.6732
R785 x2.A.n10 x2.A.n1 30.6732
R786 x2.A.n11 x2.A.n10 30.6732
R787 x2.A.n0 x2.A.n15 22.8779
R788 x2.A.n7 x2.A 19.2005
R789 x2.A.n9 x2.A 17.1525
R790 x2.A.n12 x2.A 17.1525
R791 x2.A.n17 x2.A 11.6875
R792 x2.A.n0 x2.A.n6 11.5697
R793 x2.A.n7 x2.A.n0 10.0818
R794 x2.A.n8 x2.A.n0 9.3005
R795 x2.A.n0 x2.A.n13 9.3005
R796 x2.A.n16 x2.A.n0 9.3005
R797 x2.A.n17 x2.A 7.23528
R798 x2.A x2.A.n17 5.04292
R799 x2.A x2.A.n16 4.73093
R800 x2.A x2.A.n7 4.3525
R801 x2.A.n8 x2.A 4.3525
R802 x2.A.n13 x2.A 4.3525
R803 x2.A.n6 x2.A 2.3045
R804 x2.A.n15 x2.A 2.3045
R805 x2.A.n9 x2.A.n8 2.0485
R806 x2.A.n13 x2.A.n12 2.0485
R807 x8.Y.n32 x8.Y.n30 244.069
R808 x8.Y.n5 x8.Y.n3 236.589
R809 x8.Y.n10 x8.Y.t21 212.081
R810 x8.Y.n12 x8.Y.t9 212.081
R811 x8.Y.n15 x8.Y.t23 212.081
R812 x8.Y.n17 x8.Y.t11 212.081
R813 x8.Y.n7 x8.Y.t18 212.081
R814 x8.Y.n23 x8.Y.t13 212.081
R815 x8.Y.n25 x8.Y.t20 212.081
R816 x8.Y.n26 x8.Y.t15 212.081
R817 x8.Y.n32 x8.Y.n31 204.893
R818 x8.Y.n5 x8.Y.n4 200.321
R819 x8.Y x8.Y.n27 163.264
R820 x8.Y.n24 x8.Y.n6 152
R821 x8.Y.n22 x8.Y.n21 152
R822 x8.Y.n16 x8.Y.n8 152
R823 x8.Y.n0 x8.Y.n18 152
R824 x8.Y.n14 x8.Y.n13 152
R825 x8.Y.n11 x8.Y 152
R826 x8.Y.n10 x8.Y.t16 139.78
R827 x8.Y.n12 x8.Y.t17 139.78
R828 x8.Y.n15 x8.Y.t19 139.78
R829 x8.Y.n17 x8.Y.t22 139.78
R830 x8.Y.n7 x8.Y.t8 139.78
R831 x8.Y.n23 x8.Y.t10 139.78
R832 x8.Y.n25 x8.Y.t12 139.78
R833 x8.Y.n26 x8.Y.t14 139.78
R834 x8.Y.n11 x8.Y.n10 30.6732
R835 x8.Y.n12 x8.Y.n11 30.6732
R836 x8.Y.n14 x8.Y.n12 30.6732
R837 x8.Y.n15 x8.Y.n14 30.6732
R838 x8.Y.n18 x8.Y.n15 30.6732
R839 x8.Y.n18 x8.Y.n17 30.6732
R840 x8.Y.n17 x8.Y.n16 30.6732
R841 x8.Y.n16 x8.Y.n7 30.6732
R842 x8.Y.n22 x8.Y.n7 30.6732
R843 x8.Y.n23 x8.Y.n22 30.6732
R844 x8.Y.n24 x8.Y.n23 30.6732
R845 x8.Y.n25 x8.Y.n24 30.6732
R846 x8.Y.n27 x8.Y.n25 30.6732
R847 x8.Y.n27 x8.Y.n26 30.6732
R848 x8.Y.n30 x8.Y.t2 26.5955
R849 x8.Y.n30 x8.Y.t0 26.5955
R850 x8.Y.n31 x8.Y.t3 26.5955
R851 x8.Y.n31 x8.Y.t1 26.5955
R852 x8.Y.n3 x8.Y.t5 24.9236
R853 x8.Y.n3 x8.Y.t4 24.9236
R854 x8.Y.n4 x8.Y.t7 24.9236
R855 x8.Y.n4 x8.Y.t6 24.9236
R856 x8.Y.n0 x8.Y 19.2005
R857 x8.Y x8.Y.n5 17.8856
R858 x8.Y x8.Y.n8 17.4085
R859 x8.Y.n21 x8.Y 15.3605
R860 x8.Y.n33 x8.Y 15.2156
R861 x8.Y x8.Y.n6 13.3125
R862 x8.Y.n29 x8.Y 12.3175
R863 x8.Y.n33 x8.Y.n32 11.4531
R864 x8.Y.n29 x8.Y.n1 9.96396
R865 x8.Y.n20 x8.Y.n1 9.3005
R866 x8.Y.n1 x8.Y.n28 9.3005
R867 x8.Y.n2 x8.Y.n0 9.3005
R868 x8.Y.n19 x8.Y.n2 9.3005
R869 x8.Y.n13 x8.Y.n9 6.51899
R870 x8.Y x8.Y.n9 6.28716
R871 x8.Y.n28 x8.Y.n6 5.8885
R872 x8.Y x8.Y.n19 4.3525
R873 x8.Y.n20 x8.Y 4.3525
R874 x8.Y.n28 x8.Y 4.3525
R875 x8.Y.n0 x8.Y 4.3525
R876 x8.Y x8.Y.n29 4.10616
R877 x8.Y.n21 x8.Y.n20 3.8405
R878 x8.Y.n2 x8.Y.n9 3.26701
R879 x8.Y.n13 x8.Y 2.0485
R880 x8.Y.n19 x8.Y.n8 1.7925
R881 x8.Y x8.Y.n33 1.20805
R882 x8.Y.n2 x8.Y.n1 0.663962
R883 clkb0.n5 clkb0.t23 212.081
R884 clkb0.n7 clkb0.t19 212.081
R885 clkb0.n10 clkb0.t25 212.081
R886 clkb0.n12 clkb0.t31 212.081
R887 clkb0.n2 clkb0.t26 212.081
R888 clkb0.n22 clkb0.t16 212.081
R889 clkb0.n24 clkb0.t27 212.081
R890 clkb0.n25 clkb0.t17 212.081
R891 clkb0.n46 clkb0.n31 205.28
R892 clkb0.n45 clkb0.n32 205.28
R893 clkb0.n44 clkb0.n33 205.28
R894 clkb0.n43 clkb0.n34 205.28
R895 clkb0 clkb0.n26 163.264
R896 clkb0.n23 clkb0.n1 152
R897 clkb0.n21 clkb0.n20 152
R898 clkb0.n11 clkb0.n3 152
R899 clkb0.n14 clkb0.n13 152
R900 clkb0.n9 clkb0.n8 152
R901 clkb0.n6 clkb0 152
R902 clkb0.n5 clkb0.t28 139.78
R903 clkb0.n7 clkb0.t29 139.78
R904 clkb0.n10 clkb0.t18 139.78
R905 clkb0.n12 clkb0.t20 139.78
R906 clkb0.n2 clkb0.t21 139.78
R907 clkb0.n22 clkb0.t22 139.78
R908 clkb0.n24 clkb0.t24 139.78
R909 clkb0.n25 clkb0.t30 139.78
R910 clkb0.n42 clkb0.n35 99.1759
R911 clkb0.n41 clkb0.n36 99.1749
R912 clkb0.n40 clkb0.n37 99.1749
R913 clkb0.n39 clkb0.n38 99.1749
R914 clkb0.n46 clkb0.n45 38.4005
R915 clkb0.n45 clkb0.n44 38.4005
R916 clkb0.n44 clkb0.n43 38.4005
R917 clkb0.n42 clkb0.n41 34.3584
R918 clkb0.n41 clkb0.n40 34.3584
R919 clkb0.n40 clkb0.n39 34.3584
R920 clkb0 clkb0.n42 34.0948
R921 clkb0.n6 clkb0.n5 30.6732
R922 clkb0.n7 clkb0.n6 30.6732
R923 clkb0.n9 clkb0.n7 30.6732
R924 clkb0.n10 clkb0.n9 30.6732
R925 clkb0.n13 clkb0.n10 30.6732
R926 clkb0.n13 clkb0.n12 30.6732
R927 clkb0.n12 clkb0.n11 30.6732
R928 clkb0.n11 clkb0.n2 30.6732
R929 clkb0.n21 clkb0.n2 30.6732
R930 clkb0.n22 clkb0.n21 30.6732
R931 clkb0.n23 clkb0.n22 30.6732
R932 clkb0.n24 clkb0.n23 30.6732
R933 clkb0.n26 clkb0.n24 30.6732
R934 clkb0.n26 clkb0.n25 30.6732
R935 clkb0.n43 clkb0 30.14
R936 clkb0.n39 clkb0.n30 29.011
R937 clkb0 clkb0.n46 27.6358
R938 clkb0.n31 clkb0.t1 26.5955
R939 clkb0.n31 clkb0.t7 26.5955
R940 clkb0.n32 clkb0.t0 26.5955
R941 clkb0.n32 clkb0.t6 26.5955
R942 clkb0.n33 clkb0.t3 26.5955
R943 clkb0.n33 clkb0.t5 26.5955
R944 clkb0.n34 clkb0.t2 26.5955
R945 clkb0.n34 clkb0.t4 26.5955
R946 clkb0.n35 clkb0.t13 24.9236
R947 clkb0.n35 clkb0.t12 24.9236
R948 clkb0.n36 clkb0.t15 24.9236
R949 clkb0.n36 clkb0.t14 24.9236
R950 clkb0.n37 clkb0.t9 24.9236
R951 clkb0.n37 clkb0.t8 24.9236
R952 clkb0.n38 clkb0.t11 24.9236
R953 clkb0.n38 clkb0.t10 24.9236
R954 clkb0.n15 clkb0 19.2005
R955 clkb0 clkb0.n3 17.4085
R956 clkb0.n20 clkb0 15.3605
R957 clkb0 clkb0.n1 13.3125
R958 clkb0.n29 clkb0 9.76475
R959 clkb0.n30 clkb0.n29 9.3005
R960 clkb0.n19 clkb0.n0 9.3005
R961 clkb0.n28 clkb0.n27 9.3005
R962 clkb0.n16 clkb0.n15 9.3005
R963 clkb0.n18 clkb0.n17 9.3005
R964 clkb0.n8 clkb0.n4 6.51899
R965 clkb0 clkb0.n4 6.28716
R966 clkb0.n27 clkb0.n1 5.8885
R967 clkb0 clkb0.n18 4.3525
R968 clkb0.n19 clkb0 4.3525
R969 clkb0.n27 clkb0 4.3525
R970 clkb0.n14 clkb0 4.0965
R971 clkb0.n20 clkb0.n19 3.8405
R972 clkb0 clkb0.n30 3.4005
R973 clkb0.n16 clkb0.n4 3.26701
R974 clkb0.n8 clkb0 2.0485
R975 clkb0.n18 clkb0.n3 1.7925
R976 clkb0.n29 clkb0.n28 0.663962
R977 clkb0.n15 clkb0.n14 0.2565
R978 clkb0.n17 clkb0.n16 0.221654
R979 clkb0.n17 clkb0.n0 0.221654
R980 clkb0.n28 clkb0.n0 0.221654
R981 clk0.n16 clk0.n1 205.28
R982 clk0.n15 clk0.n2 205.28
R983 clk0.n14 clk0.n3 205.28
R984 clk0.n13 clk0.n4 205.28
R985 clk0.n12 clk0.n5 99.1759
R986 clk0.n11 clk0.n6 99.1749
R987 clk0.n10 clk0.n7 99.1749
R988 clk0.n9 clk0.n8 99.1749
R989 clk0.n16 clk0.n15 38.4005
R990 clk0.n15 clk0.n14 38.4005
R991 clk0.n14 clk0.n13 38.4005
R992 clk0.n12 clk0.n11 34.3584
R993 clk0.n11 clk0.n10 34.3584
R994 clk0.n10 clk0.n9 34.3584
R995 clk0 clk0.n12 34.0948
R996 clk0.n13 clk0 30.14
R997 clk0.n9 clk0.n0 29.011
R998 clk0 clk0.n16 27.6358
R999 clk0.n1 clk0.t4 26.5955
R1000 clk0.n1 clk0.t5 26.5955
R1001 clk0.n2 clk0.t3 26.5955
R1002 clk0.n2 clk0.t0 26.5955
R1003 clk0.n3 clk0.t2 26.5955
R1004 clk0.n3 clk0.t7 26.5955
R1005 clk0.n4 clk0.t1 26.5955
R1006 clk0.n4 clk0.t6 26.5955
R1007 clk0.n5 clk0.t11 24.9236
R1008 clk0.n5 clk0.t8 24.9236
R1009 clk0.n6 clk0.t13 24.9236
R1010 clk0.n6 clk0.t12 24.9236
R1011 clk0.n7 clk0.t15 24.9236
R1012 clk0.n7 clk0.t14 24.9236
R1013 clk0.n8 clk0.t10 24.9236
R1014 clk0.n8 clk0.t9 24.9236
R1015 clk0.n0 clk0 19.193
R1016 clk0 clk0.n0 3.4005
R1017 a_n135_n688.t0 a_n135_n688.t1 49.8467
R1018 x2.Y x2.Y.n2 237.577
R1019 x2.Y.n0 x2.Y.t4 230.576
R1020 x2.Y.n0 x2.Y.t3 158.275
R1021 x2.Y.n1 x2.Y.n0 154.133
R1022 x2.Y.n3 x2.Y.t0 140.53
R1023 x2.Y.n2 x2.Y.t1 26.5955
R1024 x2.Y.n2 x2.Y.t2 26.5955
R1025 x2.Y.n3 x2.Y.n1 19.413
R1026 x2.Y.n3 x2.Y 16.5652
R1027 x2.Y x2.Y.n3 9.03579
R1028 x2.Y.n1 x2.Y 4.53383
R1029 x2.Y.n3 x2.Y 1.72748
R1030 x1.B.n17 x1.B.t1 235.56
R1031 x1.B.n14 x1.B.t11 229.369
R1032 x1.B.n3 x1.B.t8 212.081
R1033 x1.B.n4 x1.B.t3 212.081
R1034 x1.B.n1 x1.B.t10 212.081
R1035 x1.B.n11 x1.B.t5 212.081
R1036 x1.B.n12 x1.B.n11 188.516
R1037 x1.B.n14 x1.B.t6 157.07
R1038 x1.B.n15 x1.B.n14 153.897
R1039 x1.B x1.B.t0 152.889
R1040 x1.B.n10 x1.B.n9 152
R1041 x1.B.n7 x1.B.n2 152
R1042 x1.B.n6 x1.B.n5 152
R1043 x1.B.n3 x1.B.t7 139.78
R1044 x1.B.n4 x1.B.t2 139.78
R1045 x1.B.n1 x1.B.t9 139.78
R1046 x1.B.n11 x1.B.t4 139.78
R1047 x1.B.n5 x1.B.n3 30.6732
R1048 x1.B.n5 x1.B.n4 30.6732
R1049 x1.B.n4 x1.B.n2 30.6732
R1050 x1.B.n2 x1.B.n1 30.6732
R1051 x1.B.n10 x1.B.n1 30.6732
R1052 x1.B.n11 x1.B.n10 30.6732
R1053 x1.B.n0 x1.B.n15 21.4741
R1054 x1.B.n7 x1.B 19.2005
R1055 x1.B.n9 x1.B 17.1525
R1056 x1.B.n12 x1.B 17.1525
R1057 x1.B x1.B.n16 14.1918
R1058 x1.B.n0 x1.B.n6 11.5697
R1059 x1.B.n0 x1.B.n13 9.87983
R1060 x1.B.n16 x1.B.n0 9.50242
R1061 x1.B.n8 x1.B.n0 9.3005
R1062 x1.B.n7 x1.B.n0 9.3005
R1063 x1.B.n16 x1.B 4.73093
R1064 x1.B x1.B.n7 4.3525
R1065 x1.B.n8 x1.B 4.3525
R1066 x1.B.n13 x1.B 4.3525
R1067 x1.B.n15 x1.B 4.03013
R1068 x1.B.n6 x1.B 2.3045
R1069 x1.B.n17 x1.B 2.22659
R1070 x1.B.n9 x1.B.n8 2.0485
R1071 x1.B.n13 x1.B.n12 2.0485
R1072 x1.B x1.B.n17 1.55202
R1073 clk1.n12 clk1.n5 205.28
R1074 clk1.n11 clk1.n6 205.28
R1075 clk1.n10 clk1.n7 205.28
R1076 clk1.n9 clk1.n8 205.28
R1077 clk1.n16 clk1.n1 99.1759
R1078 clk1.n15 clk1.n2 99.1759
R1079 clk1.n14 clk1.n3 99.1759
R1080 clk1.n13 clk1.n4 99.1759
R1081 clk1.n12 clk1.n11 38.4005
R1082 clk1.n11 clk1.n10 38.4005
R1083 clk1.n10 clk1.n9 38.4005
R1084 clk1 clk1.n12 36.4472
R1085 clk1.n16 clk1.n15 34.3584
R1086 clk1.n15 clk1.n14 34.3584
R1087 clk1.n14 clk1.n13 34.3584
R1088 clk1.n9 clk1.n0 31.0358
R1089 clk1.n13 clk1 27.7875
R1090 clk1.n5 clk1.t4 26.5955
R1091 clk1.n5 clk1.t2 26.5955
R1092 clk1.n6 clk1.t5 26.5955
R1093 clk1.n6 clk1.t1 26.5955
R1094 clk1.n7 clk1.t6 26.5955
R1095 clk1.n7 clk1.t3 26.5955
R1096 clk1.n8 clk1.t7 26.5955
R1097 clk1.n8 clk1.t0 26.5955
R1098 clk1 clk1.n16 25.611
R1099 clk1.n1 clk1.t15 24.9236
R1100 clk1.n1 clk1.t8 24.9236
R1101 clk1.n2 clk1.t14 24.9236
R1102 clk1.n2 clk1.t11 24.9236
R1103 clk1.n3 clk1.t13 24.9236
R1104 clk1.n3 clk1.t10 24.9236
R1105 clk1.n4 clk1.t12 24.9236
R1106 clk1.n4 clk1.t9 24.9236
R1107 clk1.n0 clk1 17.2663
R1108 clk1 clk1.n0 3.4005
R1109 x5.Y.n3 x5.Y.t0 235.56
R1110 x5.Y.n0 x5.Y.t3 230.576
R1111 x5.Y.n0 x5.Y.t2 158.275
R1112 x5.Y.n1 x5.Y.n0 154.133
R1113 x5.Y x5.Y.t1 152.889
R1114 x5.Y.n2 x5.Y.n1 19.0428
R1115 x5.Y x5.Y.n2 14.1918
R1116 x5.Y.n2 x5.Y 4.73093
R1117 x5.Y.n1 x5.Y 4.53383
R1118 x5.Y.n3 x5.Y 2.22659
R1119 x5.Y x5.Y.n3 1.55202
R1120 a_n135_176.t0 a_n135_176.t1 49.8467
R1121 x1.Y.t1 x1.Y.n2 270.471
R1122 x1.Y.n3 x1.Y.t1 258.846
R1123 x1.Y.n0 x1.Y.t4 230.576
R1124 x1.Y x1.Y.n4 224.776
R1125 x1.Y.n0 x1.Y.t3 158.275
R1126 x1.Y.n1 x1.Y.n0 154.133
R1127 x1.Y.n4 x1.Y.t0 26.5955
R1128 x1.Y.n4 x1.Y.t2 26.5955
R1129 x1.Y.n2 x1.Y.n1 19.413
R1130 x1.Y.n1 x1.Y 4.53383
R1131 x1.Y x1.Y.n3 3.03935
R1132 x1.Y.n3 x1.Y 2.30266
R1133 x1.Y.n2 x1.Y 1.56597
R1134 x4.Y.n0 x4.Y.t3 230.576
R1135 x4.Y x4.Y.t0 230.518
R1136 x4.Y.n0 x4.Y.t2 158.275
R1137 x4.Y.n2 x4.Y.t1 157.62
R1138 x4.Y.n1 x4.Y.n0 154.133
R1139 x4.Y.n2 x4.Y.n1 19.0428
R1140 x4.Y.n3 x4.Y 11.6875
R1141 x4.Y.n3 x4.Y 7.23528
R1142 x4.Y x4.Y.n3 5.04292
R1143 x4.Y x4.Y.n2 4.73093
R1144 x4.Y.n1 x4.Y 4.53383
C0 x1.Y in 0.265374f
C1 x1.Y x4.Y 0.110151f
C2 in x1.B 0.288243f
C3 x1.B x4.Y 0.16164f
C4 vdda in 0.516474f
C5 x8.Y x1.B 0.015359f
C6 clk1 clk0 0.089246f
C7 vdda x4.Y 0.355849f
C8 x2.A in 0.015286f
C9 x8.Y vdda 0.741788f
C10 x2.A x4.Y 0.110994f
C11 x1.Y x1.B 0.13464f
C12 x2.B in 0.109787f
C13 x8.Y x2.A 0.437305f
C14 x1.Y vdda 0.316184f
C15 vdda x1.B 0.91356f
C16 clkb0 clk1 0.096323f
C17 x8.Y clkb1 0.076744f
C18 x2.A x1.B 0.566464f
C19 x1.Y x2.Y 0.013041f
C20 x2.A vdda 0.92531f
C21 x2.B x1.B 0.013453f
C22 x5.Y x4.Y 0.013034f
C23 x2.B vdda 0.324442f
C24 clkb1 x1.B 0.036118f
C25 vdda x2.Y 0.313587f
C26 clkb1 vdda 1.45347f
C27 x2.B x2.A 0.068737f
C28 x2.A x2.Y 0.232728f
C29 x8.Y clk0 0.558033f
C30 clkb1 x2.A 0.01075f
C31 x5.Y x1.B 0.104979f
C32 x2.B x2.Y 0.061385f
C33 x8.Y x9.Y 0.102267f
C34 x5.Y vdda 0.301599f
C35 clkb0 in 0.14011f
C36 x5.Y x2.A 0.178189f
C37 vdda clk0 0.862792f
C38 clkb0 x4.Y 0.03182f
C39 clkb0 x8.Y 1.36777f
C40 x1.B x9.Y 0.483158f
C41 x5.Y x2.Y 0.110151f
C42 x2.A clk0 0.244344f
C43 vdda x9.Y 0.852035f
C44 clkb0 x1.Y 0.067171f
C45 clkb0 x1.B 0.37645f
C46 clkb1 clk0 0.068573f
C47 clkb0 vdda 2.48076f
C48 clkb1 x9.Y 1.28706f
C49 clkb0 x2.A 0.176172f
C50 clk1 vdda 1.15341f
C51 clkb0 clkb1 0.200628f
C52 clk1 clkb1 1.56148f
C53 clkb0 clk0 1.71059f
C54 clk1 vssa 0.859199f
C55 clkb1 vssa 1.68888f
C56 clk0 vssa 1.55769f
C57 clkb0 vssa 1.803912f
C58 in vssa 0.979546f
C59 vdda vssa 6.370696f
C60 x9.Y vssa 1.23543f
C61 x5.Y vssa 0.374286f
C62 x2.Y vssa 0.593192f
C63 x2.B vssa 0.448422f
C64 x8.Y vssa 1.03794f
C65 x2.A vssa 0.793322f
C66 x4.Y vssa 0.36813f
C67 x1.Y vssa 0.579104f
C68 x1.B vssa 1.02966f
C69 clkb0.n0 vssa 0.022752f
C70 clkb0.t24 vssa 0.011771f
C71 clkb0.t27 vssa 0.019975f
C72 clkb0.t22 vssa 0.011771f
C73 clkb0.t16 vssa 0.019975f
C74 clkb0.t21 vssa 0.011771f
C75 clkb0.t26 vssa 0.019975f
C76 clkb0.n2 vssa 0.028806f
C77 clkb0.t18 vssa 0.011771f
C78 clkb0.t25 vssa 0.019975f
C79 clkb0.t29 vssa 0.011771f
C80 clkb0.t19 vssa 0.019975f
C81 clkb0.t28 vssa 0.011771f
C82 clkb0.t23 vssa 0.019975f
C83 clkb0.n5 vssa 0.026923f
C84 clkb0.n6 vssa 0.013183f
C85 clkb0.n7 vssa 0.028806f
C86 clkb0.n9 vssa 0.013183f
C87 clkb0.n10 vssa 0.028806f
C88 clkb0.t20 vssa 0.011771f
C89 clkb0.t31 vssa 0.019975f
C90 clkb0.n11 vssa 0.013183f
C91 clkb0.n12 vssa 0.028806f
C92 clkb0.n13 vssa 0.013183f
C93 clkb0.n16 vssa 0.062753f
C94 clkb0.n17 vssa 0.022752f
C95 clkb0.n21 vssa 0.013183f
C96 clkb0.n22 vssa 0.028806f
C97 clkb0.n23 vssa 0.013183f
C98 clkb0.n24 vssa 0.028806f
C99 clkb0.t30 vssa 0.011771f
C100 clkb0.t17 vssa 0.019975f
C101 clkb0.n25 vssa 0.026923f
C102 clkb0.n26 vssa 0.014085f
C103 clkb0.n28 vssa 0.045504f
C104 clkb0.n29 vssa 0.406567f
C105 clkb0.n30 vssa 0.024176f
C106 clkb0.t1 vssa 0.012841f
C107 clkb0.t7 vssa 0.012841f
C108 clkb0.n31 vssa 0.028544f
C109 clkb0.t0 vssa 0.012841f
C110 clkb0.t6 vssa 0.012841f
C111 clkb0.n32 vssa 0.028544f
C112 clkb0.t3 vssa 0.012841f
C113 clkb0.t5 vssa 0.012841f
C114 clkb0.n33 vssa 0.028544f
C115 clkb0.t2 vssa 0.012841f
C116 clkb0.t4 vssa 0.012841f
C117 clkb0.n34 vssa 0.028544f
C118 clkb0.n35 vssa 0.019009f
C119 clkb0.n36 vssa 0.019009f
C120 clkb0.n37 vssa 0.019009f
C121 clkb0.n38 vssa 0.019009f
C122 clkb0.n39 vssa 0.062442f
C123 clkb0.n40 vssa 0.056923f
C124 clkb0.n41 vssa 0.056923f
C125 clkb0.n42 vssa 0.065385f
C126 clkb0.n43 vssa 0.077689f
C127 clkb0.n44 vssa 0.074524f
C128 clkb0.n45 vssa 0.074524f
C129 clkb0.n46 vssa 0.077438f
C130 vdda.n2 vssa 0.017504f
C131 vdda.t12 vssa 0.092297f
C132 vdda.t8 vssa 0.040171f
C133 vdda.t44 vssa 0.040171f
C134 vdda.t27 vssa 0.040171f
C135 vdda.t41 vssa 0.040171f
C136 vdda.t25 vssa 0.040171f
C137 vdda.t23 vssa 0.040171f
C138 vdda.t46 vssa 0.043519f
C139 vdda.t34 vssa 0.054039f
C140 vdda.t18 vssa 0.040171f
C141 vdda.t4 vssa 0.040171f
C142 vdda.t31 vssa 0.040171f
C143 vdda.t6 vssa 0.040171f
C144 vdda.t2 vssa 0.040171f
C145 vdda.t59 vssa 0.040171f
C146 vdda.t15 vssa 0.043519f
C147 vdda.t29 vssa 0.051887f
C148 vdda.t48 vssa 0.040171f
C149 vdda.t10 vssa 0.040171f
C150 vdda.t0 vssa 0.038019f
C151 vdda.t67 vssa 0.065995f
C152 vdda.n6 vssa 0.024395f
C153 vdda.n11 vssa 0.01686f
C154 vdda.n12 vssa 0.02092f
C155 vdda.t39 vssa 0.050692f
C156 vdda.t21 vssa 0.036823f
C157 vdda.t36 vssa 0.049496f
C158 vdda.t61 vssa 0.058343f
C159 vdda.n13 vssa 0.033553f
C160 vdda.n14 vssa -0.018989f
C161 vdda.n16 vssa 0.0232f
C162 vdda.n20 vssa 0.011381f
C163 vdda.n37 vssa 0.018878f
C164 vdda.n41 vssa 0.010994f
C165 vdda.n46 vssa 0.024476f
C166 vdda.n52 vssa 0.016045f
C167 vdda.n57 vssa 0.01993f
C168 vdda.n70 vssa 0.016045f
C169 vdda.n76 vssa 0.011167f
C170 vdda.n83 vssa 0.017504f
C171 vdda.n92 vssa 0.022802f
.ends

