magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect 767 -2392 801 -2316
rect 1153 -2392 1187 -2316
rect 1153 -2482 1187 -2476
rect 1539 -2392 1573 -2316
rect 1539 -2482 1573 -2476
rect 1645 -2516 1679 -2316
rect 1645 -2606 1679 -2600
rect 2031 -2516 2065 -2316
rect 2031 -2606 2065 -2600
rect 2417 -2516 2451 -2316
rect 2417 -2606 2451 -2600
<< viali >>
rect 767 -2476 801 -2392
rect 1153 -2476 1187 -2392
rect 1539 -2476 1573 -2392
rect 1645 -2600 1679 -2516
rect 2031 -2600 2065 -2516
rect 2417 -2600 2451 -2516
<< metal1 >>
rect 931 -1829 951 -1777
rect 1003 -1829 1023 -1777
rect 1317 -1829 1337 -1777
rect 1389 -1829 1409 -1777
rect 861 -1919 867 -1867
rect 919 -1919 925 -1867
rect 861 -1991 925 -1919
rect 861 -2043 867 -1991
rect 919 -2043 925 -1991
rect 861 -2115 925 -2043
rect 861 -2167 867 -2115
rect 919 -2167 925 -2115
rect 1029 -2167 1311 -1867
rect 1415 -1919 1421 -1867
rect 1473 -1919 1479 -1867
rect 1415 -1991 1479 -1919
rect 1415 -2043 1421 -1991
rect 1473 -2043 1479 -1991
rect 1415 -2076 1479 -2043
rect 1809 -2047 1829 -1995
rect 1881 -2047 1901 -1995
rect 2195 -2047 2215 -1995
rect 2267 -2047 2287 -1995
rect 1415 -2115 1803 -2076
rect 1415 -2167 1421 -2115
rect 1473 -2167 1803 -2115
rect 1415 -2176 1803 -2167
rect 1907 -2176 2189 -2076
rect 2293 -2124 2357 -2076
rect 2293 -2176 2299 -2124
rect 2351 -2176 2357 -2124
rect 931 -2257 951 -2205
rect 1003 -2257 1023 -2205
rect 1317 -2257 1337 -2205
rect 1389 -2257 1409 -2205
rect 1809 -2257 1829 -2205
rect 1881 -2257 1901 -2205
rect 2195 -2257 2215 -2205
rect 2267 -2257 2287 -2205
rect 945 -2337 951 -2285
rect 1003 -2337 2215 -2285
rect 2267 -2337 2273 -2285
rect 731 -2392 867 -2386
rect 731 -2476 767 -2392
rect 801 -2476 867 -2392
rect 919 -2392 2487 -2386
rect 919 -2476 1153 -2392
rect 1187 -2476 1539 -2392
rect 1573 -2476 2487 -2392
rect 731 -2482 2487 -2476
rect 731 -2516 2299 -2510
rect 731 -2600 1645 -2516
rect 1679 -2600 2031 -2516
rect 2065 -2600 2299 -2516
rect 2351 -2516 2487 -2510
rect 2351 -2600 2417 -2516
rect 2451 -2600 2487 -2516
rect 731 -2606 2487 -2600
<< via1 >>
rect 951 -1829 1003 -1777
rect 1337 -1829 1389 -1777
rect 867 -1919 919 -1867
rect 867 -2043 919 -1991
rect 867 -2167 919 -2115
rect 1421 -1919 1473 -1867
rect 1421 -2043 1473 -1991
rect 1829 -2047 1881 -1995
rect 2215 -2047 2267 -1995
rect 1421 -2167 1473 -2115
rect 2299 -2176 2351 -2124
rect 951 -2257 1003 -2205
rect 1337 -2257 1389 -2205
rect 1829 -2257 1881 -2205
rect 2215 -2257 2267 -2205
rect 951 -2337 1003 -2285
rect 2215 -2337 2267 -2285
rect 867 -2476 919 -2386
rect 2299 -2600 2351 -2510
<< metal2 >>
rect 949 -1777 1005 -1771
rect 949 -1829 951 -1777
rect 1003 -1829 1005 -1777
rect 865 -1867 921 -1861
rect 865 -1919 867 -1867
rect 919 -1919 921 -1867
rect 865 -1991 921 -1919
rect 865 -2043 867 -1991
rect 919 -2043 921 -1991
rect 865 -2115 921 -2043
rect 865 -2167 867 -2115
rect 919 -2167 921 -2115
rect 865 -2386 921 -2167
rect 949 -2205 1005 -1829
rect 949 -2257 951 -2205
rect 1003 -2257 1005 -2205
rect 949 -2285 1005 -2257
rect 1335 -1777 1391 -1771
rect 1335 -1829 1337 -1777
rect 1389 -1829 1391 -1777
rect 1335 -2205 1391 -1829
rect 1419 -1867 1475 -1861
rect 1419 -1919 1421 -1867
rect 1473 -1919 1475 -1867
rect 1419 -1991 1475 -1919
rect 1419 -2043 1421 -1991
rect 1473 -2043 1475 -1991
rect 1419 -2115 1475 -2043
rect 1419 -2167 1421 -2115
rect 1473 -2167 1475 -2115
rect 1419 -2173 1475 -2167
rect 1827 -1995 1883 -1989
rect 1827 -2047 1829 -1995
rect 1881 -2047 1883 -1995
rect 1335 -2257 1337 -2205
rect 1389 -2257 1391 -2205
rect 1335 -2263 1391 -2257
rect 1827 -2205 1883 -2047
rect 1827 -2257 1829 -2205
rect 1881 -2257 1883 -2205
rect 1827 -2263 1883 -2257
rect 2213 -1995 2269 -1989
rect 2213 -2047 2215 -1995
rect 2267 -2047 2269 -1995
rect 2213 -2205 2269 -2047
rect 2213 -2257 2215 -2205
rect 2267 -2257 2269 -2205
rect 949 -2337 951 -2285
rect 1003 -2337 1005 -2285
rect 949 -2343 1005 -2337
rect 2213 -2285 2269 -2257
rect 2213 -2337 2215 -2285
rect 2267 -2337 2269 -2285
rect 2213 -2343 2269 -2337
rect 2297 -2124 2353 -2118
rect 2297 -2176 2299 -2124
rect 2351 -2176 2353 -2124
rect 865 -2476 867 -2386
rect 919 -2476 921 -2386
rect 865 -2482 921 -2476
rect 2297 -2510 2353 -2176
rect 2297 -2600 2299 -2510
rect 2351 -2600 2353 -2510
rect 2297 -2606 2353 -2600
use sky130_fd_pr__pfet_01v8_TMYSY6  XM1
timestamp 1730624594
transform 1 0 977 0 1 -2017
box -246 -369 246 369
use sky130_fd_pr__pfet_01v8_TMYSY6  XM2
timestamp 1730624594
transform 1 0 1363 0 1 -2017
box -246 -369 246 369
use sky130_fd_pr__nfet_01v8_SMGLWN  XM3
timestamp 1730624594
transform 1 0 1855 0 1 -2126
box -246 -260 246 260
use sky130_fd_pr__nfet_01v8_SMGLWN  XM4
timestamp 1730624594
transform 1 0 2241 0 1 -2126
box -246 -260 246 260
<< labels >>
flabel metal1 731 -2606 827 -2510 0 FreeSans 320 0 0 0 vssa
port 5 nsew
flabel metal1 731 -2482 827 -2386 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel via1 1337 -2257 1389 -2205 0 FreeSans 320 0 0 0 ckb
port 4 nsew
flabel via1 1829 -2257 1881 -2205 0 FreeSans 320 0 0 0 ck
port 3 nsew
flabel metal2 1421 -1919 1473 -1867 0 FreeSans 320 0 0 0 out
port 6 nsew
flabel metal2 2215 -2047 2267 -1995 0 FreeSans 320 0 0 0 in
port 2 nsew
<< end >>
