magic
tech sky130A
magscale 1 2
timestamp 1730845130
<< viali >>
rect 120 -1144 160 -1104
rect 1604 -1144 1644 -1104
rect 2054 -1144 2094 -1104
rect 3542 -1144 3582 -1104
rect 3984 -1144 4024 -1104
rect 5474 -1144 5514 -1104
rect 5916 -1144 5956 -1104
rect 7406 -1144 7446 -1104
rect 7848 -1144 7888 -1104
rect 9338 -1144 9378 -1104
rect -141 -1297 -101 -1257
rect 1791 -1297 1831 -1257
rect 3723 -1295 3763 -1255
rect 5655 -1295 5695 -1255
rect 7587 -1295 7627 -1255
<< metal1 >>
rect 104 -1150 114 -1098
rect 166 -1150 176 -1098
rect 1588 -1150 1598 -1098
rect 1650 -1150 1660 -1098
rect 2038 -1150 2048 -1098
rect 2100 -1150 2110 -1098
rect 3526 -1150 3536 -1098
rect 3588 -1150 3598 -1098
rect 3968 -1150 3978 -1098
rect 4030 -1150 4040 -1098
rect 5458 -1150 5468 -1098
rect 5520 -1150 5530 -1098
rect 5900 -1150 5910 -1098
rect 5962 -1150 5972 -1098
rect 7390 -1150 7400 -1098
rect 7452 -1150 7462 -1098
rect 7832 -1150 7842 -1098
rect 7894 -1150 7904 -1098
rect 9322 -1150 9332 -1098
rect 9384 -1150 9394 -1098
rect -157 -1303 -147 -1251
rect -95 -1303 -85 -1251
rect 1775 -1303 1785 -1251
rect 1837 -1303 1847 -1251
rect 3707 -1301 3717 -1249
rect 3769 -1301 3779 -1249
rect 5639 -1301 5649 -1249
rect 5701 -1301 5711 -1249
rect 7571 -1301 7581 -1249
rect 7633 -1301 7643 -1249
rect 1294 -1425 1304 -1373
rect 1356 -1425 1366 -1373
rect 3226 -1425 3236 -1373
rect 3288 -1425 3298 -1373
rect 5158 -1425 5168 -1373
rect 5220 -1425 5230 -1373
rect 7090 -1425 7100 -1373
rect 7152 -1425 7162 -1373
rect 9022 -1425 9032 -1373
rect 9084 -1425 9094 -1373
<< via1 >>
rect 114 -1104 166 -1098
rect 114 -1144 120 -1104
rect 120 -1144 160 -1104
rect 160 -1144 166 -1104
rect 114 -1150 166 -1144
rect 1598 -1104 1650 -1098
rect 1598 -1144 1604 -1104
rect 1604 -1144 1644 -1104
rect 1644 -1144 1650 -1104
rect 1598 -1150 1650 -1144
rect 2048 -1104 2100 -1098
rect 2048 -1144 2054 -1104
rect 2054 -1144 2094 -1104
rect 2094 -1144 2100 -1104
rect 2048 -1150 2100 -1144
rect 3536 -1104 3588 -1098
rect 3536 -1144 3542 -1104
rect 3542 -1144 3582 -1104
rect 3582 -1144 3588 -1104
rect 3536 -1150 3588 -1144
rect 3978 -1104 4030 -1098
rect 3978 -1144 3984 -1104
rect 3984 -1144 4024 -1104
rect 4024 -1144 4030 -1104
rect 3978 -1150 4030 -1144
rect 5468 -1104 5520 -1098
rect 5468 -1144 5474 -1104
rect 5474 -1144 5514 -1104
rect 5514 -1144 5520 -1104
rect 5468 -1150 5520 -1144
rect 5910 -1104 5962 -1098
rect 5910 -1144 5916 -1104
rect 5916 -1144 5956 -1104
rect 5956 -1144 5962 -1104
rect 5910 -1150 5962 -1144
rect 7400 -1104 7452 -1098
rect 7400 -1144 7406 -1104
rect 7406 -1144 7446 -1104
rect 7446 -1144 7452 -1104
rect 7400 -1150 7452 -1144
rect 7842 -1104 7894 -1098
rect 7842 -1144 7848 -1104
rect 7848 -1144 7888 -1104
rect 7888 -1144 7894 -1104
rect 7842 -1150 7894 -1144
rect 9332 -1104 9384 -1098
rect 9332 -1144 9338 -1104
rect 9338 -1144 9378 -1104
rect 9378 -1144 9384 -1104
rect 9332 -1150 9384 -1144
rect -147 -1257 -95 -1251
rect -147 -1297 -141 -1257
rect -141 -1297 -101 -1257
rect -101 -1297 -95 -1257
rect -147 -1303 -95 -1297
rect 1785 -1257 1837 -1251
rect 1785 -1297 1791 -1257
rect 1791 -1297 1831 -1257
rect 1831 -1297 1837 -1257
rect 1785 -1303 1837 -1297
rect 3717 -1255 3769 -1249
rect 3717 -1295 3723 -1255
rect 3723 -1295 3763 -1255
rect 3763 -1295 3769 -1255
rect 3717 -1301 3769 -1295
rect 5649 -1255 5701 -1249
rect 5649 -1295 5655 -1255
rect 5655 -1295 5695 -1255
rect 5695 -1295 5701 -1255
rect 5649 -1301 5701 -1295
rect 7581 -1255 7633 -1249
rect 7581 -1295 7587 -1255
rect 7587 -1295 7627 -1255
rect 7627 -1295 7633 -1255
rect 7581 -1301 7633 -1295
rect 1304 -1425 1356 -1373
rect 3236 -1425 3288 -1373
rect 5168 -1425 5220 -1373
rect 7100 -1425 7152 -1373
rect 9032 -1425 9084 -1373
<< metal2 >>
rect 114 -1098 166 -1088
rect 114 -1160 166 -1150
rect 1598 -1098 1650 -1088
rect 1598 -1160 1650 -1150
rect 2048 -1098 2100 -1088
rect 2048 -1160 2100 -1150
rect 3536 -1098 3588 -1088
rect 3536 -1160 3588 -1150
rect 3978 -1098 4030 -1088
rect 5468 -1098 5520 -1088
rect 4030 -1150 4031 -1098
rect 3978 -1160 4030 -1150
rect 5468 -1160 5520 -1150
rect 5910 -1098 5962 -1088
rect 7400 -1098 7452 -1088
rect 5962 -1150 5963 -1098
rect 5910 -1160 5962 -1150
rect 7400 -1160 7452 -1150
rect 7842 -1098 7894 -1088
rect 9332 -1098 9384 -1088
rect 7894 -1150 7895 -1098
rect 7842 -1160 7894 -1150
rect 9332 -1160 9384 -1150
rect -147 -1251 -95 -1241
rect 1785 -1251 1837 -1241
rect 3717 -1249 3769 -1239
rect -178 -1301 -147 -1251
rect -95 -1301 1785 -1251
rect -147 -1313 -95 -1303
rect 1837 -1301 3717 -1251
rect 5649 -1249 5701 -1239
rect 3769 -1301 5649 -1251
rect 7581 -1249 7633 -1239
rect 5701 -1301 7581 -1251
rect 1785 -1313 1837 -1303
rect 3717 -1311 3769 -1301
rect 5649 -1311 5701 -1301
rect 7581 -1311 7633 -1301
rect 1304 -1373 1356 -1363
rect 3236 -1373 3288 -1363
rect 5168 -1373 5220 -1363
rect 7100 -1373 7152 -1363
rect 9032 -1373 9084 -1363
rect -178 -1425 1304 -1373
rect 1356 -1425 3236 -1373
rect 3288 -1425 5168 -1373
rect 5220 -1425 7100 -1373
rect 7152 -1425 9032 -1373
rect 1304 -1435 1356 -1425
rect 3236 -1435 3288 -1425
rect 5168 -1435 5220 -1425
rect 7100 -1435 7152 -1425
rect 9032 -1435 9084 -1425
use sky130_fd_sc_hd__dfrtp_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730336909
transform 1 0 -167 0 1 -1566
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2
timestamp 1730336909
transform 1 0 1765 0 1 -1566
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3
timestamp 1730336909
transform 1 0 3697 0 1 -1566
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4
timestamp 1730336909
transform 1 0 5629 0 1 -1566
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x6
timestamp 1730336909
transform 1 0 7561 0 1 -1566
box -38 -48 1970 592
<< labels >>
flabel space -116 -990 -116 -990 0 FreeSans 160 0 0 0 VPWR
port 4 nsew
flabel space -75 -1599 -75 -1599 0 FreeSans 160 0 0 0 VGND
port 5 nsew
<< end >>
