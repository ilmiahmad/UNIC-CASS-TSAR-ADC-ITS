magic
tech sky130A
magscale 1 2
timestamp 1730671942
<< nwell >>
rect 22487 4423 22713 4649
rect 10848 2130 11074 2356
rect 10849 1191 11075 1417
<< pwell >>
rect 10806 1980 10896 1982
rect 1132 1753 10896 1980
rect 969 1576 10896 1753
rect 969 1571 1245 1576
<< psubdiff >>
rect 10846 1822 10888 1846
rect 10846 1702 10888 1726
<< nsubdiff >>
rect 22523 4579 22583 4613
rect 22617 4579 22677 4613
rect 22523 4553 22557 4579
rect 22523 4493 22557 4519
rect 22643 4553 22677 4579
rect 22643 4493 22677 4519
rect 22523 4459 22583 4493
rect 22617 4459 22677 4493
rect 10884 2286 10944 2320
rect 10978 2286 11038 2320
rect 10884 2260 10918 2286
rect 10884 2200 10918 2226
rect 11004 2260 11038 2286
rect 11004 2200 11038 2226
rect 10884 2166 10944 2200
rect 10978 2166 11038 2200
rect 10885 1347 10945 1381
rect 10979 1347 11039 1381
rect 10885 1321 10919 1347
rect 10885 1261 10919 1287
rect 11005 1321 11039 1347
rect 11005 1261 11039 1287
rect 10885 1227 10945 1261
rect 10979 1227 11039 1261
<< psubdiffcont >>
rect 10846 1726 10888 1822
<< nsubdiffcont >>
rect 22583 4579 22617 4613
rect 22523 4519 22557 4553
rect 22643 4519 22677 4553
rect 22583 4459 22617 4493
rect 10944 2286 10978 2320
rect 10884 2226 10918 2260
rect 11004 2226 11038 2260
rect 10944 2166 10978 2200
rect 10945 1347 10979 1381
rect 10885 1287 10919 1321
rect 11005 1287 11039 1321
rect 10945 1227 10979 1261
<< locali >>
rect 22523 4579 22583 4613
rect 22617 4579 22677 4613
rect 22523 4553 22557 4579
rect 22523 4493 22557 4519
rect 22643 4553 22677 4579
rect 22643 4493 22677 4519
rect 22523 4459 22583 4493
rect 22617 4459 22677 4493
rect 10884 2286 10944 2320
rect 10978 2286 11038 2320
rect 10884 2260 10918 2286
rect 10884 2200 10918 2226
rect 11004 2260 11038 2286
rect 11004 2200 11038 2226
rect 10884 2166 10944 2200
rect 10978 2166 11038 2200
rect 10846 1822 10888 1838
rect 10846 1710 10888 1726
rect 136 1512 294 1563
rect 10885 1347 10945 1381
rect 10979 1347 11039 1381
rect 10885 1321 10919 1347
rect 10885 1261 10919 1287
rect 11005 1321 11039 1347
rect 11005 1261 11039 1287
rect 10885 1227 10945 1261
rect 10979 1227 11039 1261
<< viali >>
rect 10944 2286 10978 2320
rect 10944 2166 10978 2200
rect 10846 1726 10888 1822
rect 85 1512 136 1563
rect 1074 1525 1108 1559
rect 10945 1347 10979 1381
rect 10945 1227 10979 1261
<< metal1 >>
rect 10718 2320 11038 2366
rect 10718 2286 10944 2320
rect 10978 2286 11038 2320
rect 10718 2270 11038 2286
rect 10882 2200 11038 2270
rect 10882 2166 10944 2200
rect 10978 2166 11038 2200
rect 10882 2130 11038 2166
rect 10840 1822 10894 1834
rect -98 1726 48 1822
rect 10804 1726 10846 1822
rect 10888 1726 10894 1822
rect 10840 1714 10894 1726
rect -91 1512 -85 1564
rect -33 1563 -27 1564
rect 79 1563 142 1575
rect 1066 1568 1118 1574
rect -33 1512 85 1563
rect 136 1512 142 1563
rect 1062 1519 1066 1565
rect 79 1500 142 1512
rect 1118 1519 1120 1565
rect 1066 1510 1118 1516
rect 10942 1418 11038 2130
rect 10884 1381 11038 1418
rect 10884 1347 10945 1381
rect 10979 1347 11038 1381
rect 10884 1278 11038 1347
rect -168 1182 110 1278
rect 10740 1261 11038 1278
rect 10740 1227 10945 1261
rect 10979 1227 11038 1261
rect 10740 1182 11038 1227
<< via1 >>
rect -85 1512 -33 1564
rect 1066 1559 1118 1568
rect 1066 1525 1074 1559
rect 1074 1525 1108 1559
rect 1108 1525 1118 1559
rect 1066 1516 1118 1525
<< metal2 >>
rect -98 2191 1037 2241
rect 3314 2190 3366 2602
rect 5244 2190 5296 2602
rect 7176 2190 7228 2602
rect 9108 2190 9160 2602
rect 10697 2241 10747 2602
rect 10649 2191 11065 2241
rect -87 2039 1051 2089
rect 3051 2032 3060 2088
rect 3116 2032 3125 2088
rect -84 1915 1036 1967
rect 1612 1581 1664 1966
rect -85 1564 -33 1570
rect -169 1513 -85 1564
rect 1060 1516 1066 1568
rect 1118 1516 1188 1568
rect -85 1506 -33 1512
rect 1136 1358 1188 1516
rect 3058 1514 3118 1523
rect 3058 1445 3118 1454
rect 1136 1306 1312 1358
rect 1226 918 1278 1306
rect 2802 918 2854 1358
rect 4734 910 4786 1358
rect 6666 910 6718 1358
rect 8596 910 8648 1358
rect 11015 1357 11065 2191
rect 10932 1307 11065 1357
<< via2 >>
rect 3060 2032 3116 2088
rect 3058 1454 3118 1514
<< metal3 >>
rect 3055 2088 3121 2093
rect 3055 2032 3060 2088
rect 3116 2032 3121 2088
rect 3055 2027 3121 2032
rect 3058 1519 3118 2027
rect 3053 1514 3123 1519
rect 3053 1454 3058 1514
rect 3118 1454 3123 1514
rect 3053 1449 3123 1454
use buf  buf_0
timestamp 1730671111
transform -1 0 2036 0 -1 2540
box 846 718 2026 1358
use flip_flop_5  flip_flop_5_0
timestamp 1730670220
transform 1 0 1318 0 1 3340
box -342 -1614 9531 -974
use flip_flop_5  flip_flop_5_1
timestamp 1730670220
transform -1 0 10644 0 -1 208
box -342 -1614 9531 -974
<< labels >>
flabel metal2 -60 2216 -60 2216 0 FreeSans 800 0 0 0 EN
port 0 nsew
flabel metal1 -76 1768 -76 1768 0 FreeSans 800 0 0 0 VSSD
port 3 nsew
flabel metal2 -80 2054 -80 2054 0 FreeSans 800 0 0 0 RDY
port 16 nsew
flabel metal2 -72 1940 -72 1940 0 FreeSans 800 0 0 0 CLKS
port 17 nsew
flabel metal1 -152 1228 -152 1228 0 FreeSans 800 0 0 0 VDDD
port 4 nsew
flabel metal2 -142 1538 -142 1538 0 FreeSans 800 0 0 0 FINAL
port 18 nsew
flabel metal2 3338 2548 3338 2550 0 FreeSans 800 0 0 0 CF[0]
port 19 nsew
flabel metal2 5274 2554 5274 2556 0 FreeSans 800 0 0 0 CF[1]
port 20 nsew
flabel metal2 7202 2564 7202 2566 0 FreeSans 800 0 0 0 CF[2]
port 21 nsew
flabel metal2 9132 2556 9132 2558 0 FreeSans 800 0 0 0 CF[3]
port 22 nsew
flabel metal2 10718 2552 10718 2554 0 FreeSans 800 0 0 0 CF[4]
port 23 nsew
flabel metal2 8618 966 8618 968 0 FreeSans 800 0 0 0 CF[5]
port 24 nsew
flabel metal2 6684 948 6684 950 0 FreeSans 800 0 0 0 CF[6]
port 25 nsew
flabel metal2 4754 942 4754 944 0 FreeSans 800 0 0 0 CF[7]
port 26 nsew
flabel metal2 2822 956 2822 958 0 FreeSans 800 0 0 0 CF[8]
port 27 nsew
flabel metal2 1252 956 1260 964 0 FreeSans 800 0 0 0 CF[9]
port 28 nsew
<< end >>
