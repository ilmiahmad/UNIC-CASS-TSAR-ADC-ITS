magic
tech sky130A
magscale 1 2
timestamp 1730626724
<< metal1 >>
rect 102622 -2422 102628 -2318
rect 102806 -2422 103334 -2318
rect 135331 -2422 135854 -2318
rect 136032 -2422 136038 -2318
rect 102834 -4206 102840 -4110
rect 103018 -4206 103326 -4110
rect 135334 -4206 135642 -4110
rect 135820 -4206 135826 -4110
rect 103046 -4750 103052 -4654
rect 103230 -4750 103326 -4654
rect 135334 -4750 135430 -4654
rect 135608 -4750 135614 -4654
rect 102834 -5293 102840 -5197
rect 103018 -5293 103326 -5197
rect 135430 -5198 135642 -5197
rect 135334 -5293 135642 -5198
rect 135820 -5293 135826 -5197
rect 102834 -5294 103230 -5293
rect 135334 -5294 135826 -5293
rect 102622 -5380 102628 -5322
rect 102806 -5380 103288 -5322
rect 135372 -5380 135854 -5322
rect 136032 -5380 136038 -5322
rect 102834 -5504 102840 -5408
rect 103018 -5504 103326 -5408
rect 135334 -5504 135642 -5408
rect 135820 -5504 135826 -5408
rect 103046 -5628 103052 -5532
rect 103230 -5628 103326 -5532
rect 135334 -5628 135430 -5532
rect 135608 -5628 135614 -5532
rect 103046 -15494 103052 -15398
rect 103230 -15494 103326 -15398
rect 135334 -15494 135430 -15398
rect 135608 -15494 135614 -15398
rect 102834 -15618 102840 -15522
rect 103018 -15618 103326 -15522
rect 135334 -15618 135642 -15522
rect 135820 -15618 135826 -15522
rect 102622 -15704 102628 -15646
rect 102806 -15704 103288 -15646
rect 135372 -15704 135854 -15646
rect 136032 -15704 136038 -15646
rect 102834 -15733 103326 -15732
rect 135430 -15733 135826 -15732
rect 102834 -15829 102840 -15733
rect 103018 -15828 103326 -15733
rect 103018 -15829 103230 -15828
rect 135334 -15829 135642 -15733
rect 135820 -15829 135826 -15733
rect 103046 -16372 103052 -16276
rect 103230 -16372 103326 -16276
rect 135334 -16372 135430 -16276
rect 135608 -16372 135614 -16276
rect 102834 -16916 102840 -16820
rect 103018 -16916 103326 -16820
rect 135334 -16916 135642 -16820
rect 135820 -16916 135826 -16820
rect 102622 -18708 102628 -18604
rect 102806 -18708 103329 -18604
rect 135326 -18708 135854 -18604
rect 136032 -18708 136038 -18604
<< via1 >>
rect 102628 -2422 102806 -2318
rect 135854 -2422 136032 -2318
rect 132592 -2580 132684 -2488
rect 129372 -2744 129464 -2652
rect 126152 -2908 126244 -2816
rect 122932 -3072 123024 -2980
rect 119712 -3236 119804 -3144
rect 116492 -3400 116584 -3308
rect 113272 -3564 113364 -3472
rect 110052 -3728 110144 -3636
rect 106832 -3892 106924 -3800
rect 103612 -4056 103704 -3964
rect 102840 -4206 103018 -4110
rect 135642 -4206 135820 -4110
rect 103052 -4750 103230 -4654
rect 135430 -4750 135608 -4654
rect 102840 -5293 103018 -5197
rect 135642 -5293 135820 -5197
rect 102628 -5380 102806 -5322
rect 135854 -5380 136032 -5322
rect 102840 -5504 103018 -5408
rect 135642 -5504 135820 -5408
rect 103052 -5628 103230 -5532
rect 135430 -5628 135608 -5532
rect 103052 -15494 103230 -15398
rect 135430 -15494 135608 -15398
rect 102840 -15618 103018 -15522
rect 135642 -15618 135820 -15522
rect 102628 -15704 102806 -15646
rect 135854 -15704 136032 -15646
rect 102840 -15829 103018 -15733
rect 135642 -15829 135820 -15733
rect 103052 -16372 103230 -16276
rect 135430 -16372 135608 -16276
rect 102840 -16916 103018 -16820
rect 135642 -16916 135820 -16820
rect 134956 -17062 135048 -16970
rect 131736 -17226 131828 -17134
rect 128516 -17390 128608 -17298
rect 125296 -17554 125388 -17462
rect 122076 -17718 122168 -17626
rect 118856 -17882 118948 -17790
rect 115636 -18046 115728 -17954
rect 112416 -18210 112508 -18118
rect 109196 -18374 109288 -18282
rect 105976 -18538 106068 -18446
rect 102628 -18708 102806 -18604
rect 135854 -18708 136032 -18604
<< metal2 >>
rect 102622 -2318 102806 19876
rect 102622 -2422 102628 -2318
rect 102622 -5322 102806 -2422
rect 102622 -5380 102628 -5322
rect 102622 -15646 102806 -5380
rect 102622 -15704 102628 -15646
rect 102622 -18604 102806 -15704
rect 102622 -18708 102628 -18604
rect 102622 -40902 102806 -18708
rect 102834 -4110 103018 19876
rect 102834 -4206 102840 -4110
rect 102834 -5197 103018 -4206
rect 102834 -5293 102840 -5197
rect 102834 -5408 103018 -5293
rect 102834 -5504 102840 -5408
rect 102834 -15522 103018 -5504
rect 102834 -15618 102840 -15522
rect 102834 -15733 103018 -15618
rect 102834 -15829 102840 -15733
rect 102834 -16820 103018 -15829
rect 102834 -16916 102840 -16820
rect 102834 -40902 103018 -16916
rect 103046 -4654 103230 19876
rect 132586 -2488 132690 -2482
rect 132586 -2580 132592 -2488
rect 132684 -2580 132690 -2488
rect 129366 -2652 129470 -2646
rect 129366 -2744 129372 -2652
rect 129464 -2744 129470 -2652
rect 126146 -2816 126250 -2810
rect 126146 -2908 126152 -2816
rect 126244 -2908 126250 -2816
rect 122926 -2980 123030 -2974
rect 122926 -3072 122932 -2980
rect 123024 -3072 123030 -2980
rect 119706 -3144 119810 -3138
rect 119706 -3236 119712 -3144
rect 119804 -3236 119810 -3144
rect 116486 -3308 116590 -3302
rect 116486 -3400 116492 -3308
rect 116584 -3400 116590 -3308
rect 113266 -3472 113370 -3466
rect 113266 -3564 113272 -3472
rect 113364 -3564 113370 -3472
rect 110046 -3636 110150 -3630
rect 110046 -3728 110052 -3636
rect 110144 -3728 110150 -3636
rect 106826 -3800 106930 -3794
rect 106826 -3892 106832 -3800
rect 106924 -3892 106930 -3800
rect 103046 -4750 103052 -4654
rect 103046 -5532 103230 -4750
rect 103606 -3964 103710 -3958
rect 103606 -4056 103612 -3964
rect 103704 -4056 103710 -3964
rect 103046 -5628 103052 -5532
rect 103046 -15398 103230 -5628
rect 103474 -5541 103578 -5532
rect 103474 -5883 103578 -5623
rect 103474 -5950 103578 -5941
rect 103606 -6011 103710 -4056
rect 106694 -5385 106798 -5376
rect 106694 -5883 106798 -5467
rect 106694 -5950 106798 -5941
rect 103606 -6078 103710 -6069
rect 106826 -6011 106930 -3892
rect 106826 -6078 106930 -6069
rect 109914 -5229 110018 -5220
rect 109914 -6419 110018 -5311
rect 109914 -6486 110018 -6477
rect 110046 -6547 110150 -3728
rect 113134 -5073 113238 -5064
rect 113134 -6419 113238 -5155
rect 113134 -6486 113238 -6477
rect 110046 -6614 110150 -6605
rect 113266 -6547 113370 -3564
rect 113266 -6614 113370 -6605
rect 116354 -4917 116458 -4908
rect 103046 -15494 103052 -15398
rect 103046 -16276 103230 -15494
rect 103046 -16372 103052 -16276
rect 103046 -40902 103230 -16372
rect 105970 -6917 106074 -6908
rect 105970 -18446 106074 -6975
rect 109190 -6917 109294 -6908
rect 106102 -7045 106206 -7036
rect 106102 -16807 106206 -7103
rect 106102 -16898 106206 -16889
rect 109190 -18282 109294 -6975
rect 109322 -7045 109426 -7036
rect 109322 -16651 109426 -7103
rect 116354 -7491 116458 -4999
rect 116354 -7558 116458 -7549
rect 116486 -7619 116590 -3400
rect 119574 -4761 119678 -4752
rect 119574 -7491 119678 -4843
rect 119574 -7558 119678 -7549
rect 116486 -7686 116590 -7677
rect 119706 -7619 119810 -3236
rect 119706 -7686 119810 -7677
rect 122794 -4605 122898 -4596
rect 122794 -8563 122898 -4687
rect 122794 -8754 122898 -8621
rect 122926 -8691 123030 -3072
rect 122926 -8758 123030 -8749
rect 126014 -4449 126118 -4440
rect 126014 -8563 126118 -4531
rect 126014 -8754 126118 -8621
rect 126146 -8691 126250 -2908
rect 126146 -8758 126250 -8749
rect 129234 -4293 129338 -4284
rect 109322 -16742 109426 -16733
rect 112410 -12277 112514 -12268
rect 112410 -18118 112514 -12335
rect 112542 -12405 112646 -12272
rect 112542 -16495 112646 -12463
rect 112542 -16586 112646 -16577
rect 115630 -12277 115734 -12268
rect 115630 -17954 115734 -12335
rect 115762 -12405 115866 -12272
rect 115762 -16339 115866 -12463
rect 115762 -16430 115866 -16421
rect 118850 -13349 118954 -13340
rect 118850 -17790 118954 -13407
rect 122070 -13349 122174 -13340
rect 118982 -13477 119086 -13468
rect 118982 -16183 119086 -13535
rect 118982 -16274 119086 -16265
rect 122070 -17626 122174 -13407
rect 122202 -13477 122306 -13468
rect 122202 -16027 122306 -13535
rect 129234 -13923 129338 -4375
rect 129234 -13990 129338 -13981
rect 129366 -14051 129470 -2744
rect 132454 -4137 132558 -4128
rect 132454 -13923 132558 -4219
rect 132454 -13990 132558 -13981
rect 129366 -14118 129470 -14109
rect 132586 -14051 132690 -2580
rect 132586 -14118 132690 -14109
rect 135430 -4654 135614 19876
rect 135608 -4750 135614 -4654
rect 135430 -5532 135614 -4750
rect 135608 -5628 135614 -5532
rect 122202 -16118 122306 -16109
rect 125290 -14421 125394 -14412
rect 125290 -17462 125394 -14479
rect 128510 -14421 128614 -14412
rect 125422 -14549 125526 -14540
rect 125422 -15871 125526 -14607
rect 125422 -15962 125526 -15953
rect 128510 -17298 128614 -14479
rect 128642 -14549 128746 -14540
rect 128642 -15715 128746 -14607
rect 128642 -15806 128746 -15797
rect 131730 -14957 131834 -14948
rect 131730 -17134 131834 -15015
rect 134950 -14957 135054 -14948
rect 131862 -15085 131966 -15076
rect 131862 -15559 131966 -15143
rect 131862 -15650 131966 -15641
rect 134950 -16970 135054 -15015
rect 135082 -15085 135186 -15076
rect 135082 -15403 135186 -15143
rect 135082 -15494 135186 -15485
rect 135430 -15398 135614 -5628
rect 135608 -15494 135614 -15398
rect 134950 -17062 134956 -16970
rect 135048 -17062 135054 -16970
rect 134950 -17068 135054 -17062
rect 135430 -16276 135614 -15494
rect 135608 -16372 135614 -16276
rect 131730 -17226 131736 -17134
rect 131828 -17226 131834 -17134
rect 131730 -17232 131834 -17226
rect 128510 -17390 128516 -17298
rect 128608 -17390 128614 -17298
rect 128510 -17396 128614 -17390
rect 125290 -17554 125296 -17462
rect 125388 -17554 125394 -17462
rect 125290 -17560 125394 -17554
rect 122070 -17718 122076 -17626
rect 122168 -17718 122174 -17626
rect 122070 -17724 122174 -17718
rect 118850 -17882 118856 -17790
rect 118948 -17882 118954 -17790
rect 118850 -17888 118954 -17882
rect 115630 -18046 115636 -17954
rect 115728 -18046 115734 -17954
rect 115630 -18052 115734 -18046
rect 112410 -18210 112416 -18118
rect 112508 -18210 112514 -18118
rect 112410 -18216 112514 -18210
rect 109190 -18374 109196 -18282
rect 109288 -18374 109294 -18282
rect 109190 -18380 109294 -18374
rect 105970 -18538 105976 -18446
rect 106068 -18538 106074 -18446
rect 105970 -18544 106074 -18538
rect 135430 -40903 135614 -16372
rect 135642 -4110 135826 19876
rect 135820 -4206 135826 -4110
rect 135642 -5197 135826 -4206
rect 135820 -5293 135826 -5197
rect 135642 -5408 135826 -5293
rect 135820 -5504 135826 -5408
rect 135642 -15522 135826 -5504
rect 135820 -15618 135826 -15522
rect 135642 -15733 135826 -15618
rect 135820 -15829 135826 -15733
rect 135642 -16820 135826 -15829
rect 135820 -16916 135826 -16820
rect 135642 -40903 135826 -16916
rect 135854 -2318 136038 19876
rect 136032 -2422 136038 -2318
rect 135854 -5322 136038 -2422
rect 136032 -5380 136038 -5322
rect 135854 -15646 136038 -5380
rect 136032 -15704 136038 -15646
rect 135854 -18604 136038 -15704
rect 136032 -18708 136038 -18604
rect 135854 -40903 136038 -18708
<< via2 >>
rect 103474 -5623 103578 -5541
rect 103474 -5941 103578 -5883
rect 106694 -5467 106798 -5385
rect 106694 -5941 106798 -5883
rect 103606 -6069 103710 -6011
rect 106826 -6069 106930 -6011
rect 109914 -5311 110018 -5229
rect 109914 -6477 110018 -6419
rect 113134 -5155 113238 -5073
rect 113134 -6477 113238 -6419
rect 110046 -6605 110150 -6547
rect 113266 -6605 113370 -6547
rect 116354 -4999 116458 -4917
rect 105970 -6975 106074 -6917
rect 109190 -6975 109294 -6917
rect 106102 -7103 106206 -7045
rect 106102 -16889 106206 -16807
rect 109322 -7103 109426 -7045
rect 116354 -7549 116458 -7491
rect 119574 -4843 119678 -4761
rect 119574 -7549 119678 -7491
rect 116486 -7677 116590 -7619
rect 119706 -7677 119810 -7619
rect 122794 -4687 122898 -4605
rect 122794 -8621 122898 -8563
rect 122926 -8749 123030 -8691
rect 126014 -4531 126118 -4449
rect 126014 -8621 126118 -8563
rect 126146 -8749 126250 -8691
rect 129234 -4375 129338 -4293
rect 109322 -16733 109426 -16651
rect 112410 -12335 112514 -12277
rect 112542 -12463 112646 -12405
rect 112542 -16577 112646 -16495
rect 115630 -12335 115734 -12277
rect 115762 -12463 115866 -12405
rect 115762 -16421 115866 -16339
rect 118850 -13407 118954 -13349
rect 122070 -13407 122174 -13349
rect 118982 -13535 119086 -13477
rect 118982 -16265 119086 -16183
rect 122202 -13535 122306 -13477
rect 129234 -13981 129338 -13923
rect 132454 -4219 132558 -4137
rect 132454 -13981 132558 -13923
rect 129366 -14109 129470 -14051
rect 132586 -14109 132690 -14051
rect 122202 -16109 122306 -16027
rect 125290 -14479 125394 -14421
rect 128510 -14479 128614 -14421
rect 125422 -14607 125526 -14549
rect 125422 -15953 125526 -15871
rect 128642 -14607 128746 -14549
rect 128642 -15797 128746 -15715
rect 131730 -15015 131834 -14957
rect 134950 -15015 135054 -14957
rect 131862 -15143 131966 -15085
rect 131862 -15641 131966 -15559
rect 135082 -15143 135186 -15085
rect 135082 -15485 135186 -15403
<< metal3 >>
rect 102622 -4137 136038 -4128
rect 102622 -4219 132454 -4137
rect 132558 -4219 136038 -4137
rect 102622 -4224 136038 -4219
rect 102622 -4293 136038 -4284
rect 102622 -4375 129234 -4293
rect 129338 -4375 136038 -4293
rect 102622 -4380 136038 -4375
rect 102622 -4449 136038 -4440
rect 102622 -4531 126014 -4449
rect 126118 -4531 136038 -4449
rect 102622 -4536 136038 -4531
rect 102622 -4605 136038 -4596
rect 102622 -4687 122794 -4605
rect 122898 -4687 136038 -4605
rect 102622 -4692 136038 -4687
rect 102622 -4761 136038 -4752
rect 102622 -4843 119574 -4761
rect 119678 -4843 136038 -4761
rect 102622 -4848 136038 -4843
rect 102622 -4917 136038 -4908
rect 102622 -4999 116354 -4917
rect 116458 -4999 136038 -4917
rect 102622 -5004 136038 -4999
rect 102622 -5073 136038 -5064
rect 102622 -5155 113134 -5073
rect 113238 -5155 136038 -5073
rect 102622 -5160 136038 -5155
rect 102622 -5229 136038 -5220
rect 102622 -5311 109914 -5229
rect 110018 -5311 136038 -5229
rect 102622 -5316 136038 -5311
rect 102622 -5385 136038 -5376
rect 102622 -5467 106694 -5385
rect 106798 -5467 136038 -5385
rect 102622 -5472 136038 -5467
rect 102622 -5541 136038 -5532
rect 102622 -5623 103474 -5541
rect 103578 -5623 136038 -5541
rect 102622 -5628 136038 -5623
rect 103474 -5883 103578 -5878
rect 103474 -5946 103578 -5941
rect 103606 -6011 103710 -6006
rect 103606 -6074 103710 -6069
rect 102622 -9764 136038 -9763
rect 102622 -9858 103299 -9764
rect 103401 -9858 135259 -9764
rect 135361 -9858 136038 -9764
rect 102622 -9859 136038 -9858
rect 102622 -9920 136038 -9919
rect 102622 -10014 106519 -9920
rect 106621 -10014 132039 -9920
rect 132141 -10014 136038 -9920
rect 102622 -10015 136038 -10014
rect 102622 -10076 136038 -10075
rect 102622 -10170 109739 -10076
rect 109841 -10170 128819 -10076
rect 128921 -10170 136038 -10076
rect 102622 -10171 136038 -10170
rect 102622 -10232 136038 -10231
rect 102622 -10326 112959 -10232
rect 113061 -10326 125599 -10232
rect 125701 -10326 136038 -10232
rect 102622 -10327 136038 -10326
rect 102622 -10388 136038 -10387
rect 102622 -10482 116179 -10388
rect 116281 -10482 122379 -10388
rect 122481 -10482 136038 -10388
rect 102622 -10483 136038 -10482
rect 102622 -10544 136038 -10543
rect 102622 -10638 119159 -10544
rect 119261 -10638 119399 -10544
rect 119501 -10638 136038 -10544
rect 102622 -10639 136038 -10638
rect 102622 -10700 136038 -10699
rect 102622 -10794 115939 -10700
rect 116041 -10794 122619 -10700
rect 122721 -10794 136038 -10700
rect 102622 -10795 136038 -10794
rect 102622 -10856 136038 -10855
rect 102622 -10950 112719 -10856
rect 112821 -10950 125839 -10856
rect 125941 -10950 136038 -10856
rect 102622 -10951 136038 -10950
rect 102622 -11012 136038 -11011
rect 102622 -11106 109499 -11012
rect 109601 -11106 129059 -11012
rect 129161 -11106 136038 -11012
rect 102622 -11107 136038 -11106
rect 102622 -11168 136038 -11167
rect 102622 -11262 106279 -11168
rect 106381 -11262 132279 -11168
rect 132381 -11262 136038 -11168
rect 102622 -11263 136038 -11262
rect 134950 -14957 135054 -14952
rect 134950 -15020 135054 -15015
rect 135082 -15085 135186 -15080
rect 135082 -15148 135186 -15143
rect 102622 -15403 136038 -15398
rect 102622 -15485 135082 -15403
rect 135186 -15485 136038 -15403
rect 102622 -15494 136038 -15485
rect 102622 -15559 136038 -15554
rect 102622 -15641 131862 -15559
rect 131966 -15641 136038 -15559
rect 102622 -15650 136038 -15641
rect 102622 -15715 136038 -15710
rect 102622 -15797 128642 -15715
rect 128746 -15797 136038 -15715
rect 102622 -15806 136038 -15797
rect 102622 -15871 136038 -15866
rect 102622 -15953 125422 -15871
rect 125526 -15953 136038 -15871
rect 102622 -15962 136038 -15953
rect 102622 -16027 136038 -16022
rect 102622 -16109 122202 -16027
rect 122306 -16109 136038 -16027
rect 102622 -16118 136038 -16109
rect 102622 -16183 136038 -16178
rect 102622 -16265 118982 -16183
rect 119086 -16265 136038 -16183
rect 102622 -16274 136038 -16265
rect 102622 -16339 136038 -16334
rect 102622 -16421 115762 -16339
rect 115866 -16421 136038 -16339
rect 102622 -16430 136038 -16421
rect 102622 -16495 136038 -16490
rect 102622 -16577 112542 -16495
rect 112646 -16577 136038 -16495
rect 102622 -16586 136038 -16577
rect 102622 -16651 136038 -16646
rect 102622 -16733 109322 -16651
rect 109426 -16733 136038 -16651
rect 102622 -16742 136038 -16733
rect 102622 -16807 136038 -16802
rect 102622 -16889 106102 -16807
rect 106206 -16889 136038 -16807
rect 102622 -16898 136038 -16889
<< via3 >>
rect 103299 -5817 103401 -5751
rect 106519 -5817 106621 -5751
rect 109739 -6353 109841 -6287
rect 112959 -6353 113061 -6287
rect 106279 -7235 106381 -7169
rect 109499 -7235 109601 -7169
rect 116179 -7425 116281 -7359
rect 119399 -7425 119501 -7359
rect 122619 -8497 122721 -8431
rect 125839 -8497 125941 -8431
rect 103299 -9858 103401 -9764
rect 135259 -9858 135361 -9764
rect 106519 -10014 106621 -9920
rect 132039 -10014 132141 -9920
rect 109739 -10170 109841 -10076
rect 128819 -10170 128921 -10076
rect 112959 -10326 113061 -10232
rect 125599 -10326 125701 -10232
rect 116179 -10482 116281 -10388
rect 122379 -10482 122481 -10388
rect 119159 -10638 119261 -10544
rect 119399 -10638 119501 -10544
rect 115939 -10794 116041 -10700
rect 122619 -10794 122721 -10700
rect 112719 -10950 112821 -10856
rect 125839 -10950 125941 -10856
rect 109499 -11106 109601 -11012
rect 129059 -11106 129161 -11012
rect 106279 -11262 106381 -11168
rect 132279 -11262 132381 -11168
rect 112719 -12595 112821 -12529
rect 115939 -12595 116041 -12529
rect 119159 -13667 119261 -13601
rect 122379 -13667 122481 -13601
rect 129059 -13857 129161 -13791
rect 132279 -13857 132381 -13791
rect 125599 -14739 125701 -14673
rect 128819 -14739 128921 -14673
rect 132039 -15275 132141 -15209
rect 135259 -15275 135361 -15209
<< metal4 >>
rect 103298 -5751 103402 -5750
rect 103298 -5817 103299 -5751
rect 103401 -5817 103402 -5751
rect 103298 -9764 103402 -5817
rect 106518 -5751 106622 -5750
rect 106518 -5817 106519 -5751
rect 106621 -5817 106622 -5751
rect 103298 -9858 103299 -9764
rect 103401 -9858 103402 -9764
rect 103298 -9859 103402 -9858
rect 106278 -7169 106382 -7168
rect 106278 -7235 106279 -7169
rect 106381 -7235 106382 -7169
rect 106278 -11168 106382 -7235
rect 106518 -9920 106622 -5817
rect 109738 -6287 109842 -6286
rect 109738 -6353 109739 -6287
rect 109841 -6353 109842 -6287
rect 106518 -10014 106519 -9920
rect 106621 -10014 106622 -9920
rect 106518 -10015 106622 -10014
rect 109498 -7169 109602 -7168
rect 109498 -7235 109499 -7169
rect 109601 -7235 109602 -7169
rect 109498 -11012 109602 -7235
rect 109738 -10076 109842 -6353
rect 109738 -10170 109739 -10076
rect 109841 -10170 109842 -10076
rect 109738 -10171 109842 -10170
rect 112958 -6287 113062 -6286
rect 112958 -6353 112959 -6287
rect 113061 -6353 113062 -6287
rect 112958 -10232 113062 -6353
rect 112958 -10326 112959 -10232
rect 113061 -10326 113062 -10232
rect 112958 -10327 113062 -10326
rect 116178 -7359 116282 -7358
rect 116178 -7425 116179 -7359
rect 116281 -7425 116282 -7359
rect 116178 -10388 116282 -7425
rect 116178 -10482 116179 -10388
rect 116281 -10482 116282 -10388
rect 116178 -10483 116282 -10482
rect 119398 -7359 119502 -7358
rect 119398 -7425 119399 -7359
rect 119501 -7425 119502 -7359
rect 119158 -10544 119262 -10543
rect 119158 -10638 119159 -10544
rect 119261 -10638 119262 -10544
rect 115938 -10700 116042 -10699
rect 115938 -10794 115939 -10700
rect 116041 -10794 116042 -10700
rect 109498 -11106 109499 -11012
rect 109601 -11106 109602 -11012
rect 109498 -11107 109602 -11106
rect 112718 -10856 112822 -10855
rect 112718 -10950 112719 -10856
rect 112821 -10950 112822 -10856
rect 106278 -11262 106279 -11168
rect 106381 -11262 106382 -11168
rect 106278 -11263 106382 -11262
rect 112718 -12529 112822 -10950
rect 112718 -12595 112719 -12529
rect 112821 -12595 112822 -12529
rect 112718 -12596 112822 -12595
rect 115938 -12529 116042 -10794
rect 115938 -12595 115939 -12529
rect 116041 -12595 116042 -12529
rect 115938 -12596 116042 -12595
rect 119158 -13601 119262 -10638
rect 119398 -10544 119502 -7425
rect 122618 -8431 122722 -8430
rect 122618 -8497 122619 -8431
rect 122721 -8497 122722 -8431
rect 119398 -10638 119399 -10544
rect 119501 -10638 119502 -10544
rect 119398 -10639 119502 -10638
rect 122378 -10388 122482 -10387
rect 122378 -10482 122379 -10388
rect 122481 -10482 122482 -10388
rect 119158 -13667 119159 -13601
rect 119261 -13667 119262 -13601
rect 119158 -13668 119262 -13667
rect 122378 -13601 122482 -10482
rect 122618 -10700 122722 -8497
rect 125838 -8431 125942 -8430
rect 125838 -8497 125839 -8431
rect 125941 -8497 125942 -8431
rect 122618 -10794 122619 -10700
rect 122721 -10794 122722 -10700
rect 122618 -10795 122722 -10794
rect 125598 -10232 125702 -10231
rect 125598 -10326 125599 -10232
rect 125701 -10326 125702 -10232
rect 122378 -13667 122379 -13601
rect 122481 -13667 122482 -13601
rect 122378 -13668 122482 -13667
rect 125598 -14673 125702 -10326
rect 125838 -10856 125942 -8497
rect 135258 -9764 135362 -9763
rect 135258 -9858 135259 -9764
rect 135361 -9858 135362 -9764
rect 132038 -9920 132142 -9919
rect 132038 -10014 132039 -9920
rect 132141 -10014 132142 -9920
rect 125838 -10950 125839 -10856
rect 125941 -10950 125942 -10856
rect 125838 -10951 125942 -10950
rect 128818 -10076 128922 -10075
rect 128818 -10170 128819 -10076
rect 128921 -10170 128922 -10076
rect 125598 -14739 125599 -14673
rect 125701 -14739 125702 -14673
rect 125598 -14740 125702 -14739
rect 128818 -14673 128922 -10170
rect 129058 -11012 129162 -11011
rect 129058 -11106 129059 -11012
rect 129161 -11106 129162 -11012
rect 129058 -13791 129162 -11106
rect 129058 -13857 129059 -13791
rect 129161 -13857 129162 -13791
rect 129058 -13858 129162 -13857
rect 128818 -14739 128819 -14673
rect 128921 -14739 128922 -14673
rect 128818 -14740 128922 -14739
rect 132038 -15209 132142 -10014
rect 132278 -11168 132382 -11167
rect 132278 -11262 132279 -11168
rect 132381 -11262 132382 -11168
rect 132278 -13791 132382 -11262
rect 132278 -13857 132279 -13791
rect 132381 -13857 132382 -13791
rect 132278 -13858 132382 -13857
rect 132038 -15275 132039 -15209
rect 132141 -15275 132142 -15209
rect 132038 -15276 132142 -15275
rect 135258 -15209 135362 -9858
rect 135258 -15275 135259 -15209
rect 135361 -15275 135362 -15209
rect 135258 -15276 135362 -15275
use x10b_cap_array  x10b_cap_array_0
timestamp 1730625751
transform -1 0 121209 0 -1 -40052
box -14221 -23088 17979 850
use x10b_cap_array  x10b_cap_array_1
timestamp 1730625751
transform 1 0 117451 0 1 19026
box -14221 -23088 17979 850
use cdac_sw_1  cdac_sw_1_0
timestamp 1730626724
transform 1 0 132149 0 1 -11152
box 23 -5764 3319 -3508
use cdac_sw_1  cdac_sw_1_1
timestamp 1730626724
transform 1 0 128929 0 1 -11152
box 23 -5764 3319 -3508
use cdac_sw_1  cdac_sw_1_2
timestamp 1730626724
transform -1 0 106511 0 -1 -9874
box 23 -5764 3319 -3508
use cdac_sw_2  cdac_sw_2_0
timestamp 1730626724
transform 1 0 125710 0 1 -11152
box 22 -5764 3318 -2972
use cdac_sw_2  cdac_sw_2_1
timestamp 1730626724
transform 1 0 122490 0 1 -11152
box 22 -5764 3318 -2972
use cdac_sw_4  cdac_sw_4_0
timestamp 1730626724
transform 1 0 119038 0 1 -11239
box 254 -5677 3550 -1813
use cdac_sw_4  cdac_sw_4_1
timestamp 1730626724
transform 1 0 115818 0 1 -11239
box 254 -5677 3550 -1813
use cdac_sw_8  cdac_sw_8_0
timestamp 1730626724
transform 1 0 112829 0 1 -11460
box 23 -5456 3319 552
use cdac_sw_8  cdac_sw_8_1
timestamp 1730626724
transform 1 0 109609 0 1 -11460
box 23 -5456 3319 552
use cdac_sw_16  cdac_sw_16_0
timestamp 1730626724
transform 1 0 103754 0 1 -14133
box -562 -2783 2734 7513
use cdac_sw_16  x2[0]
timestamp 1730626724
transform 1 0 106974 0 1 -14133
box -562 -2783 2734 7513
use cdac_sw_16  x3[0]
timestamp 1730626724
transform -1 0 134906 0 -1 -6893
box -562 -2783 2734 7513
use cdac_sw_16  x3[1]
timestamp 1730626724
transform -1 0 131686 0 -1 -6893
box -562 -2783 2734 7513
use cdac_sw_8  x4[2]
timestamp 1730626724
transform -1 0 129051 0 -1 -9566
box 23 -5456 3319 552
use cdac_sw_8  x4[3]
timestamp 1730626724
transform -1 0 125831 0 -1 -9566
box 23 -5456 3319 552
use cdac_sw_4  x6[4]
timestamp 1730626724
transform -1 0 122842 0 -1 -9787
box 254 -5677 3550 -1813
use cdac_sw_4  x6[5]
timestamp 1730626724
transform -1 0 119622 0 -1 -9787
box 254 -5677 3550 -1813
use cdac_sw_2  x8[6]
timestamp 1730626724
transform -1 0 116170 0 -1 -9874
box 22 -5764 3318 -2972
use cdac_sw_2  x8[7]
timestamp 1730626724
transform -1 0 112950 0 -1 -9874
box 22 -5764 3318 -2972
use cdac_sw_1  x10[8]
timestamp 1730626724
transform -1 0 109731 0 -1 -9874
box 23 -5764 3319 -3508
<< labels >>
flabel metal3 102622 -9859 102718 -9763 0 FreeSans 800 0 0 0 cf[9]
port 11 nsew
flabel metal3 102622 -10015 102718 -9919 0 FreeSans 800 0 0 0 cf[8]
port 10 nsew
flabel metal3 102622 -10171 102718 -10075 0 FreeSans 800 0 0 0 cf[7]
port 9 nsew
flabel metal3 102622 -10327 102718 -10231 0 FreeSans 800 0 0 0 cf[6]
port 8 nsew
flabel metal3 102622 -10483 102718 -10387 0 FreeSans 800 0 0 0 cf[5]
port 7 nsew
flabel metal3 102622 -10639 102718 -10543 0 FreeSans 800 0 0 0 cf[4]
port 6 nsew
flabel metal3 102622 -10795 102718 -10699 0 FreeSans 800 0 0 0 cf[3]
port 5 nsew
flabel metal3 102622 -10951 102718 -10855 0 FreeSans 800 0 0 0 cf[2]
port 4 nsew
flabel metal3 102622 -11107 102718 -11011 0 FreeSans 800 0 0 0 cf[1]
port 3 nsew
flabel metal3 102622 -11263 102718 -11167 0 FreeSans 800 0 0 0 cf[0]
port 2 nsew
flabel metal3 102622 -5628 102718 -5532 0 FreeSans 800 0 0 0 swp_in[9]
port 21 nsew
flabel metal3 102622 -5472 102718 -5376 0 FreeSans 800 0 0 0 swp_in[8]
port 20 nsew
flabel metal3 102622 -5316 102718 -5220 0 FreeSans 800 0 0 0 swp_in[7]
port 19 nsew
flabel metal3 102622 -5160 102718 -5064 0 FreeSans 800 0 0 0 swp_in[6]
port 18 nsew
flabel metal3 102622 -5004 102718 -4908 0 FreeSans 800 0 0 0 swp_in[5]
port 17 nsew
flabel metal3 102622 -4848 102718 -4752 0 FreeSans 800 0 0 0 swp_in[4]
port 16 nsew
flabel metal3 102622 -4692 102718 -4596 0 FreeSans 800 0 0 0 swp_in[3]
port 15 nsew
flabel metal3 102622 -4536 102718 -4440 0 FreeSans 800 0 0 0 swp_in[2]
port 14 nsew
flabel metal3 102622 -4380 102718 -4284 0 FreeSans 800 0 0 0 swp_in[1]
port 13 nsew
flabel metal3 102622 -4224 102718 -4128 0 FreeSans 800 0 0 0 swp_in[0]
port 12 nsew
flabel metal3 102622 -15494 102718 -15398 0 FreeSans 800 0 0 0 swn_in[9]
port 31 nsew
flabel metal3 102622 -15650 102718 -15554 0 FreeSans 800 0 0 0 swn_in[8]
port 30 nsew
flabel metal3 102622 -15806 102718 -15710 0 FreeSans 800 0 0 0 swn_in[7]
port 29 nsew
flabel metal3 102622 -15962 102718 -15866 0 FreeSans 800 0 0 0 swn_in[6]
port 28 nsew
flabel metal3 102622 -16118 102718 -16022 0 FreeSans 800 0 0 0 swn_in[5]
port 27 nsew
flabel metal3 102622 -16274 102718 -16178 0 FreeSans 800 0 0 0 swn_in[4]
port 26 nsew
flabel metal3 102622 -16430 102718 -16334 0 FreeSans 800 0 0 0 swn_in[3]
port 25 nsew
flabel metal3 102622 -16586 102718 -16490 0 FreeSans 800 0 0 0 swn_in[2]
port 24 nsew
flabel metal3 102622 -16742 102718 -16646 0 FreeSans 800 0 0 0 swn_in[1]
port 23 nsew
flabel metal3 102622 -16898 102718 -16802 0 FreeSans 800 0 0 0 swn_in[0]
port 22 nsew
flabel metal2 103046 19692 103230 19876 0 FreeSans 800 0 0 0 vdref
port 1 nsew
flabel metal2 102834 19692 103018 19876 0 FreeSans 800 0 0 0 vsref
port 33 nsew
flabel metal2 102622 19692 102806 19876 0 FreeSans 800 0 0 0 vcm
port 32 nsew
flabel metal2 119628 19692 119812 19876 0 FreeSans 800 0 0 0 vcp
port 34 nsew
flabel metal2 118848 -40901 119032 -40717 0 FreeSans 800 0 0 0 vcn
port 35 nsew
<< end >>
