magic
tech sky130A
magscale 1 2
timestamp 1731002366
<< dnwell >>
rect 773 -6771 3975 -981
rect 5554 -3232 6996 -1488
rect 5554 -6258 6996 -4516
<< nwell >>
rect 1104 -2087 1162 -2021
rect 1231 -2134 1245 -1993
rect 6056 -2088 6122 -2032
rect 6372 -2088 6438 -2032
rect 1027 -2734 1079 -2146
rect 1187 -2192 1245 -2134
rect 1231 -2678 1245 -2192
rect 6056 -2826 6122 -2770
rect 6372 -2826 6438 -2770
rect 6056 -4984 6122 -4928
rect 6372 -4984 6438 -4928
rect 1027 -5024 1079 -5018
rect 1021 -5612 1079 -5024
rect 1100 -5721 1166 -5665
rect 1107 -5723 1159 -5721
rect 6056 -5722 6122 -5666
rect 6372 -5722 6438 -5666
<< pwell >>
rect 1969 -3401 2429 -3349
rect 2357 -3487 2435 -3441
rect 1207 -3661 1245 -3519
rect 1187 -3719 1245 -3661
rect 1308 -3723 1422 -3515
rect 1969 -3564 2021 -3558
rect 1470 -3719 1744 -3615
rect 1969 -3719 2027 -3564
rect 2102 -3719 2376 -3615
rect 1975 -3725 2027 -3719
rect 922 -3802 1166 -3750
rect 1100 -3949 1166 -3945
rect 922 -4001 1166 -3949
rect 1423 -3995 1475 -3768
rect 2371 -3908 2423 -3850
rect 1732 -4001 1798 -3945
rect 2048 -4002 2114 -3945
rect 1187 -4078 1239 -4030
rect 1308 -4237 1422 -4029
rect 1783 -4181 1835 -4175
rect 922 -4309 998 -4291
rect 992 -4401 998 -4309
rect 2049 -4323 2113 -4271
rect 2358 -4311 2436 -4265
rect 2684 -4376 2742 -4266
rect 922 -4419 998 -4401
rect 2924 -4443 3047 -3309
<< ndiff >>
rect 1783 -4181 1835 -4175
<< poly >>
rect 6056 -2088 6122 -2032
rect 6372 -2088 6438 -2032
rect 6056 -2826 6122 -2770
rect 6372 -2826 6438 -2770
rect 6056 -4984 6122 -4928
rect 6372 -4984 6438 -4928
rect 6056 -5722 6122 -5666
rect 6372 -5722 6438 -5666
<< locali >>
rect 6056 -2088 6122 -2032
rect 6372 -2088 6438 -2032
rect 958 -2732 1087 -2124
rect 6056 -2826 6122 -2770
rect 6372 -2826 6438 -2770
rect 1308 -3723 1422 -3515
rect 2424 -3723 2572 -3515
rect 1308 -4237 1422 -4029
rect 2424 -4237 2572 -4029
rect 6056 -4984 6122 -4928
rect 6372 -4984 6438 -4928
rect 973 -5627 1102 -5019
rect 6056 -5722 6122 -5666
rect 6372 -5722 6438 -5666
<< viali >>
rect 6230 -2717 6264 -2141
rect 958 -3449 992 -3345
rect 958 -4407 992 -4303
rect 6230 -5613 6264 -5037
<< metal1 >>
rect 893 -987 7052 -981
rect 893 -1079 1027 -987
rect 1079 -1079 2055 -987
rect 2107 -1079 7052 -987
rect 893 -1085 7052 -1079
rect 5498 -1523 5602 -1085
rect 5488 -1627 5498 -1523
rect 5602 -1627 5612 -1523
rect 1190 -1880 6797 -1825
rect 1104 -2028 1162 -2021
rect 1104 -2080 1107 -2028
rect 1159 -2080 1162 -2028
rect 1104 -2087 1162 -2080
rect 1190 -2140 1245 -1880
rect 6056 -1977 6616 -1910
rect 6056 -2017 6123 -1977
rect 1021 -2728 1027 -2140
rect 1239 -2728 1245 -2140
rect 2606 -2084 6123 -2017
rect 1101 -2827 1107 -2775
rect 1159 -2827 1165 -2775
rect 1181 -3270 1187 -3218
rect 1239 -3270 1783 -3218
rect 1835 -3270 1841 -3218
rect 2606 -3298 2673 -2084
rect 6056 -2087 6123 -2084
rect 6056 -2088 6122 -2087
rect 6372 -2088 6438 -2032
rect 6224 -2141 6270 -2129
rect 6116 -2375 6230 -2141
rect 6264 -2375 6378 -2141
rect 5488 -2481 5498 -2377
rect 5602 -2481 6062 -2377
rect 6116 -2479 6195 -2375
rect 6299 -2479 6378 -2375
rect 6549 -2395 6616 -1977
rect 6432 -2462 6616 -2395
rect 6116 -2717 6230 -2479
rect 6264 -2717 6378 -2479
rect 6224 -2729 6270 -2717
rect 6742 -2764 6797 -1880
rect 6056 -2826 6122 -2770
rect 6371 -2819 6797 -2764
rect 6372 -2826 6438 -2819
rect 3182 -3271 3242 -3263
rect 922 -3345 1004 -3333
rect 922 -3449 958 -3345
rect 992 -3449 1004 -3345
rect 1739 -3401 2742 -3298
rect 922 -3462 1004 -3449
rect 1101 -3481 1107 -3429
rect 1159 -3481 1165 -3429
rect 1416 -3487 1482 -3431
rect 1739 -3481 1791 -3401
rect 1917 -3519 2021 -3401
rect 2049 -3481 2055 -3429
rect 2107 -3481 2113 -3429
rect 2357 -3487 2435 -3441
rect 2690 -3481 2742 -3401
rect 3182 -3456 3188 -3271
rect 3240 -3456 3242 -3271
rect 3182 -3463 3242 -3456
rect 1021 -3713 1027 -3519
rect 1079 -3713 1112 -3519
rect 1239 -3713 1245 -3519
rect 1187 -3719 1245 -3713
rect 1470 -3713 1578 -3519
rect 1630 -3713 1744 -3519
rect 1777 -3571 1783 -3519
rect 1835 -3571 1841 -3519
rect 1470 -3719 1744 -3713
rect 1917 -3719 2027 -3519
rect 2102 -3719 2376 -3519
rect 2637 -3531 2701 -3522
rect 2637 -3716 2701 -3707
rect 2734 -3719 3237 -3519
rect 3349 -3719 3852 -3519
rect 922 -3753 1166 -3750
rect 922 -3802 1107 -3753
rect 1100 -3805 1107 -3802
rect 1159 -3805 1166 -3753
rect 1100 -3807 1166 -3805
rect 1417 -3809 1481 -3757
rect 1732 -3807 1798 -3751
rect 2048 -3753 2114 -3751
rect 2048 -3805 2055 -3753
rect 2107 -3805 2114 -3753
rect 2370 -3760 2424 -3757
rect 2048 -3807 2114 -3805
rect 1423 -3850 1475 -3809
rect 2371 -3850 2423 -3760
rect 2680 -3799 3343 -3747
rect 922 -3902 2423 -3850
rect 1423 -3943 1475 -3902
rect 1100 -3949 1166 -3945
rect 922 -4001 1107 -3949
rect 1159 -4001 1166 -3949
rect 1417 -3995 1481 -3943
rect 1732 -4001 1798 -3945
rect 2048 -3950 2114 -3945
rect 2048 -4002 2055 -3950
rect 2107 -4002 2114 -3950
rect 2371 -3978 2423 -3902
rect 2680 -4005 3343 -3953
rect 1470 -4036 1744 -4033
rect 1021 -4233 1027 -4039
rect 1239 -4230 1245 -4036
rect 1470 -4230 1581 -4036
rect 1633 -4230 1744 -4036
rect 1470 -4233 1744 -4230
rect 1777 -4233 1783 -4181
rect 1835 -4233 1841 -4181
rect 922 -4303 998 -4291
rect 922 -4407 958 -4303
rect 992 -4407 998 -4303
rect 1101 -4323 1107 -4271
rect 1159 -4323 1165 -4271
rect 1416 -4321 1482 -4265
rect 922 -4419 998 -4407
rect 1736 -4355 1794 -4265
rect 1916 -4355 2020 -4033
rect 2102 -4137 2377 -4033
rect 2103 -4233 2377 -4137
rect 2637 -4045 2701 -4036
rect 2637 -4230 2701 -4221
rect 2734 -4233 3237 -4033
rect 3349 -4233 3852 -4033
rect 2048 -4305 2055 -4271
rect 2049 -4323 2055 -4305
rect 2107 -4323 2113 -4271
rect 2358 -4311 2436 -4265
rect 2684 -4355 2742 -4266
rect 1736 -4458 2742 -4355
rect 3179 -4296 3243 -4289
rect 1181 -4538 1187 -4486
rect 1239 -4538 1783 -4486
rect 1835 -4538 1841 -4486
rect 1101 -4977 1107 -4925
rect 1159 -4977 1165 -4925
rect 1021 -5612 1027 -5024
rect 1239 -5617 1252 -5029
rect 1100 -5717 1107 -5665
rect 1159 -5717 1166 -5665
rect 1100 -5721 1166 -5717
rect 1200 -5875 1252 -5617
rect 2605 -5681 2671 -4458
rect 3179 -4481 3186 -4296
rect 3238 -4481 3243 -4296
rect 3179 -4489 3243 -4481
rect 6056 -4984 6122 -4928
rect 6372 -4935 6438 -4928
rect 6372 -4987 6796 -4935
rect 6224 -5037 6270 -5025
rect 6116 -5273 6230 -5037
rect 6264 -5273 6378 -5037
rect 5492 -5378 5502 -5274
rect 5606 -5378 6062 -5274
rect 6116 -5377 6196 -5273
rect 6300 -5377 6378 -5273
rect 6432 -5358 6613 -5292
rect 6116 -5613 6230 -5377
rect 6264 -5613 6378 -5377
rect 6224 -5625 6270 -5613
rect 3243 -5681 3345 -5663
rect 6056 -5681 6122 -5666
rect 2605 -5747 6122 -5681
rect 6372 -5722 6438 -5666
rect 6056 -5775 6122 -5747
rect 6547 -5775 6613 -5358
rect 6056 -5841 6613 -5775
rect 6744 -5875 6796 -4987
rect 1200 -5927 6796 -5875
rect 5492 -6224 5502 -6120
rect 5606 -6224 5616 -6120
rect 5502 -6667 5606 -6224
rect 893 -6673 7046 -6667
rect 893 -6765 1027 -6673
rect 1079 -6765 2055 -6673
rect 2107 -6765 7046 -6673
rect 893 -6771 7046 -6765
<< via1 >>
rect 1027 -1079 1079 -987
rect 2055 -1079 2107 -987
rect 5498 -1627 5602 -1523
rect 1107 -2080 1159 -2028
rect 1027 -2728 1079 -2140
rect 1187 -2728 1239 -2140
rect 1107 -2827 1159 -2775
rect 1187 -3270 1239 -3218
rect 1783 -3270 1835 -3218
rect 5498 -2481 5602 -2377
rect 6195 -2479 6230 -2375
rect 6230 -2479 6264 -2375
rect 6264 -2479 6299 -2375
rect 1107 -3481 1159 -3429
rect 2055 -3481 2107 -3429
rect 3188 -3456 3240 -3271
rect 1027 -3713 1079 -3519
rect 1187 -3713 1239 -3519
rect 1578 -3713 1630 -3519
rect 1783 -3571 1835 -3519
rect 2637 -3707 2701 -3531
rect 1107 -3805 1159 -3753
rect 2055 -3805 2107 -3753
rect 1107 -4001 1159 -3949
rect 2055 -4002 2107 -3950
rect 1027 -4233 1079 -4039
rect 1187 -4230 1239 -4036
rect 1581 -4230 1633 -4036
rect 1783 -4233 1835 -4181
rect 1107 -4323 1159 -4271
rect 2637 -4221 2701 -4045
rect 2055 -4323 2107 -4271
rect 1187 -4538 1239 -4486
rect 1783 -4538 1835 -4486
rect 1107 -4977 1159 -4925
rect 1027 -5612 1079 -5024
rect 1187 -5617 1239 -5029
rect 1107 -5717 1159 -5665
rect 3186 -4481 3238 -4296
rect 5502 -5378 5606 -5274
rect 6196 -5377 6230 -5273
rect 6230 -5377 6264 -5273
rect 6264 -5377 6300 -5273
rect 5502 -6224 5606 -6120
rect 1027 -6765 1079 -6673
rect 2055 -6765 2107 -6673
<< metal2 >>
rect 1027 -987 1079 -981
rect 1027 -2140 1079 -1079
rect 2055 -987 2107 -981
rect 1027 -2734 1079 -2728
rect 1107 -2028 1159 -2022
rect 1107 -2775 1159 -2080
rect 1023 -3079 1079 -3070
rect 1023 -3192 1079 -3183
rect 1027 -3519 1079 -3192
rect 1027 -3719 1079 -3713
rect 1107 -3429 1159 -2827
rect 1107 -3753 1159 -3481
rect 1187 -2140 1239 -2134
rect 1187 -3218 1239 -2728
rect 1576 -3079 1632 -3070
rect 1576 -3192 1632 -3183
rect 1187 -3519 1239 -3270
rect 1187 -3719 1239 -3713
rect 1578 -3519 1630 -3192
rect 1783 -3218 1835 -3212
rect 1783 -3519 1835 -3270
rect 1783 -3577 1835 -3571
rect 2055 -3429 2107 -1079
rect 3861 -1325 3965 -1315
rect 3965 -1429 6299 -1325
rect 3861 -1438 3965 -1429
rect 5498 -1523 5602 -1513
rect 5498 -2377 5602 -1627
rect 5498 -2491 5602 -2481
rect 6195 -2375 6299 -1429
rect 6195 -2489 6299 -2479
rect 3185 -3271 3852 -3263
rect 3185 -3456 3188 -3271
rect 3240 -3456 3852 -3271
rect 3185 -3463 3852 -3456
rect 1578 -3719 1630 -3713
rect 1107 -3949 1159 -3805
rect 1027 -4039 1079 -4033
rect 1027 -4564 1079 -4233
rect 1022 -4573 1079 -4564
rect 1078 -4677 1079 -4573
rect 1022 -4686 1079 -4677
rect 1107 -4271 1159 -4001
rect 2055 -3753 2107 -3481
rect 2637 -3531 2701 -3522
rect 2637 -3716 2701 -3707
rect 2055 -3950 2107 -3805
rect 1107 -4925 1159 -4323
rect 1027 -5024 1079 -5018
rect 1027 -6673 1079 -5612
rect 1107 -5665 1159 -4977
rect 1187 -4036 1239 -4030
rect 1187 -4486 1239 -4230
rect 1187 -5029 1239 -4538
rect 1581 -4036 1633 -4030
rect 1581 -4564 1633 -4230
rect 1783 -4181 1835 -4175
rect 1783 -4486 1835 -4233
rect 1783 -4544 1835 -4538
rect 2055 -4271 2107 -4002
rect 2637 -4045 2701 -4036
rect 2637 -4230 2701 -4221
rect 1569 -4573 1644 -4564
rect 1569 -4677 1579 -4573
rect 1635 -4677 1644 -4573
rect 1569 -4687 1644 -4677
rect 1187 -5624 1239 -5617
rect 1107 -5723 1159 -5717
rect 1027 -6771 1079 -6765
rect 2055 -6673 2107 -4323
rect 3185 -4296 3852 -4289
rect 3185 -4481 3186 -4296
rect 3238 -4481 3852 -4296
rect 3185 -4489 3852 -4481
rect 5502 -5274 5606 -5264
rect 5502 -6120 5606 -5378
rect 5502 -6234 5606 -6224
rect 6196 -5273 6300 -5263
rect 3861 -6323 3965 -6314
rect 6196 -6323 6300 -5377
rect 3965 -6427 6300 -6323
rect 3861 -6437 3965 -6427
rect 2055 -6771 2107 -6765
<< via2 >>
rect 1023 -3183 1079 -3079
rect 1576 -3183 1632 -3079
rect 3861 -1429 3965 -1325
rect 1022 -4677 1078 -4573
rect 2637 -3707 2701 -3531
rect 2637 -4221 2701 -4045
rect 1579 -4677 1635 -4573
rect 3861 -6427 3965 -6323
<< metal3 >>
rect 3851 -1325 3975 -1320
rect 3851 -1429 3861 -1325
rect 3965 -1429 3975 -1325
rect 3851 -1434 3975 -1429
rect 2632 -3062 2709 -3056
rect 1018 -3079 1084 -3070
rect 1568 -3079 1638 -3070
rect 2632 -3079 2638 -3062
rect 1018 -3183 1023 -3079
rect 1079 -3183 1576 -3079
rect 1632 -3183 2638 -3079
rect 2703 -3183 2709 -3062
rect 1018 -3188 1084 -3183
rect 1568 -3189 1638 -3183
rect 2632 -3189 2709 -3183
rect 2632 -3531 2706 -3522
rect 2632 -3707 2637 -3531
rect 2701 -3707 2706 -3531
rect 2632 -3716 2706 -3707
rect 2628 -4045 2710 -4036
rect 2628 -4221 2637 -4045
rect 2701 -4221 2710 -4045
rect 2628 -4230 2710 -4221
rect 1017 -4573 1083 -4564
rect 1569 -4573 1644 -4564
rect 2630 -4565 2707 -4559
rect 2630 -4573 2636 -4565
rect 1017 -4677 1022 -4573
rect 1078 -4677 1579 -4573
rect 1635 -4677 2636 -4573
rect 1017 -4686 1083 -4677
rect 1569 -4687 1644 -4677
rect 2630 -4686 2636 -4677
rect 2701 -4686 2707 -4565
rect 2630 -4692 2707 -4686
rect 3851 -6323 3975 -6318
rect 3851 -6427 3861 -6323
rect 3965 -6427 3975 -6323
rect 3851 -6432 3975 -6427
<< via3 >>
rect 3861 -1429 3965 -1325
rect 2638 -3183 2703 -3062
rect 2637 -3707 2701 -3531
rect 2637 -4221 2701 -4045
rect 2636 -4686 2701 -4565
rect 3861 -6427 3965 -6323
<< metal4 >>
rect 3860 -1325 3966 -1324
rect 3653 -1429 3861 -1325
rect 3965 -1429 3966 -1325
rect 3860 -1430 3966 -1429
rect 2639 -3061 2699 -1807
rect 2637 -3062 2704 -3061
rect 2637 -3183 2638 -3062
rect 2703 -3183 2704 -3062
rect 2637 -3184 2704 -3183
rect 2639 -3530 2699 -3184
rect 2636 -3531 2702 -3530
rect 2636 -3707 2637 -3531
rect 2701 -3707 2702 -3531
rect 2636 -3708 2702 -3707
rect 2639 -3719 2699 -3708
rect 2636 -4045 2702 -4044
rect 2636 -4221 2637 -4045
rect 2701 -4221 2702 -4045
rect 2636 -4222 2702 -4221
rect 2639 -4564 2699 -4222
rect 2635 -4565 2702 -4564
rect 2635 -4686 2636 -4565
rect 2701 -4686 2702 -4565
rect 2635 -4687 2702 -4686
rect 2639 -5940 2699 -4687
rect 3860 -6323 3966 -6322
rect 3653 -6427 3861 -6323
rect 3965 -6427 3966 -6323
rect 3860 -6428 3966 -6427
use sky130_fd_pr__cap_mim_m3_1_V2UT89  XC1
timestamp 1730907816
transform 0 -1 2213 1 0 -6229
box -386 -1440 386 1440
use sky130_fd_pr__cap_mim_m3_1_V2UT89  XC2
timestamp 1730907816
transform 0 1 2213 -1 0 -1523
box -386 -1440 386 1440
use sky130_fd_pr__pfet_01v8_XGSNAL  XM1
timestamp 1730907816
transform 1 0 1133 0 1 -2428
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM2
timestamp 1730907816
transform 1 0 6089 0 1 -2429
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM3
timestamp 1730907816
transform 1 0 6405 0 1 -2429
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1730907816
transform 1 0 1133 0 1 -3619
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM5
timestamp 1730907816
transform 1 0 1449 0 1 -3619
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM6
timestamp 1730907816
transform 1 0 1765 0 1 -3619
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM7
timestamp 1730907816
transform 1 0 2081 0 1 -3619
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM8
timestamp 1730907816
transform 1 0 2397 0 1 -3619
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM9
timestamp 1730907816
transform 1 0 2713 0 1 -3619
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_RYGWKL  XM10
timestamp 1730907816
transform 1 0 3293 0 1 -2919
box -246 -1010 246 1010
use sky130_fd_pr__pfet_01v8_XGSNAL  XM11
timestamp 1730907816
transform 1 0 1133 0 1 -5324
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM12
timestamp 1730907816
transform 1 0 6089 0 1 -5325
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM13
timestamp 1730907816
transform 1 0 6405 0 1 -5325
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_648S5X  XM14
timestamp 1730907816
transform 1 0 1133 0 1 -4133
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM15
timestamp 1730907816
transform 1 0 1449 0 1 -4133
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM16
timestamp 1730907816
transform 1 0 1765 0 1 -4133
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM17
timestamp 1730907816
transform 1 0 2081 0 1 -4133
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM18
timestamp 1730907816
transform 1 0 2397 0 1 -4133
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM19
timestamp 1730907816
transform 1 0 2713 0 1 -4133
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_RYGWKL  XM20
timestamp 1730907816
transform 1 0 3293 0 1 -4833
box -246 -1010 246 1010
<< labels >>
flabel metal1 s 893 -1035 893 -1035 3 FreeSans 800 0 0 0 VDD
port 1 e
flabel metal2 s 3852 -3365 3852 -3365 7 FreeSans 800 0 0 0 VIP
port 4 w
flabel metal2 s 3852 -4386 3852 -4386 7 FreeSans 800 0 0 0 VIN
port 5 w
flabel metal1 s 922 -3402 922 -3402 3 FreeSans 800 0 0 0 VSS
port 6 e
flabel metal1 s 3852 -3624 3852 -3624 7 FreeSans 800 0 0 0 VCP
port 7 w
flabel metal1 s 3852 -4142 3852 -4142 7 FreeSans 800 0 0 0 VCN
port 8 w
flabel metal1 s 922 -3879 922 -3879 3 FreeSans 800 0 0 0 CLKSB
port 3 e
flabel metal1 s 922 -3780 922 -3780 3 FreeSans 800 0 0 0 CLKS
port 2 e
<< end >>
