* PEX produced on Sen 04 Nov 2024 06:58:17  CST using ./iic-pex.sh with m=1 and s=1
* NGSPICE file created from single_10b_cdac.ext - technology: sky130A

X0 cdac_sw_8_0.x2.swn cdac_sw_8_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 vdref cdac_sw_4_0.x1.x9.A cdac_sw_4_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 vsref cdac_sw_8_1.x1.x9.A cdac_sw_8_1.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 x6[4].x2.swn x6[4].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 cdac_sw_2_0.x1.x8.A cdac_sw_2_0.x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X10 x2[0].x2.swp x2[0].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 cdac_sw_2_0.x3.ck cdac_sw_2_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 vsref cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 a_122107_n4335# x6[4].x1.x8.A x6[4].x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 vdref x3[0].x1.x9.A x3[0].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 vdref x10[8].x1.x9.A x10[8].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 vsref x6[5].x1.x10.A x6[5].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 x3[1].x3.ckb x3[1].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 vdref x3[0].x3.ckb x3[0].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_116406_n15179# swn_in[4] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X25 x10b_cap_array_0.SW[5] cdac_sw_4_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X26 vdref cdac_sw_2_1.x3.ckb cdac_sw_2_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X27 cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 vdref x6[5].x2.swp x6[5].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 vcm cdac_sw_2_0.x2.swn x10b_cap_array_0.SW[7] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X36 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 vdref x6[4].x1.x10.A x6[4].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X41 a_115528_n6683# x8[6].x3.ckb x8[6].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X42 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X45 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 x6[5].x3.ckb x6[5].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X47 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X48 cdac_sw_8_1.x1.x5.A cdac_sw_8_1.x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X49 cdac_sw_4_0.x2.swp cdac_sw_4_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X50 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 vdref x6[4].x3.ckb x6[4].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X52 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 x6[4].dac_out x6[4].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X56 vdref cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X57 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 vdref x6[4].x1.x9.A x6[4].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X60 a_114650_n6256# swp_in[6] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X61 vsref cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X62 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 cdac_sw_1_1.x1.x8.A cdac_sw_1_1.x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X64 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 x4[3].x2.swp x4[3].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X66 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X71 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 x4[3].x3.ckb x4[3].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X73 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 vcp x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X77 x6[4].dac_out x6[4].x3.ck a_121090_n6892# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X78 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X79 vdref x8[7].x2.swp x8[7].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X80 vsref cdac_sw_2_0.x3.ckb cdac_sw_2_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X81 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X86 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 vdref x8[7].x1.x6.A x8[7].x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X90 vdref cdac_sw_8_1.x3.ckb cdac_sw_8_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X91 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 vcn x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 x6[5].x3.ckb x6[5].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X96 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 vdref x8[6].x1.x11.A x8[6].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X98 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X102 vdref cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X103 vdref cdac_sw_4_1.x1.x9.A cdac_sw_4_1.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X104 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 vdref cf[3] x4[3].x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X106 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X108 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 cdac_sw_1_2.x2.swn cdac_sw_1_2.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X112 vsref x4[3].x3.ckb x4[3].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X113 cdac_sw_1_0.x3.ck cdac_sw_1_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X114 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 x8[6].x1.x10.A x8[6].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X117 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 vsref x10[8].x1.x6.A x10[8].x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X121 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X122 vdref cdac_sw_1_1.x1.x8.A cdac_sw_1_1.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X123 vdref x6[5].x1.x10.A x6[5].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X124 cdac_sw_2_0.x3.ckb cdac_sw_2_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X125 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 a_128408_n9899# x4[2].x3.ckb x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X127 x10b_cap_array_0.SW[4] cdac_sw_4_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X128 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X129 cdac_sw_1_0.x2.swp cdac_sw_1_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X130 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 x6[5].x2.swn x6[5].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X132 cdac_sw_2_1.x1.x5.A cdac_sw_2_1.x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X133 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X136 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X137 vdref cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X138 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 x6[5].x3.ck x6[5].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X142 cdac_sw_2_0.x1.x3.Y cf[7] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X143 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 vsref cf[9] cdac_sw_1_2.x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X145 vdref x6[4].x1.x8.A x6[4].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X146 cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X147 cdac_sw_4_1.x1.x3.Y cf[4] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X148 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X151 vsref cdac_sw_8_0.x3.ckb cdac_sw_8_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X152 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X156 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X157 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 vdref cdac_sw_1_2.x3.ckb cdac_sw_1_2.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X159 x4[3].x2.swn x4[3].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X160 cdac_sw_1_2.x1.x5.A cdac_sw_1_2.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X161 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X162 vsref x2[0].x1.x10.A x2[0].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X163 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 cdac_sw_8_1.x3.ck cdac_sw_8_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X167 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 x4[3].x1.x11.A x4[3].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X170 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 vcn x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 vsref x6[5].x1.x5.A x6[5].x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X174 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X175 vsref cdac_sw_1_0.x1.x8.A cdac_sw_1_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X176 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X179 x10b_cap_array_0.SW[3] cdac_sw_8_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X180 cdac_sw_2_0.x1.x7.A cdac_sw_2_0.x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X181 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 cdac_sw_2_0.x1.x9.A cdac_sw_2_0.x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X184 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 x10[8].dac_out x10[8].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X188 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 vdref x8[6].x1.x8.A x8[6].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X191 vdref x2[0].x3.ckb x2[0].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X192 cdac_sw_8_0.x3.ckb cdac_sw_8_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X193 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X196 cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X197 cdac_sw_16_0.x3.ck cdac_sw_16_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X198 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 vdref x4[3].x3.ckb x4[3].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X201 vdref cdac_sw_2_1.x2.swp cdac_sw_2_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X202 cdac_sw_4_0.x2.swp cdac_sw_4_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X203 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 vsref x3[0].x3.ckb x3[0].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X205 x10[8].dac_out x10[8].x3.ck a_108210_n5938# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X206 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X207 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 x6[5].x1.x11.A x6[5].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X212 cdac_sw_8_0.x3.ck cdac_sw_8_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X213 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 vsref x6[4].x1.x10.A x6[4].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X217 vdref cdac_sw_2_0.x1.x8.A cdac_sw_2_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X218 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X219 cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X220 vsref x3[1].x1.x11.A x3[1].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X221 vsref x6[4].x3.ckb x6[4].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X222 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 a_110844_n15188# cdac_sw_8_1.x3.ck x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X225 vdref cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X226 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 vsref x6[4].x1.x9.A a_122107_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X229 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 vdref x6[4].x1.x5.A x6[4].x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X234 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 cdac_sw_4_1.x1.x5.A cdac_sw_4_1.x1.x8.A a_116499_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X236 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 vdref x8[6].x1.x10.A x8[6].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X238 cdac_sw_4_1.x3.ckb cdac_sw_4_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X239 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 x3[1].x2.swp x3[1].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X241 vsref swn_in[3] a_114064_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X242 x4[2].dac_out x4[2].x3.ck a_127530_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X243 cdac_sw_8_1.x1.x6.A cdac_sw_8_1.x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X244 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X246 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 x2[0].x3.ck x2[0].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X249 vsref cdac_sw_4_1.x1.x9.A cdac_sw_4_1.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X250 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 a_108210_n5938# swp_in[8] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X252 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 vsref x8[7].x1.x6.A x8[7].x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X255 vdref swp_in[4] a_121968_n7755# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X256 vdref cdac_sw_8_1.x2.swp cdac_sw_8_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X257 x6[5].x2.swp x6[5].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X258 vdref x6[4].x1.x10.A x6[4].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X259 vsref cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X260 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 x6[5].x3.ckb x6[5].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X262 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X263 vcm x6[5].x2.swp x6[5].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X264 x4[3].dac_out x4[3].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X265 x6[5].x2.swn x6[5].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X266 vdref cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X267 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 cdac_sw_1_0.x2.swn cdac_sw_1_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X276 cdac_sw_2_1.x2.swn cdac_sw_2_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X277 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 x4[3].x2.swp x4[3].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X282 x4[3].dac_out x4[3].x3.ck a_124310_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X283 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X284 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X285 vdref cdac_sw_1_1.x1.x9.A cdac_sw_1_1.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X286 vsref x6[5].x1.x10.A x6[5].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X287 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 x6[4].x3.ck x6[4].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X290 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X291 cdac_sw_2_0.x2.swp cdac_sw_2_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X292 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 cdac_sw_4_1.x2.swp cdac_sw_4_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X294 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X297 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X298 x6[4].x1.x4.A cf[4] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X299 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 vdref swp_in[3] a_125188_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X305 vsref x4[3].x1.x11.A x4[3].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X306 vsref x6[4].x1.x8.A x6[4].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X307 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X308 cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X309 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 vsref x6[4].x1.x7.A x6[4].x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X311 vdref cdac_sw_1_0.x3.ckb cdac_sw_1_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X312 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 x8[7].x2.swn x8[7].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X317 vsref cdac_sw_1_2.x3.ckb cdac_sw_1_2.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X318 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X320 vsref x4[3].x2.swp x4[3].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X321 cdac_sw_8_1.x2.swn cdac_sw_8_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X322 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 x6[4].x2.swp x6[4].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X325 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X328 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 vdref swp_in[3] a_125188_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X330 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X331 vdref cdac_sw_4_1.x3.ckb cdac_sw_4_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X332 x2[0].x1.x6.A x2[0].x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X333 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 a_124310_n8164# swp_in[3] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X335 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 vsref cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X338 x8[7].dac_out x8[7].x3.ck a_111430_n6256# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X339 x4[3].x3.ckb x4[3].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X340 vdref cdac_sw_8_1.x1.x8.A cdac_sw_8_1.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X341 vsref cdac_sw_2_1.x2.swp cdac_sw_2_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X342 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 vdref x8[6].x1.x11.A x8[6].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X346 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 vsref x8[6].x1.x8.A x8[6].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X348 cdac_sw_8_0.x2.swp cdac_sw_8_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X349 x6[5].x1.x11.A x6[5].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X350 vdref x2[0].x2.swp x2[0].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X351 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X353 vsref cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X354 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 cdac_sw_16_0.x2.swn cdac_sw_16_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X356 vsref x4[3].x3.ckb x4[3].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X357 a_103619_n16821# cdac_sw_16_0.x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X358 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 cdac_sw_16_0.x2.swn cdac_sw_16_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X360 vsref x6[5].x2.swp x6[5].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X361 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 vcm cdac_sw_8_1.x2.swn x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X368 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 vdref cdac_sw_2_0.x1.x9.A cdac_sw_2_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X373 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 x10b_cap_array_0.SW[3] cdac_sw_8_0.x3.ckb a_113186_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X375 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X377 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 vdref swp_in[6] a_115528_n6683# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X379 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 cdac_sw_1_2.x3.ck cdac_sw_1_2.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X381 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 x10b_cap_array_0.SW[2] cdac_sw_8_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X384 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X386 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 vsref x4[3].x1.x9.A x4[3].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X390 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X391 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 vsref x8[6].x1.x10.A x8[6].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X393 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 x6[5].x3.ck x6[5].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X395 vsref x3[0].x2.swp x3[0].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X396 vsref cdac_sw_8_1.x2.swp cdac_sw_8_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X397 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X399 x2[0].x1.x9.A x2[0].x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X400 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 x10b_cap_array_0.SW[4] cdac_sw_4_1.x3.ckb a_116406_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X407 x2[0].x2.swn x2[0].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 x6[4].x1.x11.A x6[4].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X410 vsref cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X411 vsref cdac_sw_2_1.x3.ckb cdac_sw_2_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X412 cdac_sw_1_1.x3.ckb cdac_sw_1_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X413 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 vdref x8[6].x1.x5.A x8[6].x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X415 x6[5].dac_out x6[5].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X416 vcm cdac_sw_8_0.x2.swn x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X417 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 a_121968_n7755# x6[4].x3.ckb x6[4].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X420 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 vsref x6[4].x1.x10.A x6[4].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X423 vcm cdac_sw_4_0.x2.swn x10b_cap_array_0.SW[5] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X424 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 x4[3].x3.ck x4[3].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X426 x10b_cap_array_0.SW[3] cdac_sw_8_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X427 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 vsref cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X429 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 cdac_sw_4_0.x3.ck cdac_sw_4_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X431 vsref cdac_sw_1_1.x1.x9.A cdac_sw_1_1.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X432 cdac_sw_8_0.x3.ckb cdac_sw_8_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X433 vdref x2[0].x1.x8.A x2[0].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X434 x4[3].x1.x10.A x4[3].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X435 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 vdref x6[5].x1.x4.A x6[5].x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X437 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X438 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 cdac_sw_4_1.x2.swn cdac_sw_4_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X440 vcm x4[3].x2.swp x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X441 vdref cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X442 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 vsref x4[3].x1.x11.A x4[3].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X445 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X446 vsref x4[2].x2.swp x4[2].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X447 x6[4].x3.ck x6[4].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X448 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X449 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X450 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 x8[6].x1.x11.A x8[6].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X453 cdac_sw_2_1.x3.ckb cdac_sw_2_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X454 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 a_122107_n5199# cf[4] x6[4].x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X456 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X457 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 vdref x3[0].x1.x7.A x3[0].x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X459 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 cdac_sw_2_1.x3.ck cdac_sw_2_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X463 vdref cdac_sw_1_0.x2.swp cdac_sw_1_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X464 x6[5].x2.swp x6[5].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X465 vsref x3[1].x1.x11.A x3[1].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X466 x6[5].dac_out x6[5].x3.ck a_117870_n6892# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X467 x4[2].dac_out x4[2].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X468 a_128408_n9899# x4[2].x3.ckb x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X469 cdac_sw_1_1.x2.swp cdac_sw_1_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X470 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 vcm x4[3].x2.swp x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X475 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 vsref x8[6].x1.x3.Y a_115667_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X477 x6[5].x1.x10.A x6[5].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X478 cdac_sw_4_1.x3.ckb cdac_sw_4_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X479 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 vdref x8[6].x1.x9.A x8[6].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X481 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X482 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 x3[1].x2.swp x3[1].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X484 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X485 cdac_sw_2_1.x3.ck cdac_sw_2_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X486 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X489 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 vdref x3[1].x1.x10.A x3[1].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X491 vdref swp_in[5] a_118748_n7755# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X492 a_117870_n6892# swp_in[5] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X493 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 vsref x6[5].x1.x11.A x6[5].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X496 vdref cdac_sw_4_1.x2.swp cdac_sw_4_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X497 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 vsref x8[6].x1.x7.A x8[6].x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X499 vsref x2[0].x2.swp x2[0].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X500 a_113186_n15179# swn_in[3] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X501 a_120504_n15188# cdac_sw_4_0.x3.ck x10b_cap_array_0.SW[5] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X502 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 vsref cdac_sw_16_0.x3.ckb cdac_sw_16_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X504 cdac_sw_16_0.x2.swn cdac_sw_16_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X505 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X507 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 x4[3].x3.ckb x4[3].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X510 vdref cdac_sw_8_1.x1.x9.A cdac_sw_8_1.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X511 cdac_sw_2_0.x1.x5.A cdac_sw_2_0.x1.x8.A a_126159_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X512 a_110844_n15188# cdac_sw_8_1.x3.ck x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X513 x3[1].x3.ckb x3[1].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X514 cdac_sw_2_0.x3.ckb cdac_sw_2_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X515 vdref cdac_sw_1_1.x3.ckb cdac_sw_1_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X516 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 x8[6].x2.swp x8[6].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X518 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 cdac_sw_4_0.x1.x6.A cdac_sw_4_0.x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X520 vcn vcm sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 vcm cdac_sw_4_1.x2.swn x10b_cap_array_0.SW[4] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X522 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 vdref x3[1].x2.swp x3[1].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X526 cdac_sw_4_1.x3.ck cdac_sw_4_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X527 vdref cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X528 vsref cdac_sw_2_0.x1.x9.A cdac_sw_2_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X529 vdref cdac_sw_8_0.x3.ckb cdac_sw_8_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X530 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X533 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 x6[5].x3.ckb x6[5].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X536 cdac_sw_8_1.x3.ck cdac_sw_8_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X537 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 a_125188_n9899# x4[3].x3.ckb x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X539 vsref cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X540 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 x6[4].x2.swp x6[4].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X543 vdref x2[0].x1.x10.A x2[0].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X544 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 a_127530_n8164# swp_in[2] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X548 cdac_sw_16_0.x3.ckb cdac_sw_16_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X549 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X551 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X554 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 cdac_sw_1_2.x3.ck cdac_sw_1_2.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X557 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 x4[3].x3.ckb x4[3].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X560 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 x10[8].x2.swp x10[8].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X564 cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X565 vdref x6[4].x1.x11.A x6[4].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X566 cdac_sw_4_0.x1.x4.A cdac_sw_4_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X567 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X569 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 vsref cdac_sw_1_0.x3.ckb cdac_sw_1_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X572 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 vsref cdac_sw_16_0.x2.swp cdac_sw_16_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X574 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X575 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X576 x6[5].x3.ck x6[5].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X577 a_116406_n15179# swn_in[4] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X578 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 vdref x6[4].x2.swp x6[4].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X581 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X582 cdac_sw_8_1.x1.x4.A cf[2] a_110059_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X583 vsref cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X584 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X585 vdref x4[3].x1.x10.A x4[3].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X586 a_126066_n15179# swn_in[7] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X587 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 vsref x4[2].x1.x11.A x4[2].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X589 vdref x10[8].x1.x11.A x10[8].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X590 vdref x6[4].x1.x6.A x6[4].x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X591 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 x8[6].x2.swp x8[6].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X593 cdac_sw_8_0.x3.ck cdac_sw_8_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X594 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 vcp x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 cdac_sw_4_0.x1.x9.A cdac_sw_4_0.x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X598 vdref cf[0] x3[0].x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X599 x4[3].x3.ck x4[3].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X600 vsref cdac_sw_2_1.x1.x9.A cdac_sw_2_1.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X601 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 vdref x10[8].x1.x3.Y x10[8].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X604 vdref x4[3].x3.ckb x4[3].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X605 x2[0].x3.ckb x2[0].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X606 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 vsref x4[2].x2.swp x4[2].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X608 cdac_sw_4_0.x2.swn cdac_sw_4_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X609 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 vsref cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X612 vdref x2[0].x1.x9.A x2[0].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X613 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 x4[3].x1.x10.A x4[3].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X616 x4[3].dac_out x4[3].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X617 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X618 vsref x6[5].x1.x4.A x6[5].x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X619 vdref cdac_sw_2_0.x3.ckb cdac_sw_2_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X620 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X622 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X624 x4[2].dac_out x4[2].x3.ck a_127530_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X625 vdref cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X626 cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X627 x4[2].x2.swn x4[2].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X628 vdref cdac_sw_4_0.x1.x8.A cdac_sw_4_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X629 x4[3].dac_out x4[3].x3.ck a_124310_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X630 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X631 vsref cdac_sw_1_0.x2.swp cdac_sw_1_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X632 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 vdref x8[6].x2.swp x8[6].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X634 cdac_sw_4_1.x3.ckb cdac_sw_4_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X635 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 cdac_sw_1_1.x2.swn cdac_sw_1_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X638 x6[5].x1.x10.A x6[5].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X639 cdac_sw_2_1.x2.swp cdac_sw_2_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X640 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X642 vsref cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X643 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 cdac_sw_2_1.x2.swn cdac_sw_2_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X645 a_113279_n16821# cdac_sw_8_0.x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X646 cdac_sw_2_1.x2.swp cdac_sw_2_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X647 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 vsref cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 vdref x6[5].x3.ckb x6[5].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X652 vdref x4[2].x1.x3.Y x4[2].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X653 vsref x6[4].x2.swp x6[4].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X654 x3[0].x2.swn x3[0].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X655 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X656 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 vsref cdac_sw_16_0.x3.ckb cdac_sw_16_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X658 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 x6[5].x1.x10.A x6[5].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X660 cdac_sw_4_1.x2.swp cdac_sw_4_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X661 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X667 vdref x6[4].x1.x9.A x6[4].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X668 vsref x4[2].x1.x5.A x4[2].x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X669 vdref x4[2].x1.x7.A x4[2].x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X670 a_118748_n7755# x6[5].x3.ckb x6[5].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X671 x10b_cap_array_0.SW[6] cdac_sw_2_1.x3.ckb a_122846_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X672 vsref x3[1].x1.x10.A x3[1].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X673 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 x6[4].x2.swn x6[4].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X675 cdac_sw_1_1.x3.ckb cdac_sw_1_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X676 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X678 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X680 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X681 vsref cdac_sw_2_1.x1.x8.A cdac_sw_2_1.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X682 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 vcp x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 vdref x10[8].x1.x9.A x10[8].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X685 vdref x4[3].x1.x8.A x4[3].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X686 a_124310_n8164# swp_in[3] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X687 vsref swn_in[3] a_114064_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X688 vsref cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X689 vsref x8[7].x1.x11.A x8[7].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X690 x3[1].x3.ckb x3[1].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X691 vdref cdac_sw_1_1.x2.swp cdac_sw_1_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X692 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 vdref x3[0].x3.ckb x3[0].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X694 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 x3[0].x1.x5.A x3[0].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X696 cdac_sw_4_1.x1.x9.A cdac_sw_4_1.x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X697 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X698 x4[2].x2.swn x4[2].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X699 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X700 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X701 cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X702 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 x10b_cap_array_0.SW[7] cdac_sw_2_0.x3.ckb a_126066_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X704 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X705 cdac_sw_4_1.x2.swn cdac_sw_4_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X706 vdref cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X707 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X709 vdref cdac_sw_8_0.x2.swp cdac_sw_8_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X710 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 vsref x8[7].x2.swp x8[7].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X713 cdac_sw_8_1.x2.swp cdac_sw_8_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X714 cdac_sw_8_1.x2.swn cdac_sw_8_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X715 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X716 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X717 x6[5].x3.ckb x6[5].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X718 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 x10b_cap_array_0.SW[6] cdac_sw_2_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X721 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 vdref x2[0].x1.x11.A x2[0].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X724 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 vdref x4[3].x2.swp x4[3].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X726 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 cdac_sw_16_0.x2.swp cdac_sw_16_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X728 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X730 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 x8[7].x2.swn x8[7].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X733 a_115667_n4335# x8[6].x1.x8.A x8[6].x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X734 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X735 cdac_sw_1_0.x3.ckb cdac_sw_1_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X736 cdac_sw_2_0.x2.swn cdac_sw_2_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X737 vsref cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X738 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X740 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X742 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 vdref x4[3].x1.x10.A x4[3].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X744 x4[3].x3.ckb x4[3].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X745 cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X746 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 vdref x4[2].x3.ckb x4[2].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X748 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X749 cdac_sw_4_0.x1.x5.A cdac_sw_4_0.x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X750 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 x4[3].x2.swn x4[3].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X752 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X753 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X756 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X757 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X758 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X759 vdref x8[7].x1.x3.Y x8[7].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X760 vsref cdac_sw_1_2.x2.swp cdac_sw_1_2.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X761 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X762 vsref x4[3].x1.x10.A x4[3].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X763 cdac_sw_1_0.x1.x4.A cdac_sw_1_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X764 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X767 vsref x6[4].x1.x6.A x6[4].x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X768 cdac_sw_1_0.x3.ck cdac_sw_1_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X769 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X770 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X771 x6[5].x3.ckb x6[5].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X772 vdref x3[1].x1.x10.A x3[1].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X773 x10b_cap_array_0.SW[3] cdac_sw_8_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X774 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 vdref x8[6].x1.x11.A x8[6].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X777 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 vsref x8[7].x1.x5.A x8[7].x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X779 a_125188_n9899# x4[3].x3.ckb x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X780 vsref cdac_sw_16_0.x1.x8.A cdac_sw_16_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X781 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 vdref x8[6].x1.x9.A x8[6].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X784 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X785 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X786 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X787 cdac_sw_1_0.x3.ck cdac_sw_1_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X788 vsref cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X789 vcn x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X790 cdac_sw_1_2.x2.swn cdac_sw_1_2.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X791 vsref x4[3].x3.ckb x4[3].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X792 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X793 vsref cdac_sw_1_1.x3.ckb cdac_sw_1_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X794 cdac_sw_1_1.x1.x9.A cdac_sw_1_1.x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X795 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X796 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X797 vdref x6[5].x1.x10.A x6[5].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X798 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X799 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X800 vdref x8[6].x1.x6.A x8[6].x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X801 x8[6].dac_out x8[6].x3.ck a_114650_n6256# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X802 vdref cdac_sw_2_0.x2.swp cdac_sw_2_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X803 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X804 vsref cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X805 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X806 cdac_sw_4_0.x3.ckb cdac_sw_4_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X807 cdac_sw_8_1.x1.x8.A cdac_sw_8_1.x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X808 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X809 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X810 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X811 cdac_sw_8_1.x3.ck cdac_sw_8_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X812 vsref cdac_sw_2_0.x2.swp cdac_sw_2_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X813 vdref cdac_sw_4_0.x1.x9.A cdac_sw_4_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X814 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X815 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X816 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X817 cdac_sw_4_1.x2.swp cdac_sw_4_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X818 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X819 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X820 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X821 x6[5].x1.x10.A x6[5].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X822 cdac_sw_16_0.x3.ckb cdac_sw_16_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X823 vsref x3[1].x1.x5.A x3[1].x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X824 vdref x10[8].x1.x11.A x10[8].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X825 vcm cdac_sw_2_0.x2.swn x10b_cap_array_0.SW[7] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X826 vdref cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X827 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X828 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X829 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X830 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X831 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X832 cdac_sw_1_1.x3.ckb cdac_sw_1_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X833 vsref x6[5].x3.ckb x6[5].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X834 vcm cdac_sw_8_1.x2.swn x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X835 cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X836 x4[2].dac_out x4[2].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X837 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X838 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X839 x6[4].dac_out x6[4].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X840 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X841 x4[2].x2.swp x4[2].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X842 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X843 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X844 vdref cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X845 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X846 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X847 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X848 x6[4].dac_out x6[4].x3.ck a_121090_n6892# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X849 cdac_sw_8_0.x1.x8.A cdac_sw_8_0.x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X850 cdac_sw_1_1.x2.swp cdac_sw_1_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X851 x10[8].x1.x5.A x10[8].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X852 vdref swp_in[4] a_121968_n7755# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X853 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X854 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X855 x4[2].x2.swn x4[2].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X856 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X857 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X858 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X859 x3[1].x1.x11.A x3[1].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X860 vdref x4[3].x1.x11.A x4[3].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X861 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X862 cdac_sw_1_1.x1.x4.A cdac_sw_1_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X863 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X864 vsref x4[3].x1.x8.A x4[3].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X865 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X866 vcm x6[5].x2.swp x6[5].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X867 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X868 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X869 vsref cdac_sw_8_0.x2.swp cdac_sw_8_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X870 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X871 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X872 vsref x3[0].x3.ckb x3[0].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X873 vsref cdac_sw_8_1.x3.ckb cdac_sw_8_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X874 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X875 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X876 vsref x4[2].x2.swp x4[2].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X877 vsref x2[0].x1.x11.A x2[0].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X878 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X879 vsref x3[1].x1.x9.A x3[1].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X880 vdref x4[2].x1.x10.A x4[2].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X881 cdac_sw_2_1.x3.ck cdac_sw_2_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X882 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X883 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X884 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X885 cdac_sw_4_1.x1.x6.A cdac_sw_4_1.x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X886 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X887 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X888 vsref cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X889 vsref cdac_sw_1_0.x1.x9.A cdac_sw_1_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X890 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X891 a_126944_n15188# cdac_sw_2_0.x3.ck x10b_cap_array_0.SW[7] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X892 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X893 vdref cdac_sw_4_0.x3.ckb cdac_sw_4_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X894 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X895 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X896 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X897 vdref x4[2].x3.ckb x4[2].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X898 vdref swp_in[3] a_125188_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X899 a_106839_n15957# x2[0].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X900 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X901 x4[3].x2.swn x4[3].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X902 x4[2].x1.x5.A x4[2].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X903 vsref cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X904 x6[4].x2.swn x6[4].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X905 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X906 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X907 a_127530_n8164# swp_in[2] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X908 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X909 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X910 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X911 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X912 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X913 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X914 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X915 vsref swn_in[5] a_120504_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X916 vdref cdac_sw_16_0.x3.ckb cdac_sw_16_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X917 cdac_sw_8_1.x3.ckb cdac_sw_8_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X918 cdac_sw_1_0.x3.ck cdac_sw_1_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X919 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X920 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X921 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X922 x3[1].x2.swp x3[1].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X923 cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X924 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X925 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X926 cdac_sw_1_2.x2.swp cdac_sw_1_2.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X927 vsref x4[3].x1.x10.A x4[3].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X928 x4[2].x3.ck x4[2].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X929 vsref x4[2].x3.ckb x4[2].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X930 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X931 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X932 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X933 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X934 cdac_sw_2_0.x3.ckb cdac_sw_2_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X935 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X936 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X937 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X938 cdac_sw_8_0.x2.swn cdac_sw_8_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X939 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X940 cdac_sw_1_0.x1.x5.A cdac_sw_1_0.x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X941 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X942 vdref x4[3].x1.x5.A x4[3].x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X943 cdac_sw_1_0.x2.swn cdac_sw_1_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X944 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X945 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X946 x8[7].x2.swp x8[7].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X947 x6[5].x3.ckb x6[5].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X948 vsref x3[1].x1.x10.A x3[1].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X949 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X950 vdref x6[4].x3.ckb x6[4].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X951 x3[0].x3.ck x3[0].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X952 vdref x2[0].x1.x10.A x2[0].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X953 x6[5].x2.swn x6[5].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X954 vsref x8[6].x1.x9.A a_115667_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X955 vdref cf[1] x2[0].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X956 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X957 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X958 vdref x4[2].x1.x4.A x4[2].x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X959 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X960 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X961 x4[3].x2.swp x4[3].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X962 cdac_sw_4_1.x2.swp cdac_sw_4_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X963 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X964 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X965 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X966 vsref x6[5].x1.x10.A x6[5].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X967 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X968 x6[4].x3.ck x6[4].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X969 vsref x8[6].x1.x6.A x8[6].x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X970 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X971 vsref x2[0].x3.ckb x2[0].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X972 cdac_sw_8_1.x1.x7.A cdac_sw_8_1.x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X973 vdref x6[5].x2.swp x6[5].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X974 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X975 x4[3].x2.swn x4[3].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X976 cdac_sw_8_1.x1.x9.A cdac_sw_8_1.x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X977 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X978 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X979 vsref swn_in[6] a_123724_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X980 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X981 vdref cdac_sw_1_0.x3.ckb cdac_sw_1_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X982 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X983 vsref x8[7].x2.swp x8[7].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X984 x4[3].x1.x11.A x4[3].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X985 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X986 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X987 vdref x8[7].x1.x10.A x8[7].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X988 x10b_cap_array_0.SW[3] cdac_sw_8_0.x3.ckb a_113186_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X989 x10b_cap_array_0.SW[4] cdac_sw_4_1.x3.ckb a_116406_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X990 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X991 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X992 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X993 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X994 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X995 vdref cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X996 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X997 x8[7].x2.swn x8[7].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X998 x4[2].x3.ck x4[2].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X999 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1000 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1001 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1002 vdref cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1003 x10b_cap_array_0.SW[2] cdac_sw_8_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1004 x10b_cap_array_0.SW[3] cdac_sw_8_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1005 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1006 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1007 vsref x4[3].x1.x3.Y a_125327_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1008 cdac_sw_8_0.x3.ck cdac_sw_8_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1009 cdac_sw_1_1.x2.swp cdac_sw_1_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1010 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1011 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1012 vdref x8[7].x3.ckb x8[7].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1013 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1014 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1015 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1016 x8[7].x1.x5.A x8[7].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1017 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1018 cdac_sw_1_2.x2.swn cdac_sw_1_2.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1019 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1020 vdref cdac_sw_8_1.x1.x8.A cdac_sw_8_1.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1021 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1022 vsref swn_in[4] a_117284_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1023 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1024 vcm cdac_sw_1_2.x2.swp cdac_sw_1_2.dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1025 x2[0].x3.ckb x2[0].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1026 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1027 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1028 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1029 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1030 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1031 vcn x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1032 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1033 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1034 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1035 vdref cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1036 x8[7].x3.ck x8[7].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1037 x8[6].x1.x4.A cf[6] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1038 x2[0].x1.x3.Y cf[1] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1039 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1040 vsref swn_in[3] a_114064_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1041 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1042 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1043 cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1044 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1045 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1046 a_121968_n7755# x6[4].x3.ckb x6[4].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1047 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1048 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1049 cdac_sw_1_1.x1.x5.A cdac_sw_1_1.x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1050 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1051 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1052 vdref cdac_sw_1_2.x3.ckb cdac_sw_1_2.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1053 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1054 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1055 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1056 vsref x4[2].x1.x10.A x4[2].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1057 vcm x4[3].x2.swp x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1058 cdac_sw_4_1.x3.ck cdac_sw_4_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1059 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1060 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1061 vdref x8[7].x1.x4.A x8[7].x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1062 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1063 vdref x6[5].x1.x11.A x6[5].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1064 x3[1].x2.swp x3[1].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1065 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1066 vsref cdac_sw_8_0.x1.x8.A cdac_sw_8_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1067 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1068 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1069 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1070 cdac_sw_4_1.x1.x7.A cdac_sw_4_1.x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1071 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1072 x2[0].x1.x7.A x2[0].x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1073 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1074 cdac_sw_1_2.x3.ck cdac_sw_1_2.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1075 vdref cdac_sw_4_0.x2.swp cdac_sw_4_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1076 vsref cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1077 vsref x4[2].x3.ckb x4[2].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1078 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1079 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1080 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1081 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1082 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1083 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1084 vsref x4[3].x1.x9.A x4[3].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1085 x6[5].x2.swp x6[5].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1086 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1087 vdref cdac_sw_16_0.x2.swp cdac_sw_16_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1088 cdac_sw_8_1.x2.swp cdac_sw_8_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1089 cdac_sw_1_0.x2.swn cdac_sw_1_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1090 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1091 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1092 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1093 x4[2].x3.ck x4[2].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1094 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1095 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1096 cdac_sw_2_0.x2.swp cdac_sw_2_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1097 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1098 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1099 vdref swp_in[5] a_118748_n7755# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1100 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1101 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1102 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1103 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1104 vdref x3[1].x1.x4.A x3[1].x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1105 x4[3].x2.swp x4[3].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1106 a_113186_n15179# swn_in[3] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1107 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1108 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1109 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1110 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1111 vdref x2[0].x1.x11.A x2[0].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1112 vsref x6[4].x3.ckb x6[4].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1113 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1114 x3[0].x3.ck x3[0].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1115 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1116 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1117 vdref x2[0].x1.x8.A x2[0].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1118 vsref x6[5].x1.x9.A x6[5].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1119 x4[2].x3.ckb x4[2].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1120 vdref swp_in[3] a_125188_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1121 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1122 vsref x4[2].x1.x4.A x4[2].x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1123 a_117284_n15188# cdac_sw_4_1.x3.ck x10b_cap_array_0.SW[4] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1124 cdac_sw_1_0.x1.x6.A cdac_sw_1_0.x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1125 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1126 a_125188_n9899# x4[3].x3.ckb x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1127 cdac_sw_1_2.x2.swp cdac_sw_1_2.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1128 x6[4].x3.ck x6[4].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1129 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1130 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1131 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1132 x4[2].x3.ck x4[2].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1133 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1134 x8[6].x1.x11.A x8[6].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1135 vdref x4[3].x2.swp x4[3].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1136 x3[1].x1.x10.A x3[1].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1137 vcm cdac_sw_8_0.x2.swn x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1138 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1139 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1140 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1141 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1142 vdref x10[8].x1.x7.A x10[8].x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1143 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1144 vdref cdac_sw_1_0.x2.swp cdac_sw_1_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1145 vsref cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1146 vsref cdac_sw_2_1.x2.swp cdac_sw_2_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1147 cdac_sw_1_1.x2.swp cdac_sw_1_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1148 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1149 vsref x8[7].x1.x10.A x8[7].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1150 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1151 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1152 vsref cdac_sw_4_0.x3.ckb cdac_sw_4_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1153 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1154 vsref x3[1].x1.x11.A x3[1].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1155 vcm cdac_sw_8_1.x2.swn x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1156 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1157 x2[0].x1.x10.A x2[0].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1158 vdref cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1159 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1160 vdref x4[2].x3.ckb x4[2].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1161 x4[2].x3.ck x4[2].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1162 vsref cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1163 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1164 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1165 vsref cf[6] x8[6].x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1166 vsref x3[1].x2.swp x3[1].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1167 vdref x3[1].x1.x8.A x3[1].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1168 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1169 x6[5].x2.swn x6[5].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1170 cdac_sw_8_0.x2.swp cdac_sw_8_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1171 cdac_sw_8_0.x2.swn cdac_sw_8_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1172 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1173 vsref x8[7].x3.ckb x8[7].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1174 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1175 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1176 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1177 cdac_sw_2_0.x1.x6.A cdac_sw_2_0.x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1178 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1179 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1180 vdref cdac_sw_8_1.x1.x9.A cdac_sw_8_1.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1181 vdref cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1182 vsref x6[5].x1.x11.A x6[5].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1183 x2[0].x2.swp x2[0].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1184 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1185 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1186 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1187 vsref cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1188 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1189 x6[4].x3.ck x6[4].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1190 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1191 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1192 x8[7].x3.ck x8[7].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1193 a_115667_n5199# cf[6] x8[6].x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1194 cdac_sw_2_1.x1.x4.A cf[6] a_122939_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1195 cdac_sw_4_0.x3.ckb cdac_sw_4_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1196 cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1197 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1198 x3[1].x3.ckb x3[1].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1199 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1200 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1201 cdac_sw_1_2.x3.ckb cdac_sw_1_2.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1202 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1203 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1204 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1205 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1206 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1207 vsref x4[3].x1.x11.A x4[3].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1208 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1209 x10b_cap_array_0.SW[5] cdac_sw_4_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1210 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1211 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1212 x6[5].dac_out x6[5].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1213 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1214 cdac_sw_16_0.x1.x6.A cdac_sw_16_0.x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1215 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1216 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1217 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1218 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1219 vsref cdac_sw_1_2.x3.ckb cdac_sw_1_2.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1220 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1221 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1222 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1223 cdac_sw_2_1.x2.swn cdac_sw_2_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1224 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1225 vcp x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1226 x8[7].x3.ckb x8[7].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1227 cdac_sw_1_1.x1.x6.A cdac_sw_1_1.x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1228 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1229 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1230 vsref x8[7].x1.x4.A x8[7].x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1231 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1232 vdref x3[0].x2.swp x3[0].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1233 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1234 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1235 vdref cf[4] cdac_sw_4_1.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1236 x10b_cap_array_0.SW[2] cdac_sw_8_1.x3.ckb a_109966_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1237 vsref cdac_sw_16_0.x2.swp cdac_sw_16_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1238 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1239 cdac_sw_1_2.x3.ck cdac_sw_1_2.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1240 a_110844_n15188# cdac_sw_8_1.x3.ck x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1241 cdac_sw_1_1.x3.ck cdac_sw_1_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1242 a_125327_n4335# x4[3].x1.x8.A x4[3].x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1243 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1244 x4[3].x3.ckb x4[3].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1245 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1246 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1247 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1248 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1249 vdref x6[4].x1.x11.A x6[4].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1250 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1251 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1252 cdac_sw_2_0.x2.swp cdac_sw_2_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1253 cdac_sw_2_1.x3.ckb cdac_sw_2_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1254 vdref cdac_sw_4_1.x1.x8.A cdac_sw_4_1.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1255 vdref x6[4].x2.swp x6[4].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1256 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1257 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1258 vsref cdac_sw_4_1.x3.ckb cdac_sw_4_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1259 cdac_sw_4_0.x1.x7.A cdac_sw_4_0.x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1260 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1261 a_109966_n15179# swn_in[2] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1262 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1263 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1264 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1265 vdref x8[7].x3.ckb x8[7].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1266 vdref x6[4].x1.x3.Y x6[4].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1267 vdref cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1268 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1269 vsref x8[6].x2.swp x8[6].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1270 a_118748_n7755# x6[5].x3.ckb x6[5].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1271 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1272 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1273 vsref x3[1].x1.x4.A x3[1].x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1274 x10b_cap_array_0.SW[3] cdac_sw_8_0.x3.ckb a_113186_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1275 vsref x6[5].x1.x9.A x6[5].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1276 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1277 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1278 vcm x4[3].x2.swp x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1279 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1280 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1281 x4[3].dac_out x4[3].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1282 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1283 vdref x4[3].x1.x9.A x4[3].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1284 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1285 cdac_sw_2_1.x3.ck cdac_sw_2_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1286 a_117870_n6892# swp_in[5] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1287 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1288 x10b_cap_array_0.SW[2] cdac_sw_8_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1289 cdac_sw_1_2.x3.ck cdac_sw_1_2.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1290 a_114064_n15188# cdac_sw_8_0.x3.ck x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1291 cdac_sw_4_0.x1.x4.A cf[5] a_119719_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1292 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1293 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1294 cdac_sw_4_1.x3.ckb cdac_sw_4_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1295 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1296 vdref x8[7].x1.x7.A x8[7].x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1297 x4[2].x3.ckb x4[2].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1298 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1299 x4[3].dac_out x4[3].x3.ck a_124310_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1300 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1301 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1302 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1303 x6[5].x2.swp x6[5].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1304 vsref cdac_sw_1_0.x2.swp cdac_sw_1_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1305 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1306 x10b_cap_array_0.SW[4] cdac_sw_4_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1307 cdac_sw_4_1.x1.x3.Y cf[4] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1308 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1309 x4[2].x3.ck x4[2].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1310 cdac_sw_8_1.x1.x5.A cdac_sw_8_1.x1.x8.A a_110059_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1311 vsref cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1312 x3[1].x1.x10.A x3[1].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1313 cdac_sw_8_1.x3.ckb cdac_sw_8_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1314 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1315 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1316 vdref x6[5].x1.x11.A x6[5].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1317 cdac_sw_8_0.x2.swn cdac_sw_8_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1318 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1319 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1320 vdref cf[2] x4[2].x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1321 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1322 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1323 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1324 x3[0].x2.swn x3[0].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1325 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1326 vsref x4[2].x3.ckb x4[2].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1327 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1328 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1329 x2[0].x2.swp x2[0].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1330 cdac_sw_2_0.x3.ck cdac_sw_2_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1331 vsref x3[1].x1.x8.A x3[1].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1332 vsref cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1333 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1334 vdref x6[4].x1.x9.A x6[4].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1335 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1336 cdac_sw_2_0.x1.x7.A cdac_sw_2_0.x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1337 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1338 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1339 vdref cdac_sw_2_1.x3.ckb cdac_sw_2_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1340 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1341 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1342 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1343 vsref cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1344 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1345 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1346 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1347 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1348 x6[4].x2.swn x6[4].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1349 vsref x3[0].x2.swp x3[0].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1350 vdref cdac_sw_1_2.x2.swp cdac_sw_1_2.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1351 a_124310_n8164# swp_in[3] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1352 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1353 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1354 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1355 x6[4].x3.ck x6[4].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1356 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1357 vsref cf[8] x10[8].x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1358 vdref cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1359 vdref x4[3].x1.x8.A x4[3].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1360 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1361 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1362 cdac_sw_16_0.x1.x4.A cdac_sw_16_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1363 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1364 vsref swn_in[2] a_110844_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1365 cdac_sw_16_0.x3.ck cdac_sw_16_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1366 cdac_sw_4_0.x2.swp cdac_sw_4_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1367 x3[1].x3.ckb x3[1].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1368 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1369 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1370 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1371 cdac_sw_1_2.x3.ckb cdac_sw_1_2.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1372 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1373 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1374 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1375 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1376 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1377 vcp x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1378 cdac_sw_16_0.x3.ck cdac_sw_16_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1379 vsref cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1380 vsref cdac_sw_16_0.x2.swp cdac_sw_16_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1381 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1382 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1383 x4[2].x1.x11.A x4[2].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1384 vdref x8[6].x1.x9.A x8[6].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1385 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1386 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1387 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1388 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1389 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1390 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1391 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1392 x8[7].x3.ckb x8[7].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1393 a_113186_n15179# swn_in[3] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1394 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1395 vdref x4[3].x2.swp x4[3].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1396 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1397 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1398 vsref cdac_sw_2_0.x3.ckb cdac_sw_2_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1399 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1400 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1401 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1402 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1403 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1404 vdref cdac_sw_4_1.x1.x8.A cdac_sw_4_1.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1405 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1406 x3[1].x2.swn x3[1].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1407 vdref x6[5].x1.x8.A x6[5].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1408 x4[2].dac_out x4[2].x3.ck a_127530_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1409 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1410 x2[0].x3.ckb x2[0].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1411 vsref cdac_sw_2_1.x1.x9.A cdac_sw_2_1.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1412 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1413 vdref cdac_sw_8_1.x3.ckb cdac_sw_8_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1414 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1415 x2[0].x1.x8.A x2[0].x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1416 x4[3].x3.ckb x4[3].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1417 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1418 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1419 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1420 cdac_sw_1_2.x3.ckb cdac_sw_1_2.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1421 x2[0].x3.ck x2[0].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1422 vdref cdac_sw_4_1.x1.x9.A cdac_sw_4_1.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1423 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1424 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1425 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1426 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1427 vdref cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1428 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1429 vdref cf[7] x8[7].x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1430 cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1431 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1432 vcm cdac_sw_2_1.x2.swn x10b_cap_array_0.SW[6] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1433 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1434 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1435 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1436 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1437 vdref cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1438 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1439 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1440 vsref x8[7].x3.ckb x8[7].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1441 vcm cdac_sw_8_0.x2.swn x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1442 vdref cdac_sw_1_1.x1.x8.A cdac_sw_1_1.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1443 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1444 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1445 vdref x3[1].x1.x10.A x3[1].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1446 vsref x3[0].x1.x11.A x3[0].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1447 vdref x8[6].x1.x11.A x8[6].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1448 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1449 vcn x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1450 vdref x3[1].x3.ckb x3[1].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1451 cdac_sw_4_1.x3.ck cdac_sw_4_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1452 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1453 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1454 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1455 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1456 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1457 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1458 vsref x4[3].x1.x9.A a_125327_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1459 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1460 cdac_sw_2_1.x2.swn cdac_sw_2_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1461 cdac_sw_1_2.x2.swn cdac_sw_1_2.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1462 vcp x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1463 cdac_sw_1_0.x2.swp cdac_sw_1_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1464 cdac_sw_1_2.x3.ck cdac_sw_1_2.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1465 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1466 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1467 vdref x6[5].x1.x10.A x6[5].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1468 cdac_sw_4_1.x2.swp cdac_sw_4_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1469 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1470 x3[0].x2.swp x3[0].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1471 vsref cdac_sw_8_0.x3.ckb cdac_sw_8_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1472 vdref x6[4].x1.x11.A x6[4].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1473 vsref swn_in[3] a_114064_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1474 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1475 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1476 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1477 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1478 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1479 vsref x2[0].x1.x10.A x2[0].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1480 cdac_sw_1_0.x1.x4.A cf[9] a_132599_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1481 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1482 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1483 cdac_sw_1_1.x3.ckb cdac_sw_1_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1484 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1485 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1486 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1487 x8[7].x1.x11.A x8[7].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1488 vdref x4[3].x1.x10.A x4[3].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1489 vdref swp_in[3] a_125188_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1490 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1491 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1492 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1493 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1494 vsref cdac_sw_1_2.x1.x5.A cdac_sw_1_2.x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1495 x6[5].dac_out x6[5].x3.ck a_117870_n6892# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1496 x4[2].dac_out x4[2].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1497 vsref cdac_sw_1_0.x1.x8.A cdac_sw_1_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1498 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1499 vsref cdac_sw_16_0.x1.x9.A cdac_sw_16_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1500 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1501 x6[4].x2.swn x6[4].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1502 x10b_cap_array_0.SW[2] cdac_sw_8_1.x3.ckb a_109966_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1503 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1504 cdac_sw_1_0.x2.swn cdac_sw_1_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1505 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1506 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1507 x6[4].x1.x5.A x6[4].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1508 vdref x2[0].x3.ckb x2[0].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1509 vsref cdac_sw_1_1.x2.swp cdac_sw_1_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1510 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1511 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1512 x4[2].x2.swp x4[2].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1513 cdac_sw_16_0.x3.ck cdac_sw_16_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1514 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1515 a_109966_n15179# swn_in[2] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1516 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1517 cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1518 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1519 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1520 vdref cf[7] cdac_sw_2_0.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1521 vdref cdac_sw_2_1.x2.swp cdac_sw_2_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1522 vsref cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1523 cdac_sw_4_0.x2.swp cdac_sw_4_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1524 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1525 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1526 a_120504_n15188# cdac_sw_4_0.x3.ck x10b_cap_array_0.SW[5] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1527 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1528 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1529 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1530 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1531 x4[3].x1.x4.A cf[3] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1532 cdac_sw_8_1.x2.swn cdac_sw_8_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1533 x10b_cap_array_0.SW[9] cdac_sw_1_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1534 x4[2].x2.swn x4[2].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1535 vdref swp_in[2] a_128408_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1536 vdref cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1537 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1538 x3[1].x1.x11.A x3[1].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1539 cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1540 vsref x4[3].x1.x8.A x4[3].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1541 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1542 vsref x4[3].x1.x7.A x4[3].x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1543 cdac_sw_1_0.x3.ckb cdac_sw_1_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1544 cdac_sw_16_0.x1.x5.A cdac_sw_16_0.x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1545 vdref cdac_sw_2_0.x1.x8.A cdac_sw_2_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1546 cdac_sw_16_0.x2.swp cdac_sw_16_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1547 cdac_sw_16_0.x2.swn cdac_sw_16_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1548 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1549 cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1550 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1551 vdref cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1552 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1553 vsref x4[2].x2.swp x4[2].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1554 vdref x8[6].x3.ckb x8[6].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1555 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1556 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1557 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1558 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1559 x3[0].x2.swn x3[0].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1560 x4[3].x2.swp x4[3].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1561 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1562 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1563 vcp x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1564 vdref x6[5].x1.x8.A x6[5].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1565 vdref swp_in[2] a_128408_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1566 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1567 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1568 x2[0].x3.ck x2[0].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1569 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1570 a_127530_n8164# swp_in[2] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1571 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1572 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1573 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1574 x8[6].dac_out x8[6].x3.ck a_114650_n6256# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1575 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1576 vsref cdac_sw_16_0.x1.x8.A cdac_sw_16_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1577 cdac_sw_1_1.x1.x4.A cf[8] a_129379_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1578 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1579 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1580 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1581 cdac_sw_8_0.x1.x9.A cdac_sw_8_0.x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1582 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1583 vsref x6[5].x1.x8.A x6[5].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1584 vdref cdac_sw_16_0.x3.ckb cdac_sw_16_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1585 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1586 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1587 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1588 vdref cdac_sw_8_1.x2.swp cdac_sw_8_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1589 x2[0].x1.x9.A x2[0].x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1590 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1591 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1592 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1593 cdac_sw_1_2.x2.swp cdac_sw_1_2.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1594 x10b_cap_array_0.SW[3] cdac_sw_8_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1595 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1596 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1597 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1598 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1599 vsref cdac_sw_8_1.x2.swp cdac_sw_8_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1600 cdac_sw_1_2.x3.ckb cdac_sw_1_2.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1601 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1602 cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1603 vdref cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1604 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1605 vsref x6[4].x2.swp x6[4].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1606 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1607 cdac_sw_1_2.x2.swn cdac_sw_1_2.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1608 cdac_sw_4_0.x3.ckb cdac_sw_4_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1609 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1610 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1611 vsref cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1612 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1613 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1614 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1615 cdac_sw_4_0.x1.x8.A cdac_sw_4_0.x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1616 vcm cdac_sw_8_1.x2.swn x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1617 vdref cdac_sw_2_1.x1.x8.A cdac_sw_2_1.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1618 cdac_sw_2_1.x2.swn cdac_sw_2_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1619 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1620 cdac_sw_4_0.x3.ck cdac_sw_4_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1621 vdref cdac_sw_1_1.x1.x9.A cdac_sw_1_1.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1622 x8[7].x2.swp x8[7].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1623 vsref x3[1].x1.x10.A x3[1].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1624 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1625 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1626 x3[0].x3.ck x3[0].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1627 vcp x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1628 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1629 x6[5].x2.swn x6[5].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1630 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1631 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1632 vsref x3[1].x3.ckb x3[1].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1633 cdac_sw_4_1.x2.swn cdac_sw_4_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1634 a_106839_n16821# x2[0].x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1635 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1636 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1637 cdac_sw_8_0.x3.ckb cdac_sw_8_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1638 vsref cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1639 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1640 cdac_sw_8_1.x1.x3.Y cf[2] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1641 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1642 vdref cf[9] cdac_sw_1_2.x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1643 cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1644 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1645 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1646 vsref x4[2].x1.x9.A x4[2].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1647 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1648 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1649 x8[7].x2.swn x8[7].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1650 vdref swp_in[7] a_112308_n6683# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1651 vdref cdac_sw_1_0.x3.ckb cdac_sw_1_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1652 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1653 x6[4].x3.ck x6[4].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1654 vsref x6[5].x1.x10.A x6[5].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1655 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1656 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1657 vdref x3[0].x3.ckb x3[0].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1658 cdac_sw_1_1.x3.ck cdac_sw_1_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1659 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1660 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1661 vcm x4[3].x2.swp x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1662 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1663 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1664 x4[3].x2.swn x4[3].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1665 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1666 vdref cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1667 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1668 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1669 x4[3].x1.x11.A x4[3].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1670 cdac_sw_8_0.x1.x4.A cdac_sw_8_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1671 cdac_sw_2_1.x3.ckb cdac_sw_2_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1672 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1673 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1674 vsref x8[7].x2.swp x8[7].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1675 vdref cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1676 vdref x6[5].x1.x5.A x6[5].x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1677 cdac_sw_1_1.x2.swp cdac_sw_1_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1678 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1679 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1680 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1681 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1682 cdac_sw_2_1.x1.x8.A cdac_sw_2_1.x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1683 vsref x4[3].x1.x10.A x4[3].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1684 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1685 x4[2].x2.swp x4[2].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1686 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1687 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1688 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1689 vsref cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1690 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1691 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1692 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1693 x4[2].x1.x10.A x4[2].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1694 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1695 a_126944_n15188# cdac_sw_2_0.x3.ck x10b_cap_array_0.SW[7] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1696 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1697 x10b_cap_array_0.SW[5] cdac_sw_4_0.x3.ckb a_119626_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1698 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1699 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1700 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1701 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1702 vdref x2[0].x2.swp x2[0].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1703 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1704 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1705 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1706 cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1707 vdref swp_in[5] a_118748_n7755# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1708 vcm x4[2].x2.swp x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1709 vsref swn_in[3] a_114064_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1710 cdac_sw_16_0.x2.swn cdac_sw_16_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1711 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1712 vsref x4[2].x1.x11.A x4[2].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1713 a_121090_n6892# swp_in[4] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1714 a_110844_n15188# cdac_sw_8_1.x3.ck x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1715 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1716 x3[0].x2.swp x3[0].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1717 vsref x2[0].x2.swp x2[0].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1718 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1719 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1720 vdref cdac_sw_2_0.x1.x8.A cdac_sw_2_0.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1721 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1722 x3[1].x3.ck x3[1].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1723 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1724 vdref cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1725 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1726 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1727 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1728 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1729 x6[5].x1.x11.A x6[5].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1730 vcn x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1731 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1732 vsref cdac_sw_1_2.x2.swp cdac_sw_1_2.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1733 a_125327_n5199# cf[3] x4[3].x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1734 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1735 cdac_sw_4_1.x1.x8.A cdac_sw_4_1.x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1736 a_122846_n15179# swn_in[6] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1737 a_116499_n15957# cdac_sw_4_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1738 cdac_sw_2_0.x3.ckb cdac_sw_2_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1739 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1740 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1741 vdref x3[1].x1.x11.A x3[1].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1742 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1743 vdref cdac_sw_2_0.x1.x9.A cdac_sw_2_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1744 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1745 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1746 vsref x3[0].x1.x11.A x3[0].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1747 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1748 vcm x4[2].x2.swp x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1749 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1750 cdac_sw_8_1.x3.ckb cdac_sw_8_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1751 cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1752 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1753 vcm cdac_sw_1_0.x2.swn x10b_cap_array_0.SW[9] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1754 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1755 vsref x6[5].x1.x3.Y a_118887_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1756 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1757 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1758 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1759 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1760 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1761 vdref cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1762 vsref x8[6].x3.ckb x8[6].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1763 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1764 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1765 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1766 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1767 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1768 vdref x3[0].x1.x10.A x3[0].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1769 a_125188_n9899# x4[3].x3.ckb x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1770 vsref x8[7].x1.x9.A x8[7].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1771 x3[1].x2.swp x3[1].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1772 vsref x6[5].x1.x8.A x6[5].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1773 vsref x6[5].x1.x7.A x6[5].x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1774 cdac_sw_2_0.x3.ck cdac_sw_2_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1775 vdref cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1776 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1777 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1778 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1779 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1780 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1781 cdac_sw_1_2.x3.ck cdac_sw_1_2.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1782 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1783 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1784 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1785 x3[0].x3.ckb x3[0].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1786 x6[5].x2.swp x6[5].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1787 vsref cdac_sw_2_1.x3.ckb cdac_sw_2_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1788 vdref cdac_sw_16_0.x2.swp cdac_sw_16_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1789 vsref swn_in[6] a_123724_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1790 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1791 cdac_sw_4_0.x3.ck cdac_sw_4_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1792 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1793 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1794 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1795 vsref cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1796 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1797 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1798 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1799 a_116406_n15179# swn_in[4] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1800 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1801 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1802 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1803 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1804 cdac_sw_8_0.x3.ckb cdac_sw_8_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1805 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1806 x8[7].x1.x10.A x8[7].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1807 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1808 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1809 cdac_sw_4_1.x2.swn cdac_sw_4_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1810 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1811 vsref x3[1].x1.x9.A x3[1].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1812 vdref cdac_sw_1_2.x1.x4.A cdac_sw_1_2.x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1813 x4[3].x2.swp x4[3].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1814 cdac_sw_4_0.x1.x9.A cdac_sw_4_0.x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1815 vdref cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1816 vdref cdac_sw_2_1.x1.x9.A cdac_sw_2_1.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1817 vsref cdac_sw_8_0.x1.x9.A cdac_sw_8_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1818 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1819 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1820 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1821 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1822 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1823 cdac_sw_1_1.x1.x8.A cdac_sw_1_1.x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1824 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1825 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1826 vcm x8[7].x2.swp x8[7].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1827 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1828 vsref x8[7].x1.x11.A x8[7].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1829 x3[0].x3.ck x3[0].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1830 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1831 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1832 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1833 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1834 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1835 x4[2].x3.ckb x4[2].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1836 vdref x4[3].x1.x11.A x4[3].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1837 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1838 cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1839 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1840 vdref x6[4].x1.x7.A x6[4].x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1841 a_119626_n15179# swn_in[5] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1842 x10b_cap_array_0.SW[5] cdac_sw_4_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1843 vdref cdac_sw_2_0.x3.ckb cdac_sw_2_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1844 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1845 vdref cdac_sw_1_0.x2.swp cdac_sw_1_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1846 cdac_sw_1_2.x2.swp cdac_sw_1_2.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1847 x6[4].x3.ck x6[4].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1848 vsref x3[0].x3.ckb x3[0].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1849 cdac_sw_1_1.x2.swn cdac_sw_1_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1850 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1851 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1852 x4[2].x3.ck x4[2].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1853 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1854 x3[1].x1.x10.A x3[1].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1855 cdac_sw_2_1.x1.x3.Y cf[6] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1856 cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1857 vdref x4[3].x2.swp x4[3].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1858 vdref cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1859 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1860 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1861 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1862 vdref x4[3].x1.x6.A x4[3].x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1863 vcm cdac_sw_8_1.x2.swn x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1864 cdac_sw_8_0.x1.x5.A cdac_sw_8_0.x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1865 cdac_sw_2_1.x2.swp cdac_sw_2_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1866 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1867 vdref cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1868 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1869 cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1870 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1871 vsref x3[1].x1.x11.A x3[1].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1872 x10b_cap_array_0.SW[2] cdac_sw_8_1.x3.ckb a_109966_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1873 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1874 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1875 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1876 vsref cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1877 vsref cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1878 vdref x4[2].x3.ckb x4[2].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1879 vsref x3[1].x2.swp x3[1].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1880 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1881 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1882 x3[0].x3.ck x3[0].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1883 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1884 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1885 x4[2].x1.x10.A x4[2].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1886 x4[2].dac_out x4[2].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1887 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1888 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1889 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1890 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1891 a_109966_n15179# swn_in[2] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1892 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1893 x6[5].x1.x11.A x6[5].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1894 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1895 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1896 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1897 cdac_sw_4_1.x3.ck cdac_sw_4_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1898 a_118748_n7755# x6[5].x3.ckb x6[5].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1899 cdac_sw_1_0.x1.x7.A cdac_sw_1_0.x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1900 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1901 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1902 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1903 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1904 x3[1].x2.swn x3[1].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1905 vdref x6[5].x2.swp x6[5].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1906 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1907 x3[1].x3.ck x3[1].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1908 vdref cdac_sw_8_0.x3.ckb cdac_sw_8_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1909 vdref cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1910 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1911 vsref cf[5] x6[5].x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1912 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1913 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1914 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1915 cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1916 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1917 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1918 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1919 cdac_sw_4_1.x1.x9.A cdac_sw_4_1.x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1920 cdac_sw_1_2.x3.ckb cdac_sw_1_2.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1921 vsref cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1922 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1923 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1924 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1925 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1926 vdref x2[0].x1.x10.A x2[0].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1927 vsref cdac_sw_4_0.x2.swp cdac_sw_4_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1928 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1929 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1930 vdref x6[4].x3.ckb x6[4].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1931 x2[0].x1.x11.A x2[0].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1932 cdac_sw_8_1.x2.swp cdac_sw_8_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1933 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1934 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1935 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1936 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1937 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1938 vdref cdac_sw_1_0.x1.x8.A cdac_sw_1_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1939 vdref x4[3].x1.x9.A x4[3].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1940 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1941 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1942 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1943 x8[7].x3.ckb x8[7].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1944 x10b_cap_array_0.SW[4] cdac_sw_4_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1945 vsref x3[0].x1.x10.A x3[0].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1946 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1947 vdref x3[0].x2.swp x3[0].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1948 cdac_sw_2_0.x2.swn cdac_sw_2_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1949 vdref cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1950 vcp x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1951 vsref cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1952 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1953 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1954 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1955 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1956 cdac_sw_1_2.x3.ck cdac_sw_1_2.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1957 cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1958 cdac_sw_4_0.x1.x3.Y cf[5] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1959 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1960 x8[7].x3.ck x8[7].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1961 vdref x4[2].x1.x8.A x4[2].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1962 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1963 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1964 a_127530_n8164# swp_in[2] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1965 cdac_sw_2_1.x1.x5.A cdac_sw_2_1.x1.x8.A a_122939_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1966 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1967 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1968 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1969 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1970 vsref cdac_sw_4_1.x3.ckb cdac_sw_4_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1971 vsref swn_in[5] a_120504_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1972 x3[0].x3.ckb x3[0].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1973 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1974 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1975 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1976 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1977 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1978 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1979 vsref cdac_sw_1_2.x1.x9.A cdac_sw_1_2.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1980 cdac_sw_8_0.x3.ck cdac_sw_8_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1981 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1982 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1983 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1984 cdac_sw_16_0.x1.x7.A cdac_sw_16_0.x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1985 vdref x8[7].x3.ckb x8[7].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1986 vsref x8[6].x2.swp x8[6].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1987 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1988 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1989 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1990 x8[7].x1.x10.A x8[7].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1991 cdac_sw_1_0.x1.x8.A cdac_sw_1_0.x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1992 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1993 x4[2].x3.ckb x4[2].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1994 vsref cdac_sw_1_2.x1.x4.A cdac_sw_1_2.x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1995 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1996 vdref x4[3].x1.x11.A x4[3].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1997 vdref x4[2].x2.swp x4[2].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1998 vdref cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1999 cdac_sw_1_1.x1.x7.A cdac_sw_1_1.x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2000 cdac_sw_1_1.x1.x9.A cdac_sw_1_1.x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2001 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2002 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2003 a_125188_n9899# x4[3].x3.ckb x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2004 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2005 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2006 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2007 cdac_sw_4_1.x3.ckb cdac_sw_4_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2008 x8[6].x2.swn x8[6].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2009 a_118887_n4335# x6[5].x1.x8.A x6[5].x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2010 vsref cdac_sw_1_1.x3.ckb cdac_sw_1_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2011 cdac_sw_1_1.x2.swn cdac_sw_1_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2012 cdac_sw_8_1.x1.x6.A cdac_sw_8_1.x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2013 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2014 cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2015 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2016 cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2017 vdref x4[2].x1.x10.A x4[2].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2018 x4[2].x3.ckb x4[2].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2019 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2020 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2021 a_120504_n15188# cdac_sw_4_0.x3.ck x10b_cap_array_0.SW[5] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2022 x3[0].x3.ckb x3[0].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2023 vdref cdac_sw_2_0.x2.swp cdac_sw_2_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2024 vsref cdac_sw_4_1.x2.swp cdac_sw_4_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2025 cdac_sw_2_1.x2.swp cdac_sw_2_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2026 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2027 x6[5].x2.swp x6[5].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2028 vdref x3[1].x1.x11.A x3[1].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2029 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2030 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2031 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2032 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2033 vdref x8[6].x1.x3.Y x8[6].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2034 vdref cdac_sw_1_2.x3.ckb cdac_sw_1_2.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2035 vsref x10[8].x2.swp x10[8].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2036 x4[2].x3.ck x4[2].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2037 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2038 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2039 x3[1].x1.x10.A x3[1].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2040 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2041 a_132506_n15179# swn_in[9] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2042 a_126159_n15957# cdac_sw_2_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2043 cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2044 vdref x3[0].x1.x10.A x3[0].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2045 vsref x4[3].x1.x6.A x4[3].x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2046 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2047 vdref x6[5].x1.x11.A x6[5].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2048 vdref x8[6].x1.x7.A x8[6].x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2049 cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2050 vdref x6[5].x1.x9.A x6[5].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2051 a_114064_n15188# cdac_sw_8_0.x3.ck x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2052 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2053 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2054 x3[0].x2.swn x3[0].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2055 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2056 x10[8].x2.swn x10[8].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2057 vsref x4[2].x3.ckb x4[2].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2058 x3[0].x3.ck x3[0].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2059 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2060 cdac_sw_4_0.x1.x5.A cdac_sw_4_0.x1.x8.A a_119719_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2061 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2062 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2063 vsref cf[4] x6[4].x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2064 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2065 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2066 vdref x8[7].x1.x8.A x8[7].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2067 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2068 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2069 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2070 vdref x6[5].x1.x6.A x6[5].x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2071 a_110844_n15188# cdac_sw_8_1.x3.ck x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2072 vsref swn_in[4] a_117284_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2073 cdac_sw_8_0.x1.x6.A cdac_sw_8_0.x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2074 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2075 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2076 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2077 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2078 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2079 x8[6].x2.swn x8[6].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2080 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2081 vdref cdac_sw_8_0.x2.swp cdac_sw_8_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2082 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2083 cdac_sw_8_1.x2.swp cdac_sw_8_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2084 vsref x3[0].x1.x5.A x3[0].x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2085 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2086 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2087 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2088 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2089 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2090 cdac_sw_1_2.x3.ckb cdac_sw_1_2.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2091 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2092 vdref x2[0].x1.x11.A x2[0].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2093 vsref x6[4].x3.ckb x6[4].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2094 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2095 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2096 x10b_cap_array_0.SW[2] cdac_sw_8_1.x3.ckb a_109966_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2097 x4[3].dac_out x4[3].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2098 cdac_sw_2_0.x2.swn cdac_sw_2_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2099 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2100 vdref x3[1].x1.x8.A x3[1].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2101 x2[0].x1.x6.A x2[0].x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2102 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2103 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2104 vdref cdac_sw_1_0.x1.x9.A cdac_sw_1_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2105 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2106 vdref cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2107 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2108 vcn x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2109 vdref x8[7].x1.x10.A x8[7].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2110 x8[7].x3.ckb x8[7].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2111 x4[2].dac_out x4[2].x3.ck a_127530_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2112 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2113 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2114 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2115 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2116 a_109966_n15179# swn_in[2] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2117 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2118 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2119 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2120 x4[3].dac_out x4[3].x3.ck a_124310_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2121 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2122 cdac_sw_16_0.x1.x4.A cf[0] a_103619_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2123 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2124 x3[1].x2.swn x3[1].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2125 vdref swp_in[3] a_125188_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2126 vsref swn_in[2] a_110844_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2127 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2128 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2129 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2130 x3[0].x1.x11.A x3[0].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2131 cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2132 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2133 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2134 vdref x4[2].x1.x11.A x4[2].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2135 vsref x4[2].x1.x8.A x4[2].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2136 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2137 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2138 x8[7].x3.ck x8[7].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2139 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2140 vcp x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2141 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2142 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2143 cdac_sw_1_2.x3.ckb cdac_sw_1_2.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2144 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2145 cdac_sw_1_0.x1.x3.Y cf[9] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2146 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2147 vdref x4[2].x2.swp x4[2].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2148 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2149 cdac_sw_8_0.x2.swn cdac_sw_8_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2150 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2151 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2152 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2153 cdac_sw_16_0.x2.swn cdac_sw_16_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2154 vsref cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2155 vsref cdac_sw_1_1.x3.ckb cdac_sw_1_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2156 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2157 vsref x8[7].x3.ckb x8[7].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2158 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2159 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2160 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2161 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2162 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2163 vdref x3[1].x1.x10.A x3[1].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2164 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2165 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2166 vdref cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2167 vsref cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2168 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2169 vsref x10[8].x1.x11.A x10[8].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2170 x4[2].x3.ckb x4[2].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2171 vdref x3[1].x3.ckb x3[1].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2172 x4[2].x2.swn x4[2].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2173 vdref swp_in[2] a_128408_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2174 vsref cdac_sw_2_0.x2.swp cdac_sw_2_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2175 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2176 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2177 cdac_sw_8_1.x3.ck cdac_sw_8_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2178 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2179 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2180 cdac_sw_4_1.x2.swp cdac_sw_4_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2181 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2182 a_124310_n8164# swp_in[3] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2183 x2[0].x2.swp x2[0].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2184 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2185 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2186 vcn x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2187 cdac_sw_8_1.x1.x7.A cdac_sw_8_1.x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2188 x3[0].x2.swp x3[0].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2189 cdac_sw_16_0.x3.ckb cdac_sw_16_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2190 a_117284_n15188# cdac_sw_4_1.x3.ck x10b_cap_array_0.SW[4] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2191 cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2192 vsref x4[2].x1.x10.A x4[2].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2193 x3[1].x3.ck x3[1].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2194 x3[0].x3.ckb x3[0].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2195 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2196 x2[0].x2.swn x2[0].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2197 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2198 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2199 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2200 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2201 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2202 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2203 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2204 vdref x6[4].x2.swp x6[4].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2205 x3[0].x2.swn x3[0].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2206 vdref cdac_sw_2_1.x3.ckb cdac_sw_2_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2207 cdac_sw_1_1.x3.ckb cdac_sw_1_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2208 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2209 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2210 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2211 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2212 vcm cdac_sw_8_0.x2.swn x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2213 cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2214 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2215 vsref cdac_sw_1_2.x3.ckb cdac_sw_1_2.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2216 x10[8].x2.swn x10[8].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2217 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2218 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2219 vdref x4[2].x1.x5.A x4[2].x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2220 vdref cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2221 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2222 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2223 x10b_cap_array_0.SW[4] cdac_sw_4_1.x3.ckb a_116406_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2224 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2225 cdac_sw_8_0.x3.ckb cdac_sw_8_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2226 vsref x3[0].x1.x10.A x3[0].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2227 x6[4].x2.swn x6[4].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2228 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2229 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2230 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2231 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2232 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2233 vsref x6[5].x1.x9.A a_118887_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2234 cdac_sw_1_1.x3.ck cdac_sw_1_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2235 x10b_cap_array_0.SW[3] cdac_sw_8_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2236 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2237 x8[6].x2.swn x8[6].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2238 vdref x8[7].x1.x11.A x8[7].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2239 vsref x8[7].x1.x8.A x8[7].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2240 vsref x6[5].x1.x6.A x6[5].x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2241 vsref cdac_sw_8_0.x2.swp cdac_sw_8_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2242 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2243 vsref cdac_sw_8_1.x3.ckb cdac_sw_8_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2244 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2245 x4[2].x2.swn x4[2].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2246 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2247 cdac_sw_1_1.x1.x3.Y cf[8] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2248 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2249 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2250 vsref x2[0].x1.x11.A x2[0].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2251 cdac_sw_1_0.x1.x5.A cdac_sw_1_0.x1.x8.A a_132599_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2252 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2253 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2254 vdref x8[7].x2.swp x8[7].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2255 vsref cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2256 vsref cdac_sw_2_0.x3.ckb cdac_sw_2_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2257 cdac_sw_1_0.x3.ckb cdac_sw_1_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2258 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2259 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2260 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2261 vcm cdac_sw_2_1.x2.swn x10b_cap_array_0.SW[6] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2262 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2263 vdref cdac_sw_1_2.x1.x8.A cdac_sw_1_2.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2264 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2265 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2266 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2267 cdac_sw_2_1.x3.ck cdac_sw_2_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2268 vsref cdac_sw_1_0.x1.x9.A cdac_sw_1_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2269 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2270 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2271 vdref x8[6].x3.ckb x8[6].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2272 x2[0].x3.ck x2[0].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2273 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2274 x8[7].x2.swn x8[7].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2275 x8[6].x1.x5.A x8[6].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2276 vdref swp_in[7] a_112308_n6683# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2277 x10[8].x2.swn x10[8].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2278 vsref x3[1].x1.x8.A x3[1].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2279 vcm x4[3].x2.swp x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2280 x2[0].x1.x7.A x2[0].x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2281 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2282 x3[0].x1.x11.A x3[0].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2283 x10b_cap_array_0.SW[5] cdac_sw_4_0.x3.ckb a_119626_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2284 vdref cdac_sw_16_0.x3.ckb cdac_sw_16_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2285 vdref cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2286 cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2287 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2288 x10[8].x1.x11.A x10[8].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2289 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2290 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2291 vsref x8[7].x1.x10.A x8[7].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2292 vcp x3[1].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2293 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2294 x8[6].x3.ck x8[6].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2295 x6[5].x1.x4.A cf[5] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2296 cdac_sw_2_0.x3.ckb cdac_sw_2_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2297 vsref x3[0].x2.swp x3[0].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2298 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2299 vdref cdac_sw_1_2.x2.swp cdac_sw_1_2.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2300 cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2301 cdac_sw_4_0.x1.x6.A cdac_sw_4_0.x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2302 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2303 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2304 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2305 cdac_sw_1_0.x2.swp cdac_sw_1_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2306 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2307 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2308 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2309 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2310 vdref x8[7].x1.x5.A x8[7].x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2311 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2312 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2313 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2314 cdac_sw_1_2.x3.ckb cdac_sw_1_2.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2315 vdref x10[8].x3.ckb x10[8].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2316 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2317 cdac_sw_2_0.x3.ck cdac_sw_2_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2318 cdac_sw_1_2.x2.swn cdac_sw_1_2.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2319 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2320 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2321 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2322 x6[5].dac_out x6[5].x3.ck a_117870_n6892# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2323 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2324 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2325 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2326 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2327 vdref swp_in[5] a_118748_n7755# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2328 vcm x4[2].x2.swp x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2329 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2330 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2331 x4[2].x1.x11.A x4[2].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2332 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2333 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2334 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2335 cdac_sw_16_0.x3.ckb cdac_sw_16_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2336 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2337 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2338 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2339 x8[7].x2.swp x8[7].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2340 vsref x3[1].x1.x10.A x3[1].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2341 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2342 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2343 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2344 x3[0].x3.ck x3[0].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2345 vsref cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2346 vsref x2[0].x3.ckb x2[0].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2347 x2[0].x2.swn x2[0].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2348 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2349 x10[8].x3.ck x10[8].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2350 vcm x6[4].x2.swp x6[4].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2351 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2352 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2353 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2354 vsref x3[1].x3.ckb x3[1].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2355 vsref cdac_sw_16_0.x1.x9.A cdac_sw_16_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2356 cdac_sw_1_1.x1.x5.A cdac_sw_1_1.x1.x8.A a_129379_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2357 a_114064_n15188# cdac_sw_8_0.x3.ck x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2358 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2359 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2360 vdref cdac_sw_1_0.x3.ckb cdac_sw_1_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2361 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2362 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2363 vsref x4[2].x1.x9.A x4[2].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2364 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2365 cdac_sw_2_1.x1.x6.A cdac_sw_2_1.x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2366 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2367 vdref x3[1].x1.x5.A x3[1].x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2368 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2369 vdref swp_in[3] a_125188_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2370 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2371 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2372 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2373 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2374 vdref cf[2] cdac_sw_8_1.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2375 vdref cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2376 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2377 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2378 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2379 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2380 x8[6].x3.ck x8[6].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2381 x3[1].x3.ck x3[1].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2382 a_125188_n9899# x4[3].x3.ckb x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2383 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2384 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2385 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2386 cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2387 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2388 cdac_sw_8_0.x3.ck cdac_sw_8_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2389 vdref cdac_sw_2_1.x2.swp cdac_sw_2_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2390 cdac_sw_1_1.x2.swp cdac_sw_1_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2391 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2392 cdac_sw_4_0.x2.swp cdac_sw_4_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2393 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2394 vdref x3[0].x1.x4.A x3[0].x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2395 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2396 vsref cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2397 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2398 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2399 x4[2].x2.swp x4[2].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2400 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2401 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2402 x2[0].x3.ckb x2[0].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2403 vdref cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2404 cdac_sw_4_0.x2.swn cdac_sw_4_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2405 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2406 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2407 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2408 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2409 x4[2].x2.swp x4[2].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2410 vdref cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2411 cdac_sw_8_0.x2.swp cdac_sw_8_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2412 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2413 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2414 x4[2].x2.swn x4[2].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2415 cdac_sw_8_0.x2.swp cdac_sw_8_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2416 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2417 x3[1].x1.x11.A x3[1].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2418 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2419 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2420 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2421 vdref swp_in[2] a_128408_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2422 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2423 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2424 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2425 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2426 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2427 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2428 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2429 a_116406_n15179# swn_in[4] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2430 a_119626_n15179# swn_in[5] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2431 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2432 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2433 x3[0].x2.swp x3[0].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2434 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2435 x10[8].x2.swp x10[8].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2436 cdac_sw_8_0.x1.x4.A cf[3] a_113279_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2437 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2438 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2439 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2440 x3[1].x3.ck x3[1].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2441 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2442 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2443 vsref x3[1].x1.x3.Y a_131767_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2444 vdref x4[2].x2.swp x4[2].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2445 x3[0].x1.x10.A x3[0].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2446 vsref swn_in[5] a_120504_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2447 vdref x3[1].x1.x9.A x3[1].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2448 vsref cdac_sw_1_2.x2.swp cdac_sw_1_2.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2449 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2450 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2451 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2452 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2453 vsref swn_in[2] a_110844_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2454 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2455 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2456 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2457 vcm x8[7].x2.swp x8[7].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2458 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2459 x8[7].x1.x11.A x8[7].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2460 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2461 vsref cdac_sw_8_0.x1.x8.A cdac_sw_8_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2462 vdref cdac_sw_16_0.x3.ckb cdac_sw_16_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2463 cdac_sw_2_1.x1.x9.A cdac_sw_2_1.x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2464 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2465 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2466 vsref x3[0].x1.x11.A x3[0].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2467 vdref cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2468 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2469 vsref x3[1].x1.x7.A x3[1].x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2470 vsref cdac_sw_1_2.x1.x8.A cdac_sw_1_2.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2471 x10b_cap_array_0.SW[9] cdac_sw_1_0.x3.ckb a_132506_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2472 cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2473 cdac_sw_2_1.x2.swn cdac_sw_2_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2474 vsref cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2475 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2476 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2477 x6[4].x2.swn x6[4].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2478 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2479 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2480 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2481 vsref x8[6].x3.ckb x8[6].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2482 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2483 x10b_cap_array_0.SW[8] cdac_sw_1_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2484 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2485 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2486 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2487 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2488 vsref x8[7].x1.x9.A x8[7].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2489 vdref x10[8].x1.x10.A x10[8].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2490 x3[1].x2.swp x3[1].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2491 vsref cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2492 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2493 cdac_sw_1_2.x2.swp cdac_sw_1_2.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2494 vdref cdac_sw_16_0.x2.swp cdac_sw_16_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2495 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2496 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2497 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2498 vdref cdac_sw_2_1.x1.x8.A cdac_sw_2_1.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2499 cdac_sw_4_0.x3.ck cdac_sw_4_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2500 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2501 x8[6].x3.ck x8[6].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2502 a_118887_n5199# cf[5] x6[5].x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2503 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2504 x4[2].dac_out x4[2].x3.ck a_127530_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2505 cdac_sw_2_0.x2.swp cdac_sw_2_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2506 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2507 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2508 x3[0].x3.ckb x3[0].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2509 vdref swp_in[9] a_105868_n6147# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2510 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2511 cdac_sw_4_0.x1.x7.A cdac_sw_4_0.x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2512 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2513 cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2514 a_116499_n16821# cdac_sw_4_1.x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2515 cdac_sw_2_0.x2.swp cdac_sw_2_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2516 vsref x4[2].x1.x11.A x4[2].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2517 x8[7].x2.swp x8[7].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2518 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2519 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2520 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2521 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2522 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2523 x8[7].x2.swp x8[7].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2524 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2525 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2526 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2527 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2528 x10[8].x3.ck x10[8].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2529 vsref x10[8].x3.ckb x10[8].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2530 x4[3].dac_out x4[3].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2531 a_118748_n7755# x6[5].x3.ckb x6[5].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2532 x10b_cap_array_0.SW[7] cdac_sw_2_0.x3.ckb a_126066_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2533 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2534 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2535 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2536 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2537 x4[3].x2.swp x4[3].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2538 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2539 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2540 cdac_sw_1_0.x3.ckb cdac_sw_1_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2541 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2542 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2543 vcm x4[3].x2.swp x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2544 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2545 x3[0].x3.ck x3[0].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2546 x4[3].dac_out x4[3].x3.ck a_124310_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2547 x10b_cap_array_0.SW[6] cdac_sw_2_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2548 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2549 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2550 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2551 x10[8].x3.ck x10[8].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2552 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2553 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2554 a_110844_n15188# cdac_sw_8_1.x3.ck x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2555 vsref swn_in[4] a_117284_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2556 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2557 x8[6].x3.ck x8[6].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2558 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2559 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2560 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2561 vdref x8[7].x2.swp x8[7].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2562 vdref cdac_sw_1_0.x2.swp cdac_sw_1_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2563 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2564 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2565 vsref cdac_sw_2_1.x2.swp cdac_sw_2_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2566 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2567 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2568 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2569 vsref x3[0].x1.x9.A x3[0].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2570 vsref cdac_sw_4_0.x3.ckb cdac_sw_4_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2571 cdac_sw_4_0.x2.swn cdac_sw_4_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2572 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2573 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2574 x2[0].x1.x10.A x2[0].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2575 vdref cdac_sw_8_1.x1.x8.A cdac_sw_8_1.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2576 x10b_cap_array_0.SW[8] cdac_sw_1_1.x3.ckb a_129286_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2577 vdref cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2578 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2579 vsref cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2580 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2581 vdref x4[3].x1.x3.Y x4[3].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2582 x8[6].x3.ck x8[6].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2583 vcm x8[6].x2.swp x8[6].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2584 vsref cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2585 cdac_sw_8_0.x2.swp cdac_sw_8_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2586 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2587 vsref x6[5].x2.swp x6[5].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2588 cdac_sw_8_0.x2.swn cdac_sw_8_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2589 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2590 cdac_sw_1_2.x2.swn cdac_sw_1_2.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2591 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2592 cdac_sw_8_1.x3.ckb cdac_sw_8_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2593 vdref cdac_sw_16_0.x1.x8.A cdac_sw_16_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2594 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2595 x10b_cap_array_0.SW[7] cdac_sw_2_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2596 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2597 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2598 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2599 vsref x3[0].x1.x4.A x3[0].x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2600 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2601 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2602 cdac_sw_1_0.x3.ck cdac_sw_1_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2603 vcm x4[2].x2.swp x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2604 x2[0].x2.swp x2[0].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2605 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2606 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2607 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2608 vsref cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2609 x4[2].dac_out x4[2].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2610 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2611 vdref cdac_sw_1_1.x3.ckb cdac_sw_1_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2612 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2613 vdref cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2614 x10[8].x3.ck x10[8].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2615 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2616 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2617 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2618 a_124310_n8164# swp_in[3] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2619 vdref cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2620 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2621 vsref cf[1] x3[1].x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2622 x3[0].x1.x10.A x3[0].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2623 cdac_sw_4_0.x3.ckb cdac_sw_4_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2624 vsref cdac_sw_1_2.x1.x3.Y a_106007_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2625 x10[8].x1.x10.A x10[8].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2626 cdac_sw_8_1.x3.ck cdac_sw_8_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2627 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2628 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2629 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2630 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2631 vsref x8[7].x1.x11.A x8[7].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2632 vdref x3[0].x3.ckb x3[0].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2633 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2634 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2635 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2636 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2637 cdac_sw_16_0.x3.ckb cdac_sw_16_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2638 x3[1].x3.ck x3[1].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2639 x3[0].x1.x10.A x3[0].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2640 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2641 cdac_sw_16_0.x1.x8.A cdac_sw_16_0.x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2642 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2643 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2644 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2645 vcn x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2646 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2647 vsref x2[0].x1.x8.A x2[0].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2648 vdref cdac_sw_16_0.x2.swp cdac_sw_16_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2649 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2650 vsref cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2651 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2652 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2653 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2654 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2655 cdac_sw_1_1.x3.ck cdac_sw_1_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2656 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2657 x4[2].x1.x10.A x4[2].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2658 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2659 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2660 vdref x4[3].x1.x9.A x4[3].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2661 x8[7].x3.ckb x8[7].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2662 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2663 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2664 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2665 vsref cdac_sw_4_1.x3.ckb cdac_sw_4_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2666 cdac_sw_2_1.x3.ckb cdac_sw_2_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2667 cdac_sw_8_0.x1.x8.A cdac_sw_8_0.x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2668 cdac_sw_4_1.x2.swn cdac_sw_4_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2669 vsref x10[8].x1.x10.A x10[8].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2670 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2671 a_127530_n8164# swp_in[2] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2672 cdac_sw_8_0.x3.ck cdac_sw_8_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2673 vsref x4[2].x1.x11.A x4[2].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2674 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2675 vdref cdac_sw_2_1.x1.x9.A cdac_sw_2_1.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2676 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2677 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2678 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2679 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2680 vdref x4[2].x1.x8.A x4[2].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2681 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2682 a_117284_n15188# cdac_sw_4_1.x3.ck x10b_cap_array_0.SW[4] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2683 x2[0].x3.ckb x2[0].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2684 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2685 vdref cdac_sw_8_1.x3.ckb cdac_sw_8_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2686 cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2687 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2688 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2689 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2690 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2691 a_105868_n6147# cdac_sw_1_2.x3.ckb cdac_sw_1_2.dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2692 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2693 x3[0].x3.ckb x3[0].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2694 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2695 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2696 cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2697 vsref cdac_sw_1_2.x1.x9.A cdac_sw_1_2.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2698 vcm cdac_sw_8_0.x2.swn x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2699 cdac_sw_2_1.x3.ck cdac_sw_2_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2700 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2701 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2702 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2703 x8[7].dac_out x8[7].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2704 a_129286_n15179# swn_in[8] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2705 a_104990_n5938# swp_in[9] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2706 a_131767_n4335# x3[1].x1.x8.A x3[1].x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2707 vdref x6[5].x1.x9.A x6[5].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2708 x10[8].x3.ck x10[8].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2709 x2[0].x1.x4.A x2[0].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2710 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2711 x4[2].x3.ckb x4[2].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2712 vdref cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2713 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2714 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2715 vsref cdac_sw_4_0.x3.ckb cdac_sw_4_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2716 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2717 cdac_sw_1_2.x2.swp cdac_sw_1_2.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2718 cdac_sw_1_0.x2.swp cdac_sw_1_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2719 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2720 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2721 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2722 vsref cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2723 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2724 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2725 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2726 x8[6].x3.ck x8[6].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2727 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2728 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2729 vsref cdac_sw_4_1.x2.swp cdac_sw_4_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2730 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2731 x3[0].x3.ckb x3[0].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2732 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2733 vsref cdac_sw_8_0.x3.ckb cdac_sw_8_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2734 x10[8].x3.ckb x10[8].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2735 vdref x3[1].x1.x11.A x3[1].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2736 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2737 x10b_cap_array_0.SW[2] cdac_sw_8_1.x3.ckb a_109966_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2738 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2739 vdref x3[1].x1.x9.A x3[1].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2740 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2741 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2742 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2743 vdref cdac_sw_1_2.x3.ckb cdac_sw_1_2.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2744 vdref cf[6] x8[6].x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2745 vdref x3[1].x2.swp x3[1].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2746 vsref swn_in[8] a_130164_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2747 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2748 vsref x10[8].x2.swp x10[8].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2749 x6[4].dac_out x6[4].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2750 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2751 cdac_sw_2_0.x3.ck cdac_sw_2_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2752 x8[7].x1.x10.A x8[7].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2753 vdref x3[0].x1.x10.A x3[0].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2754 a_109966_n15179# swn_in[2] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2755 vdref cdac_sw_16_0.x1.x9.A cdac_sw_16_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2756 cdac_sw_1_0.x1.x9.A cdac_sw_1_0.x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2757 vdref x6[5].x1.x11.A x6[5].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2758 vdref x3[1].x1.x6.A x3[1].x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2759 vdref swp_in[3] a_125188_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2760 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2761 cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2762 cdac_sw_1_0.x2.swn cdac_sw_1_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2763 vsref cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2764 x6[4].dac_out x6[4].x3.ck a_121090_n6892# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2765 vdref cdac_sw_1_1.x2.swp cdac_sw_1_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2766 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2767 a_111430_n6256# swp_in[7] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2768 a_110844_n15188# cdac_sw_8_1.x3.ck x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2769 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2770 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2771 vsref x8[7].x1.x11.A x8[7].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2772 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2773 vsref cdac_sw_1_1.x2.swp cdac_sw_1_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2774 x10[8].x3.ck x10[8].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2775 vdref x2[0].x3.ckb x2[0].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2776 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2777 vdref x8[7].x1.x8.A x8[7].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2778 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2779 vdref cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2780 cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2781 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2782 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2783 x3[0].x1.x10.A x3[0].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2784 cdac_sw_4_0.x2.swp cdac_sw_4_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2785 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2786 vdref x4[3].x1.x11.A x4[3].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2787 x10[8].x1.x10.A x10[8].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2788 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2789 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2790 cdac_sw_8_1.x2.swn cdac_sw_8_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2791 a_121090_n6892# swp_in[4] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2792 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2793 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2794 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2795 cdac_sw_16_0.x1.x3.Y cf[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2796 vsref x3[0].x3.ckb x3[0].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2797 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2798 cdac_sw_16_0.x2.swp cdac_sw_16_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2799 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2800 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2801 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2802 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2803 vdref swp_in[2] a_128408_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2804 a_126159_n16821# cdac_sw_2_0.x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2805 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2806 vdref x4[2].x1.x10.A x4[2].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2807 vsref x10[8].x1.x5.A x10[8].x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2808 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2809 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2810 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2811 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2812 x8[7].x3.ckb x8[7].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2813 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2814 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2815 vsref cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2816 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2817 x4[3].x1.x5.A x4[3].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2818 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2819 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2820 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2821 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2822 vsref cdac_sw_4_0.x1.x8.A cdac_sw_4_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2823 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2824 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2825 x4[2].x1.x10.A x4[2].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2826 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2827 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2828 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2829 cdac_sw_8_0.x1.x7.A cdac_sw_8_0.x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2830 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2831 x8[7].x3.ckb x8[7].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2832 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2833 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2834 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2835 cdac_sw_8_0.x1.x9.A cdac_sw_8_0.x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2836 a_128408_n9899# x4[2].x3.ckb x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2837 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2838 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2839 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2840 a_120504_n15188# cdac_sw_4_0.x3.ck x10b_cap_array_0.SW[5] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2841 vsref swn_in[7] a_126944_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2842 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2843 vcn x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2844 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2845 x3[1].x2.swn x3[1].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2846 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2847 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2848 vdref x8[6].x2.swp x8[6].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2849 x10b_cap_array_0.SW[4] cdac_sw_4_1.x3.ckb a_116406_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2850 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2851 vsref x4[2].x1.x8.A x4[2].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2852 vdref x3[0].x1.x8.A x3[0].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2853 vdref cdac_sw_8_1.x2.swp cdac_sw_8_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2854 vdref x6[5].x1.x9.A x6[5].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2855 cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2856 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2857 vsref x6[4].x1.x11.A x6[4].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2858 x10b_cap_array_0.SW[3] cdac_sw_8_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2859 cdac_sw_4_1.x3.ck cdac_sw_4_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2860 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2861 vdref x6[5].x3.ckb x6[5].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2862 vcp vcm sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2863 vsref x3[1].x2.swp x3[1].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2864 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2865 a_128408_n9899# x4[2].x3.ckb x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2866 a_130164_n15188# cdac_sw_1_1.x3.ck x10b_cap_array_0.SW[8] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2867 cdac_sw_2_1.x2.swn cdac_sw_2_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2868 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2869 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2870 a_110059_n15957# cdac_sw_8_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2871 cdac_sw_4_0.x3.ckb cdac_sw_4_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2872 vdref cdac_sw_8_0.x1.x8.A cdac_sw_8_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2873 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2874 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2875 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2876 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2877 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2878 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2879 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2880 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2881 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2882 vdref cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2883 x2[0].x1.x5.A x2[0].x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2884 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2885 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2886 x6[4].x2.swp x6[4].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2887 x4[2].x3.ckb x4[2].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2888 vdref cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2889 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2890 cdac_sw_8_1.x1.x3.Y cf[2] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2891 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2892 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2893 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2894 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2895 cdac_sw_16_0.x1.x5.A cdac_sw_16_0.x1.x8.A a_103619_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2896 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2897 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2898 vdref cdac_sw_1_2.x1.x9.A cdac_sw_1_2.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2899 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2900 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2901 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2902 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2903 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2904 x10[8].x2.swp x10[8].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2905 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2906 vdref x8[7].x1.x10.A x8[7].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2907 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2908 x3[0].x3.ckb x3[0].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2909 x10[8].x3.ckb x10[8].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2910 x3[0].x2.swn x3[0].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2911 vcm x4[3].x2.swp x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2912 vcm cdac_sw_4_0.x2.swn x10b_cap_array_0.SW[5] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2913 vsref x3[1].x1.x9.A a_131767_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2914 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2915 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2916 vsref cdac_sw_1_2.x3.ckb cdac_sw_1_2.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2917 vsref cdac_sw_1_1.x2.swp cdac_sw_1_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2918 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2919 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2920 vsref cdac_sw_4_1.x1.x8.A cdac_sw_4_1.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2921 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2922 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2923 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2924 x8[6].x2.swp x8[6].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2925 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2926 x8[7].x1.x10.A x8[7].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2927 vsref x3[0].x1.x10.A x3[0].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2928 vsref cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2929 x6[4].x2.swn x6[4].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2930 vsref x3[1].x1.x6.A x3[1].x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2931 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2932 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2933 vdref x3[0].x2.swp x3[0].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2934 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2935 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2936 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2937 a_112308_n6683# x8[7].x3.ckb x8[7].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2938 cdac_sw_8_1.x2.swn cdac_sw_8_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2939 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2940 vdref cf[8] x10[8].x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2941 cdac_sw_1_0.x1.x6.A cdac_sw_1_0.x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2942 x8[6].x2.swn x8[6].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2943 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2944 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2945 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2946 cdac_sw_1_0.x3.ckb cdac_sw_1_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2947 vdref x2[0].x2.swp x2[0].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2948 vsref x8[7].x1.x8.A x8[7].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2949 a_122939_n15957# cdac_sw_2_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2950 cdac_sw_16_0.x2.swp cdac_sw_16_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2951 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2952 vsref cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2953 vcp x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2954 vdref x4[2].x1.x10.A x4[2].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2955 vcm x4[2].x2.swp x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2956 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2957 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2958 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2959 vdref cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2960 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2961 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2962 x4[2].x1.x11.A x4[2].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2963 vdref cdac_sw_4_0.x3.ckb cdac_sw_4_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2964 cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2965 vsref x8[6].x2.swp x8[6].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2966 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2967 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2968 x2[0].x1.x10.A x2[0].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2969 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2970 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2971 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2972 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2973 vdref cdac_sw_1_2.x1.x8.A cdac_sw_1_2.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2974 vsref x4[2].x1.x10.A x4[2].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2975 vcm x6[4].x2.swp x6[4].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2976 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2977 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2978 x6[4].x1.x11.A x6[4].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2979 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2980 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2981 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2982 x8[7].x3.ckb x8[7].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2983 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2984 x3[1].x1.x4.A cf[1] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2985 cdac_sw_1_1.x2.swn cdac_sw_1_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2986 x3[1].x2.swn x3[1].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2987 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2988 x10[8].x2.swn x10[8].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2989 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2990 vdref cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2991 x10[8].x1.x11.A x10[8].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2992 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2993 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2994 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2995 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2996 cdac_sw_2_0.x1.x8.A cdac_sw_2_0.x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2997 vdref cf[6] cdac_sw_2_1.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2998 vsref cdac_sw_8_1.x2.swp cdac_sw_8_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2999 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3000 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3001 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3002 vcm cdac_sw_4_1.x2.swn x10b_cap_array_0.SW[4] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3003 vsref x10[8].x2.swp x10[8].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3004 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3005 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3006 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3007 vsref cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3008 vsref cdac_sw_2_0.x2.swp cdac_sw_2_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3009 cdac_sw_1_0.x2.swp cdac_sw_1_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3010 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3011 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3012 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3013 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3014 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3015 vsref cdac_sw_2_1.x3.ckb cdac_sw_2_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3016 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3017 vcm cdac_sw_8_0.x2.swn x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3018 cdac_sw_16_0.x1.x6.A cdac_sw_16_0.x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3019 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3020 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3021 vdref x3[0].x1.x11.A x3[0].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3022 vsref x3[0].x1.x8.A x3[0].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3023 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3024 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3025 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3026 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3027 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3028 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3029 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3030 vdref x10[8].x3.ckb x10[8].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3031 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3032 cdac_sw_1_2.x2.swn cdac_sw_1_2.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3033 cdac_sw_4_1.x2.swn cdac_sw_4_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3034 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3035 x2[0].x2.swn x2[0].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3036 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3037 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3038 vsref x6[5].x3.ckb x6[5].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3039 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3040 cdac_sw_1_1.x1.x6.A cdac_sw_1_1.x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3041 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3042 vdref cdac_sw_8_0.x1.x9.A cdac_sw_8_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3043 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3044 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3045 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3046 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3047 x3[0].x2.swp x3[0].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3048 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3049 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3050 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3051 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3052 vsref cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3053 cdac_sw_1_1.x3.ck cdac_sw_1_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3054 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3055 vsref cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3056 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3057 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3058 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3059 vdref x8[7].x1.x10.A x8[7].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3060 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3061 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3062 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3063 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3064 cdac_sw_2_1.x3.ckb cdac_sw_2_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3065 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3066 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3067 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3068 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3069 vdref cdac_sw_4_1.x3.ckb cdac_sw_4_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3070 cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3071 x8[7].x1.x11.A x8[7].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3072 vsref cdac_sw_1_2.x1.x9.A a_106007_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3073 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3074 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3075 vdref cdac_sw_1_2.x1.x5.A cdac_sw_1_2.x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3076 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3077 vcn x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3078 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3079 cdac_sw_2_1.x1.x3.Y cf[6] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3080 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3081 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3082 vsref x8[7].x1.x10.A x8[7].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3083 cdac_sw_8_0.x1.x3.Y cf[3] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3084 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3085 x8[6].x2.swp x8[6].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3086 cdac_sw_2_0.x2.swn cdac_sw_2_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3087 vsref cdac_sw_8_1.x3.ckb cdac_sw_8_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3088 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3089 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3090 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3091 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3092 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3093 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3094 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3095 vdref x10[8].x1.x4.A x10[8].x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3096 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3097 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3098 x4[2].x2.swp x4[2].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3099 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3100 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3101 vsref cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3102 cdac_sw_16_0.x2.swp cdac_sw_16_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3103 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3104 vdref cf[5] cdac_sw_4_0.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3105 vdref cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3106 x10b_cap_array_0.SW[3] cdac_sw_8_0.x3.ckb a_113186_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3107 a_114064_n15188# cdac_sw_8_0.x3.ck x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3108 vsref x2[0].x2.swp x2[0].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3109 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3110 x6[4].x2.swp x6[4].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3111 cdac_sw_1_0.x3.ck cdac_sw_1_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3112 x4[2].x2.swn x4[2].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3113 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3114 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3115 x3[1].x1.x11.A x3[1].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3116 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3117 vsref cdac_sw_1_1.x1.x8.A cdac_sw_1_1.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3118 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3119 cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3120 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3121 vdref x4[3].x1.x7.A x4[3].x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3122 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3123 x10b_cap_array_0.SW[2] cdac_sw_8_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3124 cdac_sw_2_0.x3.ckb cdac_sw_2_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3125 cdac_sw_1_0.x1.x7.A cdac_sw_1_0.x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3126 cdac_sw_2_1.x1.x7.A cdac_sw_2_1.x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3127 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3128 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3129 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3130 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3131 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3132 x10[8].x2.swp x10[8].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3133 vsref x4[2].x1.x10.A x4[2].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3134 x6[5].dac_out x6[5].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3135 cdac_sw_8_1.x3.ckb cdac_sw_8_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3136 x3[1].x3.ck x3[1].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3137 vdref x4[2].x2.swp x4[2].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3138 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3139 cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3140 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3141 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3142 x3[0].x2.swn x3[0].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3143 vdref cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3144 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3145 vdref cdac_sw_4_0.x2.swp cdac_sw_4_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3146 x2[0].x1.x11.A x2[0].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3147 vsref x3[0].x1.x11.A x3[0].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3148 vdref x6[4].x1.x10.A x6[4].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3149 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3150 vsref x10[8].x1.x11.A x10[8].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3151 cdac_sw_2_0.x3.ck cdac_sw_2_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3152 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3153 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3154 vsref cdac_sw_1_2.x1.x7.A cdac_sw_1_2.x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3155 vdref x3[1].x3.ckb x3[1].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3156 vsref cdac_sw_1_2.x1.x8.A cdac_sw_1_2.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3157 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3158 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3159 x10b_cap_array_0.SW[3] cdac_sw_8_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3160 cdac_sw_8_1.x3.ck cdac_sw_8_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3161 a_131767_n5199# cf[1] x3[1].x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3162 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3163 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3164 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3165 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3166 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3167 vsref x3[0].x1.x3.Y a_134987_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3168 vsref x10[8].x2.swp x10[8].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3169 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3170 x6[4].x3.ckb x6[4].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3171 vdref cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3172 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3173 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3174 cdac_sw_1_2.x2.swp cdac_sw_1_2.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3175 x4[2].dac_out x4[2].x3.ck a_127530_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3176 cdac_sw_4_0.x1.x3.Y cf[5] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3177 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3178 vcm x8[6].x2.swp x8[6].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3179 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3180 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3181 vdref x6[4].x2.swp x6[4].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3182 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3183 vdref cdac_sw_2_1.x1.x8.A cdac_sw_2_1.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3184 cdac_sw_8_0.x1.x5.A cdac_sw_8_0.x1.x8.A a_113279_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3185 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3186 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3187 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3188 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3189 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3190 vsref x2[0].x3.ckb x2[0].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3191 cdac_sw_8_0.x3.ckb cdac_sw_8_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3192 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3193 vsref swn_in[2] a_110844_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3194 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3195 cdac_sw_16_0.x3.ck cdac_sw_16_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3196 x10[8].x3.ckb x10[8].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3197 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3198 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3199 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3200 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3201 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3202 cdac_sw_16_0.x3.ck cdac_sw_16_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3203 vdref cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3204 x8[7].x2.swp x8[7].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3205 cdac_sw_16_0.x1.x7.A cdac_sw_16_0.x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3206 vsref cdac_sw_8_0.x1.x9.A cdac_sw_8_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3207 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3208 a_117870_n6892# swp_in[5] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3209 cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3210 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3211 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3212 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3213 vsref x10[8].x3.ckb x10[8].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3214 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3215 vsref cdac_sw_2_0.x1.x8.A cdac_sw_2_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3216 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3217 x8[7].x2.swn x8[7].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3218 vdref x4[2].x1.x9.A x4[2].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3219 cdac_sw_1_1.x1.x7.A cdac_sw_1_1.x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3220 x8[6].x3.ckb x8[6].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3221 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3222 cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3223 vdref cdac_sw_2_0.x3.ckb cdac_sw_2_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3224 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3225 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3226 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3227 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3228 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3229 vsref cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3230 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3231 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3232 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3233 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3234 x2[0].x3.ckb x2[0].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3235 cdac_sw_1_1.x2.swn cdac_sw_1_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3236 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3237 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3238 cdac_sw_4_0.x2.swn cdac_sw_4_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3239 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3240 a_113186_n15179# swn_in[3] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3241 vsref x8[7].x1.x10.A x8[7].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3242 x8[6].x3.ck x8[6].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3243 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3244 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3245 vdref x8[7].x2.swp x8[7].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3246 vsref swn_in[3] a_114064_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3247 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3248 x2[0].x3.ck x2[0].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3249 vdref cdac_sw_4_1.x2.swp cdac_sw_4_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3250 cdac_sw_2_1.x2.swp cdac_sw_2_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3251 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3252 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3253 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3254 vsref swn_in[5] a_120504_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3255 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3256 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3257 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3258 vsref x3[0].x1.x9.A x3[0].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3259 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3260 vsref x10[8].x1.x9.A x10[8].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3261 x4[2].x2.swp x4[2].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3262 x2[0].x3.ck x2[0].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3263 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3264 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3265 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3266 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3267 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3268 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3269 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3270 vsref x6[5].x2.swp x6[5].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3271 vdref x8[6].x3.ckb x8[6].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3272 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3273 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3274 x6[4].x1.x10.A x6[4].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3275 vsref x10[8].x1.x4.A x10[8].x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3276 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3277 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3278 cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3279 vdref x4[2].x1.x11.A x4[2].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3280 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3281 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3282 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3283 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3284 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3285 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3286 x3[0].x2.swp x3[0].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3287 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3288 vdref cdac_sw_4_0.x1.x8.A cdac_sw_4_0.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3289 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3290 vsref cdac_sw_1_2.x1.x10.A cdac_sw_1_2.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3291 x10[8].x3.ck x10[8].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3292 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3293 vcn x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3294 vdref cdac_sw_1_2.x2.swp cdac_sw_1_2.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3295 vdref cdac_sw_8_0.x3.ckb cdac_sw_8_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3296 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3297 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3298 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3299 x10[8].x1.x10.A x10[8].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3300 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3301 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3302 vdref x3[0].x1.x11.A x3[0].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3303 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3304 vdref x2[0].x1.x10.A x2[0].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3305 vdref cf[9] cdac_sw_1_0.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3306 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3307 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3308 vsref cdac_sw_4_0.x2.swp cdac_sw_4_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3309 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3310 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3311 x2[0].x1.x11.A x2[0].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3312 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3313 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3314 vdref x6[5].x1.x3.Y x6[5].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3315 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3316 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3317 vdref x10[8].x3.ckb x10[8].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3318 cdac_sw_8_1.x2.swp cdac_sw_8_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3319 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3320 vsref x8[7].x2.swp x8[7].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3321 x3[1].x3.ck x3[1].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3322 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3323 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3324 vsref cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3325 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3326 vsref cdac_sw_1_0.x3.ckb cdac_sw_1_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3327 vdref cdac_sw_1_0.x1.x8.A cdac_sw_1_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3328 cdac_sw_8_1.x2.swp cdac_sw_8_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3329 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3330 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3331 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3332 vdref x8[7].x1.x9.A x8[7].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3333 x4[3].dac_out x4[3].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3334 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3335 vdref x6[5].x1.x7.A x6[5].x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3336 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3337 vsref x6[4].x1.x10.A x6[4].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3338 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3339 cdac_sw_2_0.x2.swn cdac_sw_2_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3340 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3341 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3342 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3343 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3344 vsref x8[6].x1.x11.A x8[6].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3345 vsref x3[1].x3.ckb x3[1].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3346 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3347 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3348 cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3349 vsref cf[3] x4[3].x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3350 x10b_cap_array_0.SW[2] cdac_sw_8_1.x3.ckb a_109966_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3351 x4[3].dac_out x4[3].x3.ck a_124310_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3352 vsref cdac_sw_4_1.x3.ckb cdac_sw_4_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3353 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3354 vsref swn_in[4] a_117284_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3355 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3356 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3357 x6[4].x3.ckb x6[4].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3358 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3359 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3360 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3361 vsref cdac_sw_8_1.x1.x8.A cdac_sw_8_1.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3362 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3363 a_109966_n15179# swn_in[2] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3364 cdac_sw_1_0.x3.ckb cdac_sw_1_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3365 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3366 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3367 vdref x3[1].x1.x9.A x3[1].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3368 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3369 cdac_sw_16_0.x1.x9.A cdac_sw_16_0.x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3370 x10[8].x3.ckb x10[8].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3371 cdac_sw_1_0.x1.x3.Y cf[9] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3372 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3373 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3374 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3375 vsref x2[0].x1.x9.A x2[0].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3376 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3377 x8[6].x3.ckb x8[6].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3378 x10b_cap_array_0.SW[3] cdac_sw_8_0.x3.ckb a_113186_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3379 cdac_sw_16_0.x2.swn cdac_sw_16_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3380 vdref cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3381 vdref x8[7].x1.x11.A x8[7].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3382 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3383 vcm cdac_sw_8_1.x2.swn x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3384 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3385 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3386 x4[2].dac_out x4[2].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3387 cdac_sw_1_1.x2.swn cdac_sw_1_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3388 a_106007_n4335# cdac_sw_1_2.x1.x8.A cdac_sw_1_2.x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3389 x10b_cap_array_0.SW[2] cdac_sw_8_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3390 x2[0].x3.ck x2[0].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3391 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3392 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3393 x8[6].x3.ckb x8[6].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3394 vdref cdac_sw_16_0.x1.x8.A cdac_sw_16_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3395 vdref cf[8] cdac_sw_1_1.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3396 vdref cdac_sw_2_0.x2.swp cdac_sw_2_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3397 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3398 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3399 a_124310_n8164# swp_in[3] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3400 vsref cdac_sw_4_1.x2.swp cdac_sw_4_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3401 cdac_sw_2_1.x2.swp cdac_sw_2_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3402 x6[4].x3.ckb x6[4].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3403 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3404 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3405 cdac_sw_1_2.x2.swp cdac_sw_1_2.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3406 cdac_sw_8_0.x2.swn cdac_sw_8_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3407 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3408 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3409 x2[0].x2.swp x2[0].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3410 vdref swp_in[2] a_128408_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3411 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3412 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3413 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3414 x8[6].x3.ck x8[6].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3415 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3416 x2[0].x2.swp x2[0].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3417 x2[0].x2.swn x2[0].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3418 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3419 cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3420 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3421 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3422 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3423 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3424 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3425 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3426 x10[8].x3.ckb x10[8].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3427 vdref x3[1].x1.x11.A x3[1].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3428 cdac_sw_4_0.x3.ckb cdac_sw_4_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3429 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3430 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3431 vdref cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3432 vdref cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3433 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3434 vdref x3[1].x2.swp x3[1].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3435 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3436 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3437 cdac_sw_4_0.x3.ck cdac_sw_4_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3438 vsref x8[6].x3.ckb x8[6].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3439 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3440 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3441 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3442 vdref x3[0].x1.x10.A x3[0].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3443 a_128408_n9899# x4[2].x3.ckb x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3444 vdref x10[8].x1.x10.A x10[8].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3445 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3446 vdref cdac_sw_1_2.x1.x6.A cdac_sw_1_2.x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3447 cdac_sw_8_0.x3.ckb cdac_sw_8_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3448 x6[4].x1.x10.A x6[4].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3449 cdac_sw_4_0.x3.ck cdac_sw_4_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3450 vsref cdac_sw_4_0.x2.swp cdac_sw_4_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3451 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3452 x3[1].x2.swn x3[1].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3453 vsref x2[0].x1.x8.A x2[0].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3454 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3455 vdref x3[0].x1.x9.A x3[0].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3456 vdref cf[5] x6[5].x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3457 a_127530_n8164# swp_in[2] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3458 vsref cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3459 vdref x10[8].x3.ckb x10[8].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3460 x10[8].x3.ck x10[8].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3461 vdref cdac_sw_8_0.x2.swp cdac_sw_8_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3462 vsref cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3463 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3464 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3465 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3466 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3467 x10[8].x1.x10.A x10[8].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3468 cdac_sw_1_1.x1.x3.Y cf[8] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3469 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3470 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3471 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3472 vsref x6[4].x1.x5.A x6[4].x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3473 a_117284_n15188# cdac_sw_4_1.x3.ck x10b_cap_array_0.SW[4] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3474 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3475 vsref cdac_sw_8_0.x2.swp cdac_sw_8_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3476 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3477 vdref x2[0].x1.x11.A x2[0].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3478 vdref cdac_sw_1_0.x1.x8.A cdac_sw_1_0.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3479 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3480 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3481 cdac_sw_2_1.x3.ckb cdac_sw_2_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3482 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3483 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3484 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3485 vsref x10[8].x3.ckb x10[8].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3486 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3487 cdac_sw_2_1.x1.x8.A cdac_sw_2_1.x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3488 vcm cdac_sw_8_0.x2.swn x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3489 cdac_sw_2_0.x2.swn cdac_sw_2_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3490 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3491 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3492 cdac_sw_2_1.x3.ck cdac_sw_2_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3493 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3494 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3495 x8[7].dac_out x8[7].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3496 vdref cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3497 vdref cdac_sw_1_0.x1.x9.A cdac_sw_1_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3498 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3499 cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3500 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3501 vcp x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3502 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3503 cdac_sw_4_1.x3.ckb cdac_sw_4_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3504 a_113186_n15179# swn_in[3] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3505 vsref cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3506 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3507 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3508 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3509 cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3510 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3511 x6[5].x2.swn x6[5].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3512 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3513 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3514 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3515 x10b_cap_array_0.SW[5] cdac_sw_4_0.x3.ckb a_119626_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3516 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3517 vdref cdac_sw_1_2.x1.x9.A cdac_sw_1_2.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3518 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3519 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3520 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3521 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3522 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3523 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3524 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3525 cdac_sw_4_1.x1.x4.A cdac_sw_4_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3526 cdac_sw_2_0.x3.ckb cdac_sw_2_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3527 x4[2].dac_out x4[2].x3.ck a_127530_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3528 cdac_sw_1_0.x2.swp cdac_sw_1_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3529 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3530 vdref x8[6].x2.swp x8[6].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3531 vsref cdac_sw_1_1.x3.ckb cdac_sw_1_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3532 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3533 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3534 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3535 vdref x3[0].x1.x8.A x3[0].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3536 vdref x10[8].x1.x8.A x10[8].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3537 cdac_sw_4_1.x3.ck cdac_sw_4_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3538 vsref cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3539 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3540 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3541 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3542 a_112308_n6683# x8[7].x3.ckb x8[7].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3543 a_122846_n15179# swn_in[6] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3544 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3545 x8[6].x3.ckb x8[6].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3546 vsref cdac_sw_8_0.x3.ckb cdac_sw_8_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3547 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3548 vdref x6[5].x3.ckb x6[5].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3549 x8[6].x2.swn x8[6].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3550 x6[5].x1.x5.A x6[5].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3551 cdac_sw_8_1.x3.ck cdac_sw_8_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3552 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3553 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3554 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3555 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3556 x8[7].x2.swn x8[7].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3557 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3558 vsref x2[0].x1.x10.A x2[0].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3559 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3560 a_111430_n6256# swp_in[7] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3561 vcm x4[2].x2.swp x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3562 x2[0].x2.swn x2[0].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3563 vsref cdac_sw_4_0.x1.x9.A cdac_sw_4_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3564 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3565 a_114064_n15188# cdac_sw_8_0.x3.ck x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3566 cdac_sw_16_0.x3.ckb cdac_sw_16_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3567 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3568 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3569 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3570 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3571 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3572 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3573 x6[4].x2.swp x6[4].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3574 vdref cdac_sw_16_0.x1.x9.A cdac_sw_16_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3575 vdref cdac_sw_1_1.x1.x8.A cdac_sw_1_1.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3576 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3577 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3578 x6[4].x3.ckb x6[4].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3579 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3580 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3581 vcm x6[4].x2.swp x6[4].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3582 vdref cdac_sw_2_1.x3.ckb cdac_sw_2_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3583 vdref x10[8].x2.swp x10[8].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3584 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3585 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3586 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3587 cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3588 cdac_sw_4_0.x3.ck cdac_sw_4_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3589 a_126066_n15179# swn_in[7] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3590 a_119719_n15957# cdac_sw_4_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3591 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3592 vdref cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3593 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3594 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3595 cdac_sw_8_0.x3.ckb cdac_sw_8_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3596 cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3597 cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3598 vsref x8[6].x1.x11.A x8[6].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3599 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3600 x10[8].x3.ckb x10[8].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3601 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3602 cdac_sw_4_0.x2.swp cdac_sw_4_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3603 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3604 vdref x8[7].x3.ckb x8[7].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3605 x3[0].x2.swn x3[0].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3606 vdref cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3607 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3608 x10[8].x2.swn x10[8].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3609 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3610 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3611 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3612 vdref cf[4] x6[4].x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3613 cdac_sw_4_0.x2.swn cdac_sw_4_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3614 a_110059_n16821# cdac_sw_8_1.x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3615 cdac_sw_4_0.x2.swp cdac_sw_4_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3616 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3617 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3618 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3619 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3620 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3621 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3622 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3623 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3624 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3625 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3626 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3627 vsref x10[8].x1.x10.A x10[8].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3628 vsref x3[0].x1.x10.A x3[0].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3629 cdac_sw_8_0.x2.swp cdac_sw_8_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3630 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3631 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3632 vdref x8[6].x1.x10.A x8[6].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3633 vsref cdac_sw_1_2.x1.x6.A cdac_sw_1_2.x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3634 x8[6].x2.swn x8[6].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3635 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3636 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3637 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3638 vsref cdac_sw_2_0.x3.ckb cdac_sw_2_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3639 vsref x3[0].x1.x9.A a_134987_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3640 vsref swn_in[7] a_126944_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3641 vdref x3[0].x1.x5.A x3[0].x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3642 vsref x10[8].x3.ckb x10[8].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3643 vdref swp_in[2] a_128408_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3644 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3645 vsref cdac_sw_4_0.x1.x8.A cdac_sw_4_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3646 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3647 vsref swn_in[2] a_110844_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3648 a_119626_n15179# swn_in[5] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3649 cdac_sw_4_1.x3.ckb cdac_sw_4_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3650 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3651 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3652 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3653 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3654 cdac_sw_2_1.x1.x9.A cdac_sw_2_1.x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3655 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3656 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3657 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3658 vdref cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3659 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3660 vsref cdac_sw_4_1.x1.x9.A cdac_sw_4_1.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3661 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3662 x10b_cap_array_0.SW[6] cdac_sw_2_1.x3.ckb a_122846_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3663 vdref cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3664 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3665 x6[4].x1.x11.A x6[4].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3666 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3667 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3668 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3669 vsref x8[6].x1.x5.A x8[6].x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3670 a_128408_n9899# x4[2].x3.ckb x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3671 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3672 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3673 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3674 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3675 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3676 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3677 cdac_sw_1_2.x1.x4.A cf[9] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3678 x3[1].x2.swn x3[1].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3679 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3680 x3[0].x1.x11.A x3[0].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3681 cdac_sw_4_1.x3.ck cdac_sw_4_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3682 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3683 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3684 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3685 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3686 cdac_sw_1_0.x2.swp cdac_sw_1_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3687 a_122939_n16821# cdac_sw_2_1.x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3688 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3689 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3690 cdac_sw_1_1.x3.ckb cdac_sw_1_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3691 vsref cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3692 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3693 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3694 cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3695 cdac_sw_2_0.x1.x3.Y cf[7] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3696 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3697 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3698 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3699 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3700 vcm cdac_sw_8_0.x2.swn x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3701 cdac_sw_4_1.x1.x5.A cdac_sw_4_1.x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3702 cdac_sw_2_0.x2.swp cdac_sw_2_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3703 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3704 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3705 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3706 cdac_sw_1_2.dac_out cdac_sw_1_2.x3.ck a_104990_n5938# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3707 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3708 x10b_cap_array_0.SW[3] cdac_sw_8_0.x3.ckb a_113186_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3709 x8[6].x1.x11.A x8[6].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3710 vdref x10[8].x1.x11.A x10[8].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3711 vsref x3[0].x1.x8.A x3[0].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3712 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3713 vsref x3[0].x1.x7.A x3[0].x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3714 vsref x10[8].x1.x8.A x10[8].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3715 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3716 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3717 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3718 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3719 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3720 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3721 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3722 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3723 x10b_cap_array_0.SW[2] cdac_sw_8_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3724 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3725 vsref x6[5].x3.ckb x6[5].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3726 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3727 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3728 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3729 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3730 x3[0].x2.swp x3[0].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3731 vsref x8[6].x1.x9.A x8[6].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3732 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3733 x3[1].x2.swp x3[1].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3734 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3735 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3736 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3737 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3738 cdac_sw_2_0.x1.x9.A cdac_sw_2_0.x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3739 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3740 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3741 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3742 vdref cdac_sw_4_1.x3.ckb cdac_sw_4_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3743 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3744 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3745 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3746 vdref cdac_sw_2_1.x2.swp cdac_sw_2_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3747 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3748 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3749 x10[8].x2.swn x10[8].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3750 vdref swp_in[8] a_109088_n6147# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3751 cdac_sw_4_0.x2.swn cdac_sw_4_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3752 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3753 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3754 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3755 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3756 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3757 vdref x6[4].x1.x4.A x6[4].x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3758 vsref cdac_sw_2_1.x2.swp cdac_sw_2_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3759 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3760 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3761 vdref cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3762 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3763 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3764 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3765 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3766 cdac_sw_8_0.x2.swp cdac_sw_8_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3767 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3768 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3769 x8[6].x2.swp x8[6].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3770 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3771 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3772 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3773 cdac_sw_1_0.x1.x8.A cdac_sw_1_0.x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3774 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3775 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3776 vsref x8[7].x3.ckb x8[7].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3777 vcn x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3778 x4[2].dac_out x4[2].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3779 a_132599_n15957# cdac_sw_1_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3780 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3781 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3782 vsref x3[1].x2.swp x3[1].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3783 x6[4].dac_out x6[4].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3784 cdac_sw_1_0.x3.ck cdac_sw_1_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3785 x8[6].x2.swn x8[6].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3786 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3787 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3788 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3789 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3790 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3791 vdref cdac_sw_1_1.x3.ckb cdac_sw_1_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3792 vsref cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3793 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3794 vcm x4[2].x2.swp x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3795 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3796 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3797 x6[4].x2.swp x6[4].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3798 x6[4].dac_out x6[4].x3.ck a_121090_n6892# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3799 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3800 cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3801 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3802 vsref x8[6].x1.x10.A x8[6].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3803 x6[5].x3.ck x6[5].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3804 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3805 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3806 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3807 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3808 cdac_sw_8_1.x1.x8.A cdac_sw_8_1.x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3809 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3810 vdref swp_in[4] a_121968_n7755# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3811 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3812 a_121090_n6892# swp_in[4] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3813 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3814 x10[8].x2.swp x10[8].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3815 vsref x6[4].x1.x11.A x6[4].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3816 cdac_sw_2_0.x1.x4.A cdac_sw_2_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3817 vcm x6[5].x2.swp x6[5].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3818 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3819 vsref cdac_sw_8_1.x2.swp cdac_sw_8_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3820 x10[8].x2.swn x10[8].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3821 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3822 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3823 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3824 x3[0].x1.x11.A x3[0].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3825 vsref cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3826 vdref cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3827 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3828 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3829 vsref x6[4].x2.swp x6[4].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3830 x10[8].x1.x11.A x10[8].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3831 vsref cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3832 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3833 vsref x10[8].x1.x11.A x10[8].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3834 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3835 a_113186_n15179# swn_in[3] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3836 cdac_sw_1_1.x3.ckb cdac_sw_1_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3837 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3838 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3839 x8[6].x2.swp x8[6].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3840 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3841 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3842 cdac_sw_1_0.x2.swn cdac_sw_1_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3843 x8[7].x3.ck x8[7].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3844 vdref x3[0].x2.swp x3[0].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3845 cdac_sw_8_0.x1.x6.A cdac_sw_8_0.x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3846 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3847 a_127530_n8164# swp_in[2] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3848 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3849 vsref cf[0] x3[0].x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3850 a_106007_n5199# cf[9] cdac_sw_1_2.x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3851 cdac_sw_4_1.x2.swn cdac_sw_4_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3852 vsref cdac_sw_1_1.x1.x9.A cdac_sw_1_1.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3853 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3854 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3855 vsref x10[8].x1.x3.Y a_109227_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3856 a_123724_n15188# cdac_sw_2_1.x3.ck x10b_cap_array_0.SW[6] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3857 cdac_sw_2_0.x2.swp cdac_sw_2_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3858 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3859 x6[4].x3.ckb x6[4].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3860 vsref cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3861 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3862 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3863 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3864 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3865 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3866 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3867 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3868 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3869 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3870 cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3871 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3872 a_129379_n15957# cdac_sw_1_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3873 cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3874 x4[2].x1.x11.A x4[2].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3875 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3876 vsref x8[6].x2.swp x8[6].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3877 vdref x8[6].x1.x10.A x8[6].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3878 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3879 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3880 x8[7].x2.swp x8[7].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3881 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3882 vcp x3[0].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3883 cdac_sw_8_1.x2.swn cdac_sw_8_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3884 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3885 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3886 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3887 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3888 vsref x4[2].x1.x3.Y a_128547_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3889 a_114064_n15188# cdac_sw_8_0.x3.ck x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3890 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3891 vdref x4[2].x1.x9.A x4[2].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3892 cdac_sw_4_1.x1.x6.A cdac_sw_4_1.x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3893 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3894 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3895 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3896 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3897 vcm x10[8].x2.swp x10[8].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3898 vsref cdac_sw_4_0.x3.ckb cdac_sw_4_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3899 vdref cf[0] cdac_sw_16_0.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3900 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3901 vsref x6[4].x1.x9.A x6[4].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3902 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3903 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3904 vsref x4[2].x1.x7.A x4[2].x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3905 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3906 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3907 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3908 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3909 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3910 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3911 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3912 vdref cdac_sw_4_1.x2.swp cdac_sw_4_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3913 vsref x2[0].x2.swp x2[0].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3914 cdac_sw_8_0.x2.swp cdac_sw_8_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3915 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3916 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3917 cdac_sw_8_1.x3.ckb cdac_sw_8_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3918 cdac_sw_1_0.x3.ck cdac_sw_1_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3919 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3920 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3921 a_109088_n6147# x10[8].x3.ckb x10[8].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3922 vsref cdac_sw_16_0.x3.ckb cdac_sw_16_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3923 cdac_sw_16_0.x2.swn cdac_sw_16_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3924 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3925 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3926 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3927 x4[2].x2.swp x4[2].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3928 vsref x6[4].x1.x4.A x6[4].x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3929 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3930 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3931 vsref x10[8].x1.x9.A x10[8].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3932 cdac_sw_2_0.x3.ckb cdac_sw_2_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3933 vdref cdac_sw_1_1.x3.ckb cdac_sw_1_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3934 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3935 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3936 x8[6].dac_out x8[6].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3937 x10b_cap_array_0.SW[2] cdac_sw_8_1.x3.ckb a_109966_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3938 x10b_cap_array_0.SW[3] cdac_sw_8_0.x3.ckb a_113186_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3939 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3940 vcm cdac_sw_4_0.x2.swn x10b_cap_array_0.SW[5] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3941 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3942 cdac_sw_1_0.x1.x9.A cdac_sw_1_0.x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3943 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3944 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3945 a_134987_n4335# x3[0].x1.x8.A x3[0].x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3946 vdref cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3947 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3948 vsref cdac_sw_2_0.x1.x9.A cdac_sw_2_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3949 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3950 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3951 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3952 x6[4].x1.x10.A x6[4].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3953 x10b_cap_array_0.SW[2] cdac_sw_8_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3954 cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3955 a_109966_n15179# swn_in[2] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3956 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3957 vsref x2[0].x1.x10.A x2[0].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3958 cdac_sw_8_1.x3.ck cdac_sw_8_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3959 vdref x8[6].x1.x4.A x8[6].x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3960 x10[8].x2.swp x10[8].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3961 x3[0].x2.swp x3[0].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3962 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3963 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3964 x2[0].x1.x4.A cf[1] a_106839_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3965 vdref cdac_sw_1_1.x2.swp cdac_sw_1_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3966 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3967 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3968 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3969 vsref swn_in[3] a_114064_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3970 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3971 vdref x3[1].x1.x3.Y x3[1].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3972 cdac_sw_16_0.x3.ckb cdac_sw_16_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3973 cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3974 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3975 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3976 vsref x4[3].x2.swp x4[3].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3977 vdref cdac_sw_1_2.x2.swp cdac_sw_1_2.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3978 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3979 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3980 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3981 x6[5].x3.ck x6[5].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3982 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3983 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3984 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3985 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3986 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3987 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3988 x8[7].x1.x11.A x8[7].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3989 vdref x3[0].x1.x11.A x3[0].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3990 vsref swn_in[2] a_110844_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3991 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3992 cdac_sw_16_0.x1.x3.Y cf[0] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3993 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3994 vdref x3[1].x1.x7.A x3[1].x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3995 cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3996 a_121968_n7755# x6[4].x3.ckb x6[4].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3997 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3998 x2[0].x2.swn x2[0].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3999 vsref cdac_sw_1_0.x3.ckb cdac_sw_1_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4000 cdac_sw_2_0.x1.x5.A cdac_sw_2_0.x1.x3.Y vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4001 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4002 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4003 x4[3].x2.swn x4[3].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4004 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4005 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4006 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4007 x4[3].dac_out x4[3].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4008 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4009 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4010 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4011 vsref x8[7].x1.x3.Y a_112447_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4012 x8[6].x1.x10.A x8[6].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4013 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4014 vdref swp_in[2] a_128408_n9899# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4015 vsref cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4016 vdref x8[7].x1.x9.A x8[7].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4017 vdref x3[0].x1.x6.A x3[0].x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4018 cdac_sw_1_1.x3.ck cdac_sw_1_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4019 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4020 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4021 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4022 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4023 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4024 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4025 x4[3].dac_out x4[3].x3.ck a_124310_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4026 cdac_sw_8_0.x3.ck cdac_sw_8_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4027 a_114650_n6256# swp_in[6] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4028 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4029 vsref x8[6].x1.x11.A x8[6].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4030 vsref cdac_sw_8_1.x1.x8.A cdac_sw_8_1.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4031 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4032 x8[7].x3.ck x8[7].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4033 cdac_sw_8_0.x1.x7.A cdac_sw_8_0.x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4034 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4035 vdref x8[6].x1.x8.A x8[6].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4036 x2[0].x3.ckb x2[0].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4037 vdref cdac_sw_8_1.x3.ckb cdac_sw_8_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4038 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4039 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4040 x3[1].x3.ckb x3[1].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4041 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4042 vdref x4[2].x1.x11.A x4[2].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4043 x6[4].x3.ckb x6[4].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4044 vdref cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4045 vdref cdac_sw_2_0.x3.ckb cdac_sw_2_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4046 cdac_sw_1_0.x3.ckb cdac_sw_1_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4047 x8[7].x2.swp x8[7].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4048 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4049 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4050 a_128408_n9899# x4[2].x3.ckb x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4051 vcm cdac_sw_4_1.x2.swn x10b_cap_array_0.SW[4] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4052 cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4053 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4054 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4055 vsref cdac_sw_1_0.x2.swp cdac_sw_1_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4056 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4057 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4058 x2[0].x3.ck x2[0].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4059 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4060 x8[6].x3.ckb x8[6].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4061 vsref x8[6].x1.x10.A x8[6].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4062 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4063 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4064 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4065 vsref x10[8].x1.x11.A x10[8].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4066 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4067 vdref x3[1].x3.ckb x3[1].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4068 a_113186_n15179# swn_in[3] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4069 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4070 a_124310_n8164# swp_in[3] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4071 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4072 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4073 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4074 vsref cdac_sw_4_1.x2.swp cdac_sw_4_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4075 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4076 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4077 vdref x3[0].x1.x9.A x3[0].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4078 x6[4].x3.ckb x6[4].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4079 vdref cdac_sw_16_0.x1.x8.A cdac_sw_16_0.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4080 cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4081 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4082 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4083 vsref cdac_sw_8_1.x1.x9.A cdac_sw_8_1.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4084 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4085 vdref x6[5].x2.swp x6[5].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4086 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4087 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4088 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4089 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4090 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4091 cdac_sw_2_0.x3.ck cdac_sw_2_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4092 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4093 a_109227_n4335# x10[8].x1.x8.A x10[8].x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4094 x10[8].x3.ckb x10[8].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4095 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4096 vdref x6[4].x1.x10.A x6[4].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4097 vcm cdac_sw_8_1.x2.swn x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4098 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4099 vsref x4[3].x1.x11.A x4[3].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4100 vdref cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4101 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4102 vdref cdac_sw_1_1.x2.swp cdac_sw_1_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4103 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4104 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4105 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4106 cdac_sw_16_0.x3.ckb cdac_sw_16_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4107 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4108 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4109 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4110 vdref cf[1] x3[1].x1.x3.Y vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4111 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4112 vdref x6[4].x3.ckb x6[4].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4113 x10b_cap_array_0.SW[5] cdac_sw_4_0.x3.ckb a_119626_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4114 vdref x2[0].x3.ckb x2[0].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4115 vdref cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4116 vdref cdac_sw_1_2.x1.x3.Y cdac_sw_1_2.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4117 vdref x10[8].x1.x10.A x10[8].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4118 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4119 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4120 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4121 x6[4].x1.x10.A x6[4].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4122 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4123 x8[6].x3.ckb x8[6].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4124 cdac_sw_8_1.x2.swn cdac_sw_8_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4125 vdref x8[7].x1.x11.A x8[7].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4126 vsref x8[6].x1.x4.A x8[6].x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4127 cdac_sw_2_1.x1.x6.A cdac_sw_2_1.x1.x4.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4128 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4129 vdref x10[8].x1.x9.A x10[8].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4130 cdac_sw_16_0.x2.swp cdac_sw_16_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4131 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4132 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4133 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4134 x4[3].x2.swn x4[3].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4135 a_128547_n4335# x4[2].x1.x8.A x4[2].x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4136 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4137 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4138 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4139 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4140 x6[5].dac_out x6[5].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4141 vcm x4[2].x2.swp x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4142 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4143 cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4144 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4145 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4146 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4147 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4148 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4149 vdref x8[6].x3.ckb x8[6].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4150 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4151 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4152 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4153 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4154 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4155 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4156 x8[6].x1.x10.A x8[6].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4157 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4158 vsref x3[0].x1.x6.A x3[0].x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4159 vcm x6[4].x2.swp x6[4].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4160 cdac_sw_1_1.x2.swn cdac_sw_1_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4161 vdref x4[2].x1.x11.A x4[2].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4162 cdac_sw_4_0.x2.swn cdac_sw_4_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4163 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4164 vsref x4[3].x1.x5.A x4[3].x1.x7.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4165 vsref x2[0].x1.x9.A x2[0].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4166 a_115528_n6683# x8[6].x3.ckb x8[6].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4167 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4168 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4169 vdref x4[2].x1.x9.A x4[2].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4170 cdac_sw_2_0.x1.x6.A cdac_sw_2_0.x1.x4.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4171 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4172 x6[5].x2.swn x6[5].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4173 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4174 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4175 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4176 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4177 vdref cf[3] cdac_sw_8_0.x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4178 vdref cdac_sw_8_1.x2.swp cdac_sw_8_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4179 vsref cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4180 vsref x8[6].x1.x8.A x8[6].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4181 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4182 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4183 vdref x6[4].x1.x8.A x6[4].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4184 x3[1].x3.ckb x3[1].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4185 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4186 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4187 vdref cdac_sw_1_2.x1.x9.A cdac_sw_1_2.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4188 vdref x4[2].x1.x6.A x4[2].x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4189 x4[2].dac_out x4[2].x3.ck a_127530_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4190 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4191 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4192 x10b_cap_array_0.SW[5] cdac_sw_4_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4193 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4194 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4195 vdref cdac_sw_16_0.x1.x11.A cdac_sw_16_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4196 vdref cdac_sw_2_0.x2.swp cdac_sw_2_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4197 cdac_sw_1_0.x2.swp cdac_sw_1_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4198 cdac_sw_2_1.x2.swp cdac_sw_2_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4199 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4200 x6[5].dac_out x6[5].x3.ck a_117870_n6892# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4201 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4202 cdac_sw_4_0.x3.ckb cdac_sw_4_0.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4203 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4204 vsref x6[5].x2.swp x6[5].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4205 x3[1].x1.x5.A x3[1].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4206 vdref cdac_sw_8_0.x1.x8.A cdac_sw_8_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4207 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4208 vcn x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4209 cdac_sw_1_2.dac_out cdac_sw_1_2.x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4210 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4211 x4[3].x2.swn x4[3].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4212 cdac_sw_8_1.x1.x10.A cdac_sw_8_1.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4213 cdac_sw_2_1.x2.swn cdac_sw_2_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4214 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4215 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4216 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4217 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4218 vdref x10[8].x1.x8.A x10[8].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4219 vsref swn_in[1] a_107624_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4220 x4[3].x1.x11.A x4[3].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4221 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4222 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4223 x2[0].x2.swn x2[0].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4224 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4225 x8[6].x3.ckb x8[6].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4226 a_117870_n6892# swp_in[5] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4227 cdac_sw_4_1.x2.swp cdac_sw_4_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4228 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4229 x3[0].x1.x4.A cf[0] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4230 x10b_cap_array_0.SW[2] cdac_sw_8_1.x3.ckb a_109966_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4231 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4232 vdref cdac_sw_1_0.x1.x10.A cdac_sw_1_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4233 x8[7].x2.swn x8[7].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4234 vsref x3[1].x3.ckb x3[1].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4235 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4236 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4237 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4238 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4239 cdac_sw_4_0.x3.ck cdac_sw_4_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4240 a_119626_n15179# swn_in[5] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4241 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4242 a_112447_n4335# x8[7].x1.x8.A x8[7].x1.x5.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4243 a_109966_n15179# swn_in[2] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4244 a_110844_n15188# cdac_sw_8_1.x3.ck x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4245 cdac_sw_4_1.x1.x4.A cf[4] a_116499_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4246 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4247 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4248 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4249 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4250 x6[4].x3.ckb x6[4].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4251 cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4252 vdref x4[3].x3.ckb x4[3].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4253 vdref x10[8].x2.swp x10[8].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4254 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4255 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4256 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4257 vsref swn_in[3] a_114064_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4258 vsref cdac_sw_1_1.x2.swp cdac_sw_1_1.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4259 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4260 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4261 vsref cdac_sw_4_1.x1.x8.A cdac_sw_4_1.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4262 cdac_sw_8_0.x1.x3.Y cf[3] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4263 cdac_sw_2_0.x2.swn cdac_sw_2_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4264 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4265 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4266 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4267 cdac_sw_4_1.x2.swn cdac_sw_4_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4268 vsref cdac_sw_2_1.x1.x11.A cdac_sw_2_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4269 x10[8].x3.ckb x10[8].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4270 vsref x6[4].x1.x10.A x6[4].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4271 x4[3].x3.ck x4[3].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4272 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4273 vsref cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4274 vsref cdac_sw_8_0.x2.swp cdac_sw_8_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4275 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4276 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4277 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4278 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4279 vdref x8[7].x1.x11.A x8[7].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4280 cdac_sw_8_1.x2.swn cdac_sw_8_1.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4281 cdac_sw_16_0.x2.swp cdac_sw_16_0.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4282 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4283 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4284 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4285 vdref x8[7].x1.x9.A x8[7].x1.x4.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4286 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4287 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4288 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4289 vsref x2[0].x1.x11.A x2[0].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4290 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4291 vdref x2[0].x2.swp x2[0].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4292 vsref x6[4].x3.ckb x6[4].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4293 a_104404_n15188# cdac_sw_16_0.x3.ck x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4294 cdac_sw_16_0.x2.swp cdac_sw_16_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4295 vsref x10[8].x1.x10.A x10[8].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4296 cdac_sw_2_1.x3.ck cdac_sw_2_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4297 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4298 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4299 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4300 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4301 vdref x8[6].x1.x10.A x8[6].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4302 x8[6].x3.ckb x8[6].x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4303 x10b_cap_array_0.SW[4] cdac_sw_4_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4304 vsref x6[5].x1.x11.A x6[5].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4305 x3[1].x2.swp x3[1].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4306 x8[7].dac_out x8[7].x3.ck a_111430_n6256# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4307 cdac_sw_2_1.x1.x7.A cdac_sw_2_1.x1.x5.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4308 cdac_sw_4_1.x3.ckb cdac_sw_4_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4309 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4310 vdref cdac_sw_4_0.x3.ckb cdac_sw_4_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4311 cdac_sw_1_1.x1.x11.A cdac_sw_1_1.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4312 x2[0].x1.x10.A x2[0].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4313 a_119719_n16821# cdac_sw_4_0.x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4314 vsref x10[8].x1.x9.A a_109227_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4315 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4316 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4317 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4318 vdref x10[8].x1.x5.A x10[8].x1.x7.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4319 x10b_cap_array_0.SW[0] cdac_sw_16_0.x3.ckb a_103526_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4320 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4321 vdref cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4322 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4323 x6[5].x2.swp x6[5].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4324 cdac_sw_8_1.x3.ckb cdac_sw_8_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4325 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4326 vdref cdac_sw_1_2.x1.x11.A cdac_sw_1_2.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4327 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4328 x10b_cap_array_0.SW[1] x2[0].x3.ckb a_106746_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4329 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4330 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4331 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4332 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4333 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4334 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4335 vsref x8[6].x3.ckb x8[6].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4336 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4337 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4338 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4339 a_107624_n15188# x2[0].x3.ck x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4340 x4[3].dac_out x4[3].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4341 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4342 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4343 vdref x10[8].x1.x10.A x10[8].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4344 x10b_cap_array_0.SW[7] cdac_sw_2_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4345 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4346 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4347 x4[3].x2.swp x4[3].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4348 a_114064_n15188# cdac_sw_8_0.x3.ck x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4349 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4350 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4351 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4352 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4353 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4354 x3[1].x2.swn x3[1].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4355 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4356 vsref x4[2].x1.x9.A a_128547_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4357 x4[3].dac_out x4[3].x3.ck a_124310_n8164# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4358 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4359 vsref cdac_sw_2_0.x2.swp cdac_sw_2_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4360 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4361 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4362 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4363 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4364 vsref cdac_sw_2_1.x3.ckb cdac_sw_2_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4365 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4366 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4367 vdref cdac_sw_8_0.x1.x8.A cdac_sw_8_0.x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4368 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4369 vdref x6[4].x1.x11.A x6[4].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4370 a_130750_n10708# swp_in[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4371 vsref cdac_sw_4_0.x1.x9.A cdac_sw_4_0.x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4372 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4373 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4374 vsref x6[4].x1.x8.A x6[4].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4375 vsref x4[2].x1.x6.A x4[2].x1.x8.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4376 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4377 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4378 vdref x3[1].x2.swp x3[1].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4379 vsref cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4380 cdac_sw_16_0.x1.x8.A cdac_sw_16_0.x1.x6.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4381 cdac_sw_4_1.x2.swp cdac_sw_4_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4382 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4383 a_103619_n15957# cdac_sw_16_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4384 vdref x2[0].x1.x8.A x2[0].x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4385 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4386 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4387 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4388 cdac_sw_16_0.x3.ck cdac_sw_16_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4389 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4390 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4391 x10[8].x1.x4.A cf[8] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4392 vdref cdac_sw_8_0.x1.x9.A cdac_sw_8_0.x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4393 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4394 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4395 vsref x4[3].x2.swp x4[3].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4396 cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4397 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4398 x8[6].x1.x11.A x8[6].x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4399 vdref x4[3].x1.x10.A x4[3].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4400 vcm cdac_sw_4_0.x2.swn x10b_cap_array_0.SW[5] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4401 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4402 x6[4].x2.swp x6[4].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4403 vsref x10[8].x1.x8.A x10[8].x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4404 cdac_sw_1_1.x3.ck cdac_sw_1_1.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4405 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4406 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4407 vsref x10[8].x1.x7.A x10[8].x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4408 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4409 vcm cdac_sw_8_1.x2.swn x10b_cap_array_0.SW[2] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4410 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4411 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4412 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4413 a_134987_n5199# cf[0] x3[0].x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4414 vdref cdac_sw_4_1.x3.ckb cdac_sw_4_1.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4415 cdac_sw_2_1.x3.ckb cdac_sw_2_1.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4416 vdref cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4417 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4418 vdref swp_in[4] a_121968_n7755# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4419 cdac_sw_8_0.x3.ck cdac_sw_8_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4420 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4421 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4422 x6[5].x2.swn x6[5].x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4423 x10[8].x2.swp x10[8].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4424 cdac_sw_4_0.x2.swn cdac_sw_4_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4425 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4426 vcm x6[5].x2.swp x6[5].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4427 a_124310_n8164# swp_in[3] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4428 vcn x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4429 cdac_sw_1_1.x2.swp cdac_sw_1_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4430 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4431 x2[0].x3.ckb x2[0].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4432 vcp x3[1].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4433 vsref cdac_sw_8_1.x3.ckb cdac_sw_8_1.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4434 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4435 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4436 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4437 x4[3].x3.ck x4[3].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4438 x4[2].x1.x4.A cf[2] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4439 vsref x4[3].x3.ckb x4[3].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4440 vsref swn_in[2] a_110844_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4441 x2[0].x1.x8.A x2[0].x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4442 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4443 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4444 vcm cdac_sw_16_0.x2.swn x10b_cap_array_0.SW[0] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4445 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4446 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4447 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4448 a_133970_n10708# swp_in[0] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4449 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4450 vdref swp_in[1] a_131628_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4451 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4452 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4453 x8[6].x2.swp x8[6].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4454 vsref cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4455 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4456 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4457 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4458 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4459 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4460 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4461 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4462 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4463 x4[3].x3.ck x4[3].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4464 vsref cdac_sw_1_1.x1.x8.A cdac_sw_1_1.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4465 vdref cdac_sw_4_0.x3.ckb cdac_sw_4_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4466 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4467 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4468 x8[6].x2.swn x8[6].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4469 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4470 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4471 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4472 vsref x8[7].x1.x9.A a_112447_n5199# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4473 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4474 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4475 cdac_sw_4_1.x3.ck cdac_sw_4_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4476 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4477 vdref x4[3].x1.x4.A x4[3].x1.x6.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4478 x3[0].dac_out x3[0].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4479 vdref cdac_sw_8_0.x1.x10.A cdac_sw_8_0.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4480 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4481 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4482 vsref x8[6].x1.x10.A x8[6].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4483 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4484 x6[5].x3.ck x6[5].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4485 a_106746_n15179# swn_in[1] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4486 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4487 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4488 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4489 vdref x8[6].x2.swp x8[6].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4490 vdref cdac_sw_8_0.x3.ckb cdac_sw_8_0.x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4491 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4492 vsref x3[0].x2.swp x3[0].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4493 vdref cdac_sw_4_0.x2.swp cdac_sw_4_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4494 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4495 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4496 x2[0].x1.x11.A x2[0].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4497 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4498 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4499 x6[4].x1.x11.A x6[4].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4500 vcm cdac_sw_4_1.x2.swn x10b_cap_array_0.SW[4] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4501 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4502 vdref swp_in[0] a_134848_n14187# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4503 cdac_sw_2_0.x3.ck cdac_sw_2_0.x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4504 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4505 vsref x6[4].x1.x11.A x6[4].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4506 vdref cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4507 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4508 vdref x6[5].x3.ckb x6[5].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4509 cdac_sw_1_1.x3.ckb cdac_sw_1_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4510 cdac_sw_8_1.x2.swp cdac_sw_8_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4511 vsref x6[4].x2.swp x6[4].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4512 x4[3].x3.ck x4[3].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4513 a_132599_n16821# cdac_sw_1_0.x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4514 x10[8].x2.swn x10[8].x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4515 cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4516 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4517 cdac_sw_1_0.x2.swn cdac_sw_1_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4518 vcm x3[1].x2.swp x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4519 vdref cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4520 vsref x6[4].x1.x3.Y a_122107_n4335# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4521 x10[8].x1.x11.A x10[8].x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4522 x4[3].x1.x10.A x4[3].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4523 a_103526_n15179# swn_in[0] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4524 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4525 vcn x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4526 vsref x10[8].x1.x10.A x10[8].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4527 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4528 x8[7].x3.ck x8[7].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4529 vsref x2[0].x3.ckb x2[0].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4530 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4531 vdref x10[8].x2.swp x10[8].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4532 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4533 cdac_sw_16_0.x3.ck cdac_sw_16_0.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4534 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4535 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4536 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4537 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4538 x8[7].x1.x4.A cf[7] vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4539 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4540 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4541 vcm x2[0].x2.swn x10b_cap_array_0.SW[1] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4542 vdref swp_in[6] a_115528_n6683# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4543 x10b_cap_array_0.SW[3] cdac_sw_8_0.x3.ckb a_113186_n15179# vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4544 cdac_sw_2_0.x1.x4.A cf[7] a_126159_n15957# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4545 cdac_sw_8_1.x1.x9.A cdac_sw_8_1.x1.x7.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4546 vsref x8[7].x1.x7.A x8[7].x1.x9.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4547 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4548 vsref swn_in[9] a_133384_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4549 vcm x3[0].x2.swp x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4550 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4551 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4552 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4553 x6[5].x2.swp x6[5].x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4554 cdac_sw_16_0.x1.x9.A cdac_sw_16_0.x1.x7.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4555 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4556 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4557 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4558 x10b_cap_array_0.SW[2] cdac_sw_8_1.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4559 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4560 vsref cdac_sw_2_0.x1.x8.A cdac_sw_2_0.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4561 vdref x2[0].x1.x9.A x2[0].x1.x11.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4562 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4563 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4564 cdac_sw_2_1.x1.x10.A cdac_sw_2_1.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4565 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4566 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4567 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4568 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4569 a_109227_n5199# cf[8] x10[8].x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4570 x4[2].dac_out x4[2].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4571 a_131628_n14187# x3[1].x3.ckb x3[1].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4572 vsref cdac_sw_1_0.x1.x11.A cdac_sw_1_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4573 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4574 vsref x4[3].x1.x10.A x4[3].x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4575 vsref cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4576 cdac_sw_1_1.x2.swp cdac_sw_1_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4577 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4578 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4579 a_114064_n15188# cdac_sw_8_0.x3.ck x10b_cap_array_0.SW[3] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4580 cdac_sw_1_1.x2.swn cdac_sw_1_1.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4581 vdref cdac_sw_4_0.x1.x8.A cdac_sw_4_0.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4582 vsref x6[5].x1.x11.A x6[5].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4583 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4584 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4585 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4586 vsref cf[2] x4[2].x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4587 x10b_cap_array_0.SW[0] cdac_sw_16_0.x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4588 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4589 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4590 vdref cdac_sw_4_1.x2.swp cdac_sw_4_1.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4591 cdac_sw_2_1.x2.swp cdac_sw_2_1.x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4592 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4593 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4594 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4595 a_121968_n7755# x6[4].x3.ckb x6[4].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4596 cdac_sw_8_0.x2.swn cdac_sw_8_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4597 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4598 vsref cdac_sw_8_1.x1.x11.A cdac_sw_8_1.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4599 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4600 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4601 x2[0].x1.x3.Y cf[1] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4602 vcn x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4603 vsref x6[4].x1.x9.A x6[4].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4604 vdref x6[5].x1.x10.A x6[5].x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4605 x3[1].x3.ckb x3[1].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4606 x8[6].x2.swp x8[6].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4607 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4608 x2[0].x2.swp x2[0].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4609 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4610 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4611 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4612 vsref cdac_sw_16_0.x3.ckb cdac_sw_16_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4613 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4614 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4615 a_121090_n6892# swp_in[4] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4616 cdac_sw_4_1.x1.x10.A cdac_sw_4_1.x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4617 a_129379_n16821# cdac_sw_1_1.x1.x3.Y vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4618 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4619 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4620 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4621 vsref cdac_sw_1_2.x2.swp cdac_sw_1_2.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4622 x4[3].x3.ck x4[3].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4623 a_128547_n5199# cf[2] x4[2].x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4624 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4625 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4626 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4627 x6[5].x3.ckb x6[5].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4628 cdac_sw_8_1.x1.x4.A cdac_sw_8_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4629 cdac_sw_4_0.x3.ckb cdac_sw_4_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4630 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4631 x6[4].x2.swp x6[4].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4632 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4633 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4634 x3[1].dac_out x3[1].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4635 cdac_sw_4_0.x1.x8.A cdac_sw_4_0.x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4636 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4637 vsref cdac_sw_2_1.x1.x8.A cdac_sw_2_1.x1.x10.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4638 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4639 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4640 vdref cdac_sw_4_0.x2.swp cdac_sw_4_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4641 cdac_sw_4_1.x1.x7.A cdac_sw_4_1.x1.x5.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4642 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4643 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4644 vcn x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4645 a_127530_n8164# swp_in[2] vsref vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4646 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4647 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4648 a_128408_n9899# x4[2].x3.ckb x4[2].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4649 vsref cdac_sw_4_0.x2.swp cdac_sw_4_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4650 vsref x8[6].x1.x9.A x8[6].x1.x11.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4651 x10[8].x2.swp x10[8].x1.x11.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4652 x4[3].x3.ckb x4[3].x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4653 a_123724_n15188# cdac_sw_2_1.x3.ck x10b_cap_array_0.SW[6] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4654 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4655 vsref x4[3].x1.x4.A x4[3].x1.x6.A vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4656 vdref cdac_sw_8_0.x1.x11.A cdac_sw_8_0.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4657 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4658 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4659 cdac_sw_16_0.x1.x10.A cdac_sw_16_0.x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4660 vsref x4[3].x2.swp x4[3].x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4661 x10b_cap_array_0.SW[1] x2[0].x2.swp vcm vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4662 vsref swn_in[2] a_110844_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4663 x3[0].dac_out x3[0].x3.ck a_133970_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4664 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4665 x6[5].x3.ck x6[5].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4666 x3[1].dac_out x3[1].x3.ck a_130750_n10708# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4667 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4668 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4669 vsref cdac_sw_1_0.x3.ckb cdac_sw_1_0.x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4670 vdref cdac_sw_8_0.x2.swp cdac_sw_8_0.x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4671 vsref cdac_sw_16_0.x2.swp cdac_sw_16_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4672 cdac_sw_8_1.x2.swp cdac_sw_8_1.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4673 cdac_sw_1_0.x2.swn cdac_sw_1_0.x2.swp vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4674 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4675 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4676 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4677 cdac_sw_1_1.x3.ck cdac_sw_1_1.x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4678 vdref x3[0].x1.x11.A x3[0].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4679 vdref x10[8].x1.x11.A x10[8].x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4680 vcp x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4681 vdref cdac_sw_1_2.x1.x7.A cdac_sw_1_2.x1.x9.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4682 a_113186_n15179# swn_in[3] vdref vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4683 a_134848_n14187# x3[0].x3.ckb x3[0].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4684 vsref cdac_sw_2_0.x1.x10.A cdac_sw_2_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4685 cdac_sw_2_0.x2.swp cdac_sw_2_0.x1.x11.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4686 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4687 a_133384_n15188# cdac_sw_1_0.x3.ck x10b_cap_array_0.SW[9] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4688 cdac_sw_2_0.x2.swn cdac_sw_2_0.x2.swp vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4689 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4690 a_113279_n15957# cdac_sw_8_0.x1.x9.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4691 cdac_sw_2_1.x3.ckb cdac_sw_2_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4692 vdref cdac_sw_4_1.x1.x8.A cdac_sw_4_1.x1.x10.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4693 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4694 vsref cdac_sw_4_0.x1.x10.A cdac_sw_4_0.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4695 vsref x6[5].x3.ckb x6[5].x3.ck vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4696 vdref x3[0].x1.x3.Y x3[0].x1.x5.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4697 vdref x4[3].x3.ckb x4[3].x3.ck vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4698 x4[3].x3.ck x4[3].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4699 cdac_sw_4_0.x1.x11.A cdac_sw_4_0.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4700 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4701 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4702 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4703 vsref cf[7] x8[7].x1.x3.Y vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4704 vdref x10[8].x2.swp x10[8].x2.swn vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4705 x8[6].x1.x10.A x8[6].x1.x8.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4706 vcm cdac_sw_1_1.x2.swn x10b_cap_array_0.SW[8] vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4707 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4708 vcn x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4709 vdref cdac_sw_4_1.x1.x11.A cdac_sw_4_1.x2.swp vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4710 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4711 vdref x10[8].x1.x6.A x10[8].x1.x8.A vdref sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4712 x4[3].x1.x10.A x4[3].x1.x8.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4713 vsref x2[0].x1.x11.A x2[0].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4714 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4715 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4716 x2[0].x1.x5.A x2[0].x1.x8.A a_106839_n16821# vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4717 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4718 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4719 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4720 vsref x8[6].x1.x11.A x8[6].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4721 a_125188_n9899# x4[3].x3.ckb x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4722 cdac_sw_1_0.x3.ckb cdac_sw_1_0.x1.x10.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4723 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4724 vsref swn_in[0] a_104404_n15188# vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4725 cdac_sw_2_1.x1.x4.A cdac_sw_2_1.x1.x9.A vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4726 x8[7].x3.ck x8[7].x3.ckb vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4727 vdref cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x3.ckb vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4728 x6[5].x3.ck x6[5].x3.ckb vdref vdref sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4729 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4730 a_112447_n5199# cf[7] x8[7].x1.x4.A vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4731 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4732 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4733 vcp x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4734 vsref cdac_sw_1_1.x1.x10.A cdac_sw_1_1.x3.ckb vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4735 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4736 vsref x6[4].x1.x11.A x6[4].x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4737 cdac_sw_4_1.x1.x8.A cdac_sw_4_1.x1.x6.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4738 vsref cdac_sw_1_0.x2.swp cdac_sw_1_0.x2.swn vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4739 vcn x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4740 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4741 x8[6].dac_out x8[6].x2.swn vcm vsref sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4742 a_125188_n9899# x4[3].x3.ckb x4[3].dac_out vdref sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4743 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4744 vcn x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4745 vcp x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4746 vcp x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4747 vsref cdac_sw_2_0.x1.x11.A cdac_sw_2_0.x2.swp vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4748 cdac_sw_8_1.x3.ckb cdac_sw_8_1.x1.x10.A vsref vsref sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4749 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4750 vcp x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4751 vcp cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 vcn vsref 0.398342p
C1 vcp vsref 0.398342p
C2 swn_in[9] vsref 17.743198f
C3 swn_in[8] vsref 17.8092f
C4 swp_in[0] vsref 43.1834f
C5 swp_in[1] vsref 43.117302f
C6 swn_in[7] vsref 19.517801f
C7 swn_in[6] vsref 19.583801f
C8 swn_in[5] vsref 22.952099f
C9 swn_in[4] vsref 23.0181f
C10 swn_in[3] vsref 28.8857f
C11 swn_in[2] vsref 28.951698f
C12 swp_in[2] vsref 28.951698f
C13 swp_in[3] vsref 28.8857f
C14 swp_in[4] vsref 23.0181f
C15 swp_in[5] vsref 22.952099f
C16 swp_in[6] vsref 19.583801f
C17 swp_in[7] vsref 19.517801f
C18 swn_in[1] vsref 43.117302f
C19 swn_in[0] vsref 43.1834f
C20 swp_in[8] vsref 17.8092f
C21 swp_in[9] vsref 17.743198f
C22 vcm vsref 0.236244p
C23 cf[0] vsref 29.3552f
C24 cf[1] vsref 29.3552f
C25 cf[2] vsref 24.063599f
C26 cf[3] vsref 24.063599f
C27 cf[4] vsref 24.0349f
C28 cf[5] vsref 24.0349f
C29 cf[6] vsref 24.0061f
C30 cf[7] vsref 24.0061f
C31 cf[8] vsref 23.9917f
C32 cf[9] vsref 23.9917f
C33 vdref vsref 0.857427p
C34 m1_118408_n27032# vsref 0.091357f $ **FLOATING
C35 m1_120148_5902# vsref 0.091357f $ **FLOATING
C36 cdac_sw_1_0.x1.x11.A vsref 2.51762f $ **FLOATING
C37 cdac_sw_1_0.x1.x7.A vsref 0.615623f $ **FLOATING
C38 cdac_sw_1_0.x1.x5.A vsref 0.736451f $ **FLOATING
C39 cdac_sw_1_0.x1.x3.Y vsref 0.60393f $ **FLOATING
C40 cdac_sw_1_1.x1.x11.A vsref 2.51762f $ **FLOATING
C41 cdac_sw_1_1.x1.x7.A vsref 0.615623f $ **FLOATING
C42 cdac_sw_1_1.x1.x5.A vsref 0.736451f $ **FLOATING
C43 cdac_sw_1_1.x1.x3.Y vsref 0.60393f $ **FLOATING
C44 cdac_sw_2_0.x1.x11.A vsref 2.51762f $ **FLOATING
C45 cdac_sw_2_0.x1.x7.A vsref 0.615623f $ **FLOATING
C46 cdac_sw_2_0.x1.x5.A vsref 0.736451f $ **FLOATING
C47 cdac_sw_2_0.x1.x3.Y vsref 0.60393f $ **FLOATING
C48 cdac_sw_2_1.x1.x11.A vsref 2.51762f $ **FLOATING
C49 cdac_sw_2_1.x1.x7.A vsref 0.615623f $ **FLOATING
C50 cdac_sw_2_1.x1.x5.A vsref 0.736451f $ **FLOATING
C51 cdac_sw_2_1.x1.x3.Y vsref 0.60393f $ **FLOATING
C52 cdac_sw_4_0.x1.x11.A vsref 2.51762f $ **FLOATING
C53 cdac_sw_4_0.x1.x7.A vsref 0.615623f $ **FLOATING
C54 cdac_sw_4_0.x1.x5.A vsref 0.736451f $ **FLOATING
C55 cdac_sw_4_0.x1.x3.Y vsref 0.60393f $ **FLOATING
C56 cdac_sw_4_1.x1.x11.A vsref 2.51762f $ **FLOATING
C57 cdac_sw_4_1.x1.x7.A vsref 0.615623f $ **FLOATING
C58 cdac_sw_4_1.x1.x5.A vsref 0.736451f $ **FLOATING
C59 cdac_sw_4_1.x1.x3.Y vsref 0.60393f $ **FLOATING
C60 cdac_sw_8_0.x1.x11.A vsref 2.51762f $ **FLOATING
C61 cdac_sw_8_0.x1.x7.A vsref 0.615623f $ **FLOATING
C62 cdac_sw_8_0.x1.x5.A vsref 0.736451f $ **FLOATING
C63 cdac_sw_8_0.x1.x3.Y vsref 0.60393f $ **FLOATING
C64 cdac_sw_8_1.x1.x11.A vsref 2.51762f $ **FLOATING
C65 cdac_sw_8_1.x1.x7.A vsref 0.615623f $ **FLOATING
C66 cdac_sw_8_1.x1.x5.A vsref 0.736451f $ **FLOATING
C67 cdac_sw_8_1.x1.x3.Y vsref 0.60393f $ **FLOATING
C68 x2[0].x1.x11.A vsref 2.51762f $ **FLOATING
C69 x2[0].x1.x7.A vsref 0.615623f $ **FLOATING
C70 x2[0].x1.x5.A vsref 0.736451f $ **FLOATING
C71 x2[0].x1.x3.Y vsref 0.60393f $ **FLOATING
C72 cdac_sw_16_0.x1.x11.A vsref 2.51762f $ **FLOATING
C73 cdac_sw_16_0.x1.x7.A vsref 0.615623f $ **FLOATING
C74 cdac_sw_16_0.x1.x5.A vsref 0.736451f $ **FLOATING
C75 cdac_sw_16_0.x1.x3.Y vsref 0.60393f $ **FLOATING
C76 cdac_sw_1_0.x1.x10.A vsref 2.51762f $ **FLOATING
C77 cdac_sw_1_0.x1.x8.A vsref 2.14748f $ **FLOATING
C78 cdac_sw_1_0.x1.x6.A vsref 0.615623f $ **FLOATING
C79 cdac_sw_1_0.x1.x4.A vsref 0.736451f $ **FLOATING
C80 cdac_sw_1_0.x1.x9.A vsref 2.26866f $ **FLOATING
C81 cdac_sw_1_1.x1.x10.A vsref 2.51762f $ **FLOATING
C82 cdac_sw_1_1.x1.x8.A vsref 2.14748f $ **FLOATING
C83 cdac_sw_1_1.x1.x6.A vsref 0.615623f $ **FLOATING
C84 cdac_sw_1_1.x1.x4.A vsref 0.736451f $ **FLOATING
C85 cdac_sw_1_1.x1.x9.A vsref 2.26866f $ **FLOATING
C86 cdac_sw_2_0.x1.x10.A vsref 2.51762f $ **FLOATING
C87 cdac_sw_2_0.x1.x8.A vsref 2.14748f $ **FLOATING
C88 cdac_sw_2_0.x1.x6.A vsref 0.615623f $ **FLOATING
C89 cdac_sw_2_0.x1.x4.A vsref 0.736451f $ **FLOATING
C90 cdac_sw_2_0.x1.x9.A vsref 2.26866f $ **FLOATING
C91 cdac_sw_2_1.x1.x10.A vsref 2.51762f $ **FLOATING
C92 cdac_sw_2_1.x1.x8.A vsref 2.14748f $ **FLOATING
C93 cdac_sw_2_1.x1.x6.A vsref 0.615623f $ **FLOATING
C94 cdac_sw_2_1.x1.x4.A vsref 0.736451f $ **FLOATING
C95 cdac_sw_2_1.x1.x9.A vsref 2.26866f $ **FLOATING
C96 cdac_sw_4_0.x1.x10.A vsref 2.51762f $ **FLOATING
C97 cdac_sw_4_0.x1.x8.A vsref 2.14748f $ **FLOATING
C98 cdac_sw_4_0.x1.x6.A vsref 0.615623f $ **FLOATING
C99 cdac_sw_4_0.x1.x4.A vsref 0.736451f $ **FLOATING
C100 cdac_sw_4_0.x1.x9.A vsref 2.26866f $ **FLOATING
C101 cdac_sw_4_1.x1.x10.A vsref 2.51762f $ **FLOATING
C102 cdac_sw_4_1.x1.x8.A vsref 2.14748f $ **FLOATING
C103 cdac_sw_4_1.x1.x6.A vsref 0.615623f $ **FLOATING
C104 cdac_sw_4_1.x1.x4.A vsref 0.736451f $ **FLOATING
C105 cdac_sw_4_1.x1.x9.A vsref 2.26866f $ **FLOATING
C106 cdac_sw_8_0.x1.x10.A vsref 2.51762f $ **FLOATING
C107 cdac_sw_8_0.x1.x8.A vsref 2.14748f $ **FLOATING
C108 cdac_sw_8_0.x1.x6.A vsref 0.615623f $ **FLOATING
C109 cdac_sw_8_0.x1.x4.A vsref 0.736451f $ **FLOATING
C110 cdac_sw_8_0.x1.x9.A vsref 2.26866f $ **FLOATING
C111 cdac_sw_8_1.x1.x10.A vsref 2.51762f $ **FLOATING
C112 cdac_sw_8_1.x1.x8.A vsref 2.14748f $ **FLOATING
C113 cdac_sw_8_1.x1.x6.A vsref 0.615623f $ **FLOATING
C114 cdac_sw_8_1.x1.x4.A vsref 0.736451f $ **FLOATING
C115 cdac_sw_8_1.x1.x9.A vsref 2.26866f $ **FLOATING
C116 x2[0].x1.x10.A vsref 2.51762f $ **FLOATING
C117 x2[0].x1.x8.A vsref 2.14748f $ **FLOATING
C118 x2[0].x1.x6.A vsref 0.615623f $ **FLOATING
C119 x2[0].x1.x4.A vsref 0.736451f $ **FLOATING
C120 x2[0].x1.x9.A vsref 2.26866f $ **FLOATING
C121 cdac_sw_16_0.x1.x10.A vsref 2.51762f $ **FLOATING
C122 cdac_sw_16_0.x1.x8.A vsref 2.14748f $ **FLOATING
C123 cdac_sw_16_0.x1.x6.A vsref 0.615623f $ **FLOATING
C124 cdac_sw_16_0.x1.x4.A vsref 0.736451f $ **FLOATING
C125 cdac_sw_16_0.x1.x9.A vsref 2.26866f $ **FLOATING
C126 cdac_sw_1_0.x2.swn vsref 2.78825f $ **FLOATING
C127 cdac_sw_1_0.x2.swp vsref 4.63322f $ **FLOATING
C128 a_133384_n15188# vsref 0.295532f $ **FLOATING
C129 cdac_sw_1_0.x3.ck vsref 3.14422f $ **FLOATING
C130 x10b_cap_array_0.SW[9] vsref 0.499508p $ **FLOATING
C131 cdac_sw_1_0.x3.ckb vsref 5.12291f $ **FLOATING
C132 a_132506_n15179# vsref 0.588398f $ **FLOATING
C133 cdac_sw_1_1.x2.swn vsref 2.78825f $ **FLOATING
C134 cdac_sw_1_1.x2.swp vsref 4.63322f $ **FLOATING
C135 a_130164_n15188# vsref 0.295532f $ **FLOATING
C136 cdac_sw_1_1.x3.ck vsref 3.14422f $ **FLOATING
C137 x10b_cap_array_0.SW[8] vsref 0.259038p $ **FLOATING
C138 cdac_sw_1_1.x3.ckb vsref 5.12291f $ **FLOATING
C139 a_129286_n15179# vsref 0.588398f $ **FLOATING
C140 cdac_sw_2_0.x2.swn vsref 3.409f $ **FLOATING
C141 a_134848_n14187# vsref 16.1733f $ **FLOATING
C142 a_133970_n10708# vsref 8.6969f $ **FLOATING
C143 x3[0].dac_out vsref 52.5439f $ **FLOATING
C144 a_131628_n14187# vsref 16.1733f $ **FLOATING
C145 a_130750_n10708# vsref 8.6969f $ **FLOATING
C146 cdac_sw_2_0.x2.swp vsref 5.35635f $ **FLOATING
C147 a_126944_n15188# vsref 0.940559f $ **FLOATING
C148 cdac_sw_2_0.x3.ck vsref 3.76497f $ **FLOATING
C149 x10b_cap_array_0.SW[7] vsref 0.140663p $ **FLOATING
C150 cdac_sw_2_0.x3.ckb vsref 5.84648f $ **FLOATING
C151 a_126066_n15179# vsref 1.90105f $ **FLOATING
C152 cdac_sw_2_1.x2.swn vsref 3.409f $ **FLOATING
C153 cdac_sw_2_1.x2.swp vsref 5.35635f $ **FLOATING
C154 a_123724_n15188# vsref 0.940559f $ **FLOATING
C155 cdac_sw_2_1.x3.ck vsref 3.76497f $ **FLOATING
C156 x10b_cap_array_0.SW[6] vsref 80.502f $ **FLOATING
C157 cdac_sw_2_1.x3.ckb vsref 5.84648f $ **FLOATING
C158 a_122846_n15179# vsref 1.90105f $ **FLOATING
C159 cdac_sw_4_0.x2.swn vsref 4.65051f $ **FLOATING
C160 cdac_sw_4_0.x2.swp vsref 6.80262f $ **FLOATING
C161 a_120504_n15188# vsref 2.0817f $ **FLOATING
C162 cdac_sw_4_0.x3.ck vsref 5.00691f $ **FLOATING
C163 x10b_cap_array_0.SW[5] vsref 58.667103f $ **FLOATING
C164 cdac_sw_4_0.x3.ckb vsref 7.29232f $ **FLOATING
C165 a_119626_n15179# vsref 3.93995f $ **FLOATING
C166 cdac_sw_4_1.x2.swn vsref 4.65051f $ **FLOATING
C167 cdac_sw_4_1.x2.swp vsref 6.80262f $ **FLOATING
C168 a_117284_n15188# vsref 2.0817f $ **FLOATING
C169 cdac_sw_4_1.x3.ck vsref 5.00691f $ **FLOATING
C170 x10b_cap_array_0.SW[4] vsref 45.7835f $ **FLOATING
C171 cdac_sw_4_1.x3.ckb vsref 7.29232f $ **FLOATING
C172 a_116406_n15179# vsref 3.93995f $ **FLOATING
C173 cdac_sw_8_0.x2.swn vsref 7.13352f $ **FLOATING
C174 cdac_sw_8_0.x2.swp vsref 9.69516f $ **FLOATING
C175 a_114064_n15188# vsref 4.28676f $ **FLOATING
C176 cdac_sw_8_0.x3.ck vsref 7.49036f $ **FLOATING
C177 x10b_cap_array_0.SW[3] vsref 44.920498f $ **FLOATING
C178 cdac_sw_8_0.x3.ckb vsref 10.1849f $ **FLOATING
C179 a_113186_n15179# vsref 8.01774f $ **FLOATING
C180 cdac_sw_8_1.x2.swn vsref 7.13352f $ **FLOATING
C181 cdac_sw_8_1.x2.swp vsref 9.69516f $ **FLOATING
C182 a_110844_n15188# vsref 4.28676f $ **FLOATING
C183 cdac_sw_8_1.x3.ck vsref 7.49036f $ **FLOATING
C184 x10b_cap_array_0.SW[2] vsref 40.3181f $ **FLOATING
C185 cdac_sw_8_1.x3.ckb vsref 10.1849f $ **FLOATING
C186 a_109966_n15179# vsref 8.01774f $ **FLOATING
C187 x3[1].dac_out vsref 54.380604f $ **FLOATING
C188 x2[0].x2.swn vsref 12.0995f $ **FLOATING
C189 a_128408_n9899# vsref 8.01774f $ **FLOATING
C190 a_127530_n8164# vsref 4.28676f $ **FLOATING
C191 x4[2].dac_out vsref 40.3181f $ **FLOATING
C192 a_125188_n9899# vsref 8.01774f $ **FLOATING
C193 a_124310_n8164# vsref 4.28676f $ **FLOATING
C194 x4[3].dac_out vsref 44.920498f $ **FLOATING
C195 a_121968_n7755# vsref 3.93995f $ **FLOATING
C196 a_121090_n6892# vsref 2.0817f $ **FLOATING
C197 x6[4].dac_out vsref 45.7835f $ **FLOATING
C198 a_118748_n7755# vsref 3.93995f $ **FLOATING
C199 a_117870_n6892# vsref 2.0817f $ **FLOATING
C200 x6[5].dac_out vsref 58.667103f $ **FLOATING
C201 a_115528_n6683# vsref 1.90105f $ **FLOATING
C202 a_114650_n6256# vsref 0.940559f $ **FLOATING
C203 x8[6].dac_out vsref 80.502f $ **FLOATING
C204 a_112308_n6683# vsref 1.90105f $ **FLOATING
C205 a_111430_n6256# vsref 0.940559f $ **FLOATING
C206 x2[0].x2.swp vsref 15.4802f $ **FLOATING
C207 a_107624_n15188# vsref 8.6969f $ **FLOATING
C208 x2[0].x3.ck vsref 12.4572f $ **FLOATING
C209 x10b_cap_array_0.SW[1] vsref 54.380604f $ **FLOATING
C210 x2[0].x3.ckb vsref 15.9699f $ **FLOATING
C211 a_106746_n15179# vsref 16.1733f $ **FLOATING
C212 cdac_sw_16_0.x2.swn vsref 12.0995f $ **FLOATING
C213 cdac_sw_16_0.x2.swp vsref 15.4802f $ **FLOATING
C214 a_104404_n15188# vsref 8.6969f $ **FLOATING
C215 cdac_sw_16_0.x3.ck vsref 12.4572f $ **FLOATING
C216 x10b_cap_array_0.SW[0] vsref 52.5439f $ **FLOATING
C217 cdac_sw_16_0.x3.ckb vsref 15.9699f $ **FLOATING
C218 a_103526_n15179# vsref 16.1733f $ **FLOATING
C219 x8[7].dac_out vsref 0.140663p $ **FLOATING
C220 a_109088_n6147# vsref 0.588398f $ **FLOATING
C221 a_108210_n5938# vsref 0.295532f $ **FLOATING
C222 x10[8].dac_out vsref 0.259038p $ **FLOATING
C223 a_105868_n6147# vsref 0.588398f $ **FLOATING
C224 a_104990_n5938# vsref 0.295532f $ **FLOATING
C225 cdac_sw_1_2.dac_out vsref 0.499508p $ **FLOATING
C226 x3[0].x1.x4.A vsref 0.736451f $ **FLOATING
C227 x3[0].x3.ck vsref 12.4572f $ **FLOATING
C228 x3[0].x1.x6.A vsref 0.615623f $ **FLOATING
C229 x3[0].x1.x10.A vsref 2.51762f $ **FLOATING
C230 x3[0].x3.ckb vsref 15.9699f $ **FLOATING
C231 x3[1].x1.x4.A vsref 0.736451f $ **FLOATING
C232 x3[1].x3.ck vsref 12.4572f $ **FLOATING
C233 x3[1].x1.x6.A vsref 0.615623f $ **FLOATING
C234 x3[1].x1.x10.A vsref 2.51762f $ **FLOATING
C235 x3[1].x3.ckb vsref 15.9699f $ **FLOATING
C236 x4[2].x1.x4.A vsref 0.736451f $ **FLOATING
C237 x4[2].x3.ck vsref 7.49036f $ **FLOATING
C238 x4[2].x1.x6.A vsref 0.615623f $ **FLOATING
C239 x4[2].x1.x10.A vsref 2.51762f $ **FLOATING
C240 x4[2].x3.ckb vsref 10.1849f $ **FLOATING
C241 x4[3].x1.x4.A vsref 0.736451f $ **FLOATING
C242 x4[3].x3.ck vsref 7.49036f $ **FLOATING
C243 x4[3].x1.x6.A vsref 0.615623f $ **FLOATING
C244 x4[3].x1.x10.A vsref 2.51762f $ **FLOATING
C245 x4[3].x3.ckb vsref 10.1849f $ **FLOATING
C246 x6[4].x1.x4.A vsref 0.736451f $ **FLOATING
C247 x6[4].x3.ck vsref 5.00691f $ **FLOATING
C248 x6[4].x1.x6.A vsref 0.615623f $ **FLOATING
C249 x6[4].x1.x10.A vsref 2.51762f $ **FLOATING
C250 x6[4].x3.ckb vsref 7.29232f $ **FLOATING
C251 x6[5].x1.x4.A vsref 0.736451f $ **FLOATING
C252 x6[5].x3.ck vsref 5.00691f $ **FLOATING
C253 x6[5].x1.x6.A vsref 0.615623f $ **FLOATING
C254 x6[5].x1.x10.A vsref 2.51762f $ **FLOATING
C255 x6[5].x3.ckb vsref 7.29232f $ **FLOATING
C256 x8[6].x1.x4.A vsref 0.736451f $ **FLOATING
C257 x8[6].x3.ck vsref 3.76497f $ **FLOATING
C258 x8[6].x1.x6.A vsref 0.615623f $ **FLOATING
C259 x8[6].x1.x10.A vsref 2.51762f $ **FLOATING
C260 x8[6].x3.ckb vsref 5.84648f $ **FLOATING
C261 x8[7].x1.x4.A vsref 0.736451f $ **FLOATING
C262 x8[7].x3.ck vsref 3.76497f $ **FLOATING
C263 x8[7].x1.x6.A vsref 0.615623f $ **FLOATING
C264 x8[7].x1.x10.A vsref 2.51762f $ **FLOATING
C265 x8[7].x3.ckb vsref 5.84648f $ **FLOATING
C266 x10[8].x1.x4.A vsref 0.736451f $ **FLOATING
C267 x10[8].x3.ck vsref 3.14422f $ **FLOATING
C268 x10[8].x1.x6.A vsref 0.615623f $ **FLOATING
C269 x10[8].x1.x10.A vsref 2.51762f $ **FLOATING
C270 x10[8].x3.ckb vsref 5.12291f $ **FLOATING
C271 cdac_sw_1_2.x1.x4.A vsref 0.736451f $ **FLOATING
C272 cdac_sw_1_2.x3.ck vsref 3.14422f $ **FLOATING
C273 cdac_sw_1_2.x1.x6.A vsref 0.615623f $ **FLOATING
C274 cdac_sw_1_2.x1.x10.A vsref 2.51762f $ **FLOATING
C275 cdac_sw_1_2.x3.ckb vsref 5.12291f $ **FLOATING
C276 x3[0].x2.swn vsref 12.0995f $ **FLOATING
C277 x3[1].x2.swn vsref 12.0995f $ **FLOATING
C278 x4[2].x2.swn vsref 7.13352f $ **FLOATING
C279 x4[3].x2.swn vsref 7.13352f $ **FLOATING
C280 x6[4].x2.swn vsref 4.65051f $ **FLOATING
C281 x6[5].x2.swn vsref 4.65051f $ **FLOATING
C282 x8[6].x2.swn vsref 3.409f $ **FLOATING
C283 x8[7].x2.swn vsref 3.409f $ **FLOATING
C284 x10[8].x2.swn vsref 2.78825f $ **FLOATING
C285 cdac_sw_1_2.x2.swn vsref 2.78825f $ **FLOATING
C286 x3[0].x1.x3.Y vsref 0.60393f $ **FLOATING
C287 x3[0].x1.x8.A vsref 2.14748f $ **FLOATING
C288 x3[0].x1.x5.A vsref 0.736451f $ **FLOATING
C289 x3[0].x1.x7.A vsref 0.615623f $ **FLOATING
C290 x3[0].x1.x9.A vsref 2.26866f $ **FLOATING
C291 x3[0].x1.x11.A vsref 2.51762f $ **FLOATING
C292 x3[0].x2.swp vsref 15.4802f $ **FLOATING
C293 x3[1].x1.x3.Y vsref 0.60393f $ **FLOATING
C294 x3[1].x1.x8.A vsref 2.14748f $ **FLOATING
C295 x3[1].x1.x5.A vsref 0.736451f $ **FLOATING
C296 x3[1].x1.x7.A vsref 0.615623f $ **FLOATING
C297 x3[1].x1.x9.A vsref 2.26866f $ **FLOATING
C298 x3[1].x1.x11.A vsref 2.51762f $ **FLOATING
C299 x3[1].x2.swp vsref 15.4802f $ **FLOATING
C300 x4[2].x1.x3.Y vsref 0.60393f $ **FLOATING
C301 x4[2].x1.x8.A vsref 2.14748f $ **FLOATING
C302 x4[2].x1.x5.A vsref 0.736451f $ **FLOATING
C303 x4[2].x1.x7.A vsref 0.615623f $ **FLOATING
C304 x4[2].x1.x9.A vsref 2.26866f $ **FLOATING
C305 x4[2].x1.x11.A vsref 2.51762f $ **FLOATING
C306 x4[2].x2.swp vsref 9.69516f $ **FLOATING
C307 x4[3].x1.x3.Y vsref 0.60393f $ **FLOATING
C308 x4[3].x1.x8.A vsref 2.14748f $ **FLOATING
C309 x4[3].x1.x5.A vsref 0.736451f $ **FLOATING
C310 x4[3].x1.x7.A vsref 0.615623f $ **FLOATING
C311 x4[3].x1.x9.A vsref 2.26866f $ **FLOATING
C312 x4[3].x1.x11.A vsref 2.51762f $ **FLOATING
C313 x4[3].x2.swp vsref 9.69516f $ **FLOATING
C314 x6[4].x1.x3.Y vsref 0.60393f $ **FLOATING
C315 x6[4].x1.x8.A vsref 2.14748f $ **FLOATING
C316 x6[4].x1.x5.A vsref 0.736451f $ **FLOATING
C317 x6[4].x1.x7.A vsref 0.615623f $ **FLOATING
C318 x6[4].x1.x9.A vsref 2.26866f $ **FLOATING
C319 x6[4].x1.x11.A vsref 2.51762f $ **FLOATING
C320 x6[4].x2.swp vsref 6.80262f $ **FLOATING
C321 x6[5].x1.x3.Y vsref 0.60393f $ **FLOATING
C322 x6[5].x1.x8.A vsref 2.14748f $ **FLOATING
C323 x6[5].x1.x5.A vsref 0.736451f $ **FLOATING
C324 x6[5].x1.x7.A vsref 0.615623f $ **FLOATING
C325 x6[5].x1.x9.A vsref 2.26866f $ **FLOATING
C326 x6[5].x1.x11.A vsref 2.51762f $ **FLOATING
C327 x6[5].x2.swp vsref 6.80262f $ **FLOATING
C328 x8[6].x1.x3.Y vsref 0.60393f $ **FLOATING
C329 x8[6].x1.x8.A vsref 2.14748f $ **FLOATING
C330 x8[6].x1.x5.A vsref 0.736451f $ **FLOATING
C331 x8[6].x1.x7.A vsref 0.615623f $ **FLOATING
C332 x8[6].x1.x9.A vsref 2.26866f $ **FLOATING
C333 x8[6].x1.x11.A vsref 2.51762f $ **FLOATING
C334 x8[6].x2.swp vsref 5.35635f $ **FLOATING
C335 x8[7].x1.x3.Y vsref 0.60393f $ **FLOATING
C336 x8[7].x1.x8.A vsref 2.14748f $ **FLOATING
C337 x8[7].x1.x5.A vsref 0.736451f $ **FLOATING
C338 x8[7].x1.x7.A vsref 0.615623f $ **FLOATING
C339 x8[7].x1.x9.A vsref 2.26866f $ **FLOATING
C340 x8[7].x1.x11.A vsref 2.51762f $ **FLOATING
C341 x8[7].x2.swp vsref 5.35635f $ **FLOATING
C342 x10[8].x1.x3.Y vsref 0.60393f $ **FLOATING
C343 x10[8].x1.x8.A vsref 2.14748f $ **FLOATING
C344 x10[8].x1.x5.A vsref 0.736451f $ **FLOATING
C345 x10[8].x1.x7.A vsref 0.615623f $ **FLOATING
C346 x10[8].x1.x9.A vsref 2.26866f $ **FLOATING
C347 x10[8].x1.x11.A vsref 2.51762f $ **FLOATING
C348 x10[8].x2.swp vsref 4.63322f $ **FLOATING
C349 cdac_sw_1_2.x1.x3.Y vsref 0.60393f $ **FLOATING
C350 cdac_sw_1_2.x1.x8.A vsref 2.14748f $ **FLOATING
C351 cdac_sw_1_2.x1.x5.A vsref 0.736451f $ **FLOATING
C352 cdac_sw_1_2.x1.x7.A vsref 0.615623f $ **FLOATING
C353 cdac_sw_1_2.x1.x9.A vsref 2.26866f $ **FLOATING
C354 cdac_sw_1_2.x1.x11.A vsref 2.51762f $ **FLOATING
C355 cdac_sw_1_2.x2.swp vsref 4.63322f $ **FLOATING
