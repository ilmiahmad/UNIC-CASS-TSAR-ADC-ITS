magic
tech sky130A
magscale 1 2
timestamp 1731085074
<< locali >>
rect -106 1173 9858 1175
rect -106 1139 26 1173
rect 3154 1139 3312 1173
rect 6440 1139 6598 1173
rect 9726 1139 9858 1173
rect -106 1105 9858 1139
rect -106 -427 -36 1105
rect 9788 -427 9858 1105
rect -107 -1577 -37 -863
rect 9787 -1577 9857 -863
rect -107 -1647 9857 -1577
<< viali >>
rect 26 1139 3154 1173
rect 3312 1139 6440 1173
rect 6598 1139 9726 1173
rect 6502 -331 6536 1043
rect -107 -1747 9893 -1647
<< metal1 >>
rect -118 1173 9870 1280
rect -118 1169 26 1173
rect 14 1139 26 1169
rect 3154 1169 3312 1173
rect 3154 1139 3166 1169
rect 14 1133 3166 1139
rect 3300 1139 3312 1169
rect 6440 1139 6598 1173
rect 9726 1169 9870 1173
rect 9726 1139 9738 1169
rect 3300 1133 9738 1139
rect 3366 1037 3376 1097
rect 6376 1037 6386 1097
rect 6434 1043 6604 1133
rect 6434 956 6502 1043
rect -11 -244 90 956
rect 3080 -244 3090 956
rect 3148 -244 3158 956
rect 3308 -244 3318 956
rect 3376 -244 3386 956
rect 6382 -244 6502 956
rect -11 -463 39 -244
rect -71 -563 -61 -463
rect 39 -563 49 -463
rect -11 -1037 39 -563
rect 93 -727 143 -285
rect 6496 -331 6502 -244
rect 6536 956 6604 1043
rect 6536 -244 6656 956
rect 9662 -244 9761 956
rect 6536 -331 6542 -244
rect 6496 -343 6542 -331
rect 6665 -463 6715 -285
rect 9711 -463 9761 -244
rect 6606 -563 6616 -463
rect 6715 -563 6725 -463
rect 9701 -563 9711 -463
rect 9811 -563 9821 -463
rect 83 -827 93 -727
rect 193 -827 203 -727
rect 93 -1005 143 -827
rect 6665 -1005 6715 -563
rect 9711 -1037 9761 -563
rect -11 -1437 89 -1037
rect 3095 -1437 3369 -1037
rect 6365 -1437 6375 -1037
rect 6433 -1437 6443 -1037
rect 6593 -1437 6603 -1037
rect 6661 -1437 6671 -1037
rect 9661 -1437 9761 -1037
rect 3147 -1641 3317 -1437
rect 3365 -1569 3375 -1509
rect 6375 -1569 6385 -1509
rect -119 -1647 9905 -1641
rect -119 -1747 -107 -1647
rect 9893 -1747 9905 -1647
rect -119 -1753 9905 -1747
<< via1 >>
rect 3376 1037 6376 1097
rect 3090 -244 3148 956
rect 3318 -244 3376 956
rect -61 -563 39 -463
rect 6616 -563 6715 -463
rect 9711 -563 9811 -463
rect 93 -827 193 -727
rect 6375 -1437 6433 -1037
rect 6603 -1437 6661 -1037
rect 3375 -1569 6375 -1509
<< metal2 >>
rect -106 1097 6376 1107
rect -106 1037 3376 1097
rect -106 1027 6376 1037
rect 3090 956 3376 966
rect 3148 -244 3318 956
rect 3090 -254 3376 -244
rect -61 -463 6715 -453
rect 39 -563 6616 -463
rect -61 -573 6715 -563
rect 9711 -463 9858 -453
rect 9811 -563 9858 -463
rect 9711 -573 9858 -563
rect -107 -727 193 -717
rect -107 -827 93 -727
rect -107 -837 193 -827
rect 6375 -1037 6661 -1027
rect 6433 -1437 6603 -1037
rect 6375 -1447 6661 -1437
rect -107 -1509 6375 -1499
rect -107 -1569 3375 -1509
rect -107 -1579 6375 -1569
use sky130_fd_pr__pfet_01v8_lvt_NZTZAV  XM1
timestamp 1729870836
transform 1 0 1590 0 1 356
box -1696 -819 1696 819
use sky130_fd_pr__pfet_01v8_lvt_NZTZAV  XM2
timestamp 1729870836
transform 1 0 4876 0 1 356
box -1696 -819 1696 819
use sky130_fd_pr__nfet_01v8_lvt_PHPD3W  XM3
timestamp 1729870836
transform 1 0 1589 0 1 -1237
box -1696 -410 1696 410
use sky130_fd_pr__pfet_01v8_lvt_NZTZAV  XM6
timestamp 1729870836
transform 1 0 8162 0 1 356
box -1696 -819 1696 819
use sky130_fd_pr__nfet_01v8_lvt_PHPD3W  XM7
timestamp 1729870836
transform 1 0 4875 0 1 -1237
box -1696 -410 1696 410
use sky130_fd_pr__nfet_01v8_lvt_PHPD3W  XM8
timestamp 1729870836
transform 1 0 8161 0 1 -1237
box -1696 -410 1696 410
<< labels >>
flabel metal2 -97 1032 -33 1095 0 FreeSans 32 0 0 0 vip
port 1 nsew
flabel metal2 -92 -1572 -28 -1509 0 FreeSans 32 0 0 0 vin
port 3 nsew
flabel viali -92 -1727 -26 -1665 0 FreeSans 32 0 0 0 vss
port 7 nsew
flabel metal2 -87 -815 -22 -739 0 FreeSans 32 0 0 0 in
port 2 nsew
flabel metal2 9783 -550 9848 -474 0 FreeSans 32 0 0 0 out
port 8 nsew
<< end >>
