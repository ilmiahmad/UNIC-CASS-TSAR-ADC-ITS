magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect 776 -1954 810 -1878
rect 776 -2044 810 -2038
rect 1162 -1954 1196 -1878
rect 1162 -2044 1196 -2038
rect 1268 -2078 1302 -1878
rect 1268 -2168 1302 -2162
rect 1654 -2078 1688 -1878
rect 1654 -2168 1688 -2162
<< viali >>
rect 776 -2038 810 -1954
rect 1162 -2038 1196 -1954
rect 1268 -2162 1302 -2078
rect 1654 -2162 1688 -2078
<< metal1 >>
rect 940 -1391 960 -1339
rect 1012 -1391 1032 -1339
rect 870 -1481 876 -1429
rect 928 -1481 934 -1429
rect 870 -1553 934 -1481
rect 870 -1605 876 -1553
rect 928 -1605 934 -1553
rect 870 -1677 934 -1605
rect 870 -1729 876 -1677
rect 928 -1729 934 -1677
rect 1038 -1481 1044 -1429
rect 1096 -1481 1102 -1429
rect 1038 -1553 1102 -1481
rect 1038 -1605 1044 -1553
rect 1096 -1605 1102 -1553
rect 1038 -1638 1102 -1605
rect 1432 -1609 1452 -1557
rect 1504 -1609 1524 -1557
rect 1038 -1677 1426 -1638
rect 1038 -1729 1044 -1677
rect 1096 -1729 1426 -1677
rect 1038 -1738 1426 -1729
rect 1530 -1686 1594 -1638
rect 1530 -1738 1536 -1686
rect 1588 -1738 1594 -1686
rect 940 -1819 960 -1767
rect 1012 -1819 1032 -1767
rect 1432 -1819 1452 -1767
rect 1504 -1819 1524 -1767
rect 870 -1899 876 -1847
rect 928 -1899 1536 -1847
rect 1588 -1899 1594 -1847
rect 740 -1954 1724 -1948
rect 740 -2038 776 -1954
rect 810 -2038 1162 -1954
rect 1196 -2038 1724 -1954
rect 740 -2044 1724 -2038
rect 740 -2078 1724 -2072
rect 740 -2162 1268 -2078
rect 1302 -2162 1654 -2078
rect 1688 -2162 1724 -2078
rect 740 -2168 1724 -2162
rect 740 -2248 876 -2196
rect 928 -2248 1724 -2196
rect 740 -2254 1724 -2248
<< via1 >>
rect 960 -1391 1012 -1339
rect 876 -1481 928 -1429
rect 876 -1605 928 -1553
rect 876 -1729 928 -1677
rect 1044 -1481 1096 -1429
rect 1044 -1605 1096 -1553
rect 1452 -1609 1504 -1557
rect 1044 -1729 1096 -1677
rect 1536 -1738 1588 -1686
rect 960 -1819 1012 -1767
rect 1452 -1819 1504 -1767
rect 876 -1899 928 -1847
rect 1536 -1899 1588 -1847
rect 876 -2248 928 -2196
<< metal2 >>
rect 958 -1339 1014 -1333
rect 958 -1391 960 -1339
rect 1012 -1391 1014 -1339
rect 874 -1429 930 -1423
rect 874 -1481 876 -1429
rect 928 -1481 930 -1429
rect 874 -1553 930 -1481
rect 874 -1605 876 -1553
rect 928 -1605 930 -1553
rect 874 -1677 930 -1605
rect 874 -1729 876 -1677
rect 928 -1729 930 -1677
rect 874 -1847 930 -1729
rect 958 -1767 1014 -1391
rect 1042 -1429 1098 -1423
rect 1042 -1481 1044 -1429
rect 1096 -1481 1098 -1429
rect 1042 -1553 1098 -1481
rect 1042 -1605 1044 -1553
rect 1096 -1605 1098 -1553
rect 1042 -1677 1098 -1605
rect 1042 -1729 1044 -1677
rect 1096 -1729 1098 -1677
rect 1042 -1735 1098 -1729
rect 1450 -1557 1506 -1551
rect 1450 -1609 1452 -1557
rect 1504 -1609 1506 -1557
rect 958 -1819 960 -1767
rect 1012 -1819 1014 -1767
rect 958 -1825 1014 -1819
rect 1450 -1767 1506 -1609
rect 1450 -1819 1452 -1767
rect 1504 -1819 1506 -1767
rect 1450 -1825 1506 -1819
rect 1534 -1686 1590 -1680
rect 1534 -1738 1536 -1686
rect 1588 -1738 1590 -1686
rect 874 -1899 876 -1847
rect 928 -1899 930 -1847
rect 874 -2196 930 -1899
rect 1534 -1847 1590 -1738
rect 1534 -1899 1536 -1847
rect 1588 -1899 1590 -1847
rect 1534 -1905 1590 -1899
rect 874 -2248 876 -2196
rect 928 -2248 930 -2196
rect 874 -2254 930 -2248
use sky130_fd_pr__pfet_01v8_TMYSY6  XM1
timestamp 1730624594
transform 1 0 986 0 1 -1579
box -246 -369 246 369
use sky130_fd_pr__nfet_01v8_SMGLWN  XM2
timestamp 1730624594
transform 1 0 1478 0 1 -1688
box -246 -260 246 260
<< labels >>
flabel metal1 740 -2044 836 -1948 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel via1 960 -1819 1012 -1767 0 FreeSans 320 0 0 0 swp
port 2 nsew
flabel via1 1452 -1819 1504 -1767 0 FreeSans 320 0 0 0 swn
port 3 nsew
flabel metal1 740 -2168 836 -2072 0 FreeSans 320 0 0 0 vssa
port 4 nsew
flabel metal1 740 -2254 798 -2196 0 FreeSans 320 0 0 0 in
port 5 nsew
flabel metal2 1044 -1481 1096 -1429 0 FreeSans 320 0 0 0 out
port 6 nsew
<< end >>
