magic
tech sky130A
magscale 1 2
timestamp 1730796434
<< error_p >>
rect 82658 18621 83058 18789
rect 81517 18238 81541 18493
rect 81545 18210 81569 18465
rect 82918 18389 83058 18621
rect 83226 18749 83626 18789
rect 83226 18621 83586 18749
rect 83587 18708 83626 18749
rect 83226 18389 83366 18621
rect 82105 18269 82157 18321
rect 82099 18263 82163 18269
rect 82105 18257 82111 18263
rect 82151 18257 82157 18263
rect 82182 18259 82185 18317
rect 81020 17780 81032 17832
rect 81048 17770 81060 17822
rect 82658 17789 83058 17957
rect 81537 17678 81589 17701
rect 81509 17650 81617 17673
rect 80470 17491 80492 17599
rect 80498 17519 80520 17571
rect 82658 17568 82826 17789
rect 82918 17557 83058 17789
rect 83226 17789 83626 17957
rect 83226 17557 83366 17789
rect 81600 17418 81611 17470
rect 81628 17390 81639 17498
rect 81401 16475 81412 16583
rect 81429 16503 81440 16555
rect 79674 16184 79814 16416
rect 79414 16016 79814 16184
rect 79982 16184 80122 16416
rect 80214 16184 80382 16405
rect 82520 16402 82542 16454
rect 82548 16374 82570 16482
rect 81423 16300 81531 16323
rect 81451 16272 81503 16295
rect 79982 16016 80382 16184
rect 81980 16151 81992 16203
rect 82008 16141 82020 16193
rect 80855 15656 80858 15714
rect 80883 15710 80889 15716
rect 80929 15710 80935 15716
rect 80877 15704 80941 15710
rect 80883 15652 80935 15704
rect 79674 15352 79814 15584
rect 79414 15224 79453 15265
rect 79454 15224 79814 15352
rect 79414 15184 79814 15224
rect 79982 15352 80122 15584
rect 81471 15508 81495 15763
rect 81499 15480 81523 15735
rect 79982 15184 80382 15352
use cdac_10b  cdac_10b_0
timestamp 1730796434
transform 1 0 -18 0 1 30
box -246 -63 67002 60828
use sh_bsw_diff  sh_bsw_diff_0
timestamp 1730796434
transform 1 0 79399 0 1 14689
box -349 -425 4657 5031
use tdc  tdc_0
timestamp 1730796434
transform 1 0 -31840 0 1 13821
box -4836 -3709 9311 2246
<< end >>
