* PEX produced on Sel 12 Nov 2024 06:38:04  CST using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from phase_detector.ext - technology: sky130A

.subckt phase_detector OUT OUTN INN INP VDD VSS
X0 OUT.t0 OUTN.t3 a_15_691.t1 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_n964_406.t1 INP.t0 VSS.t4 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2 VDD.t10 INN.t0 a_n955_1460.t1 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X3 VDD.t13 sky130_fd_sc_hd__nand2_1_1.A.t3 sky130_fd_sc_hd__nand2_1_0.B.t1 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X4 VDD.t1 sky130_fd_sc_hd__nand2_1_1.A.t4 OUTN.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 sky130_fd_sc_hd__nand2_1_0.B.t0 sky130_fd_sc_hd__nand2_1_1.A.t5 a_n964_406.t0 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X6 OUTN.t2 OUT.t3 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_1302_406.t1 INN.t1 VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X8 a_n955_1460.t0 INP.t1 sky130_fd_sc_hd__nand2_1_0.B.t2 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X9 OUT.t2 sky130_fd_sc_hd__nand2_1_0.B.t3 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 sky130_fd_sc_hd__nand2_1_1.A.t2 sky130_fd_sc_hd__nand2_1_0.B.t4 a_1302_406.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X11 VDD.t5 OUTN.t4 OUT.t1 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 VDD.t6 INP.t2 a_893_1460.t0 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X13 VDD.t3 sky130_fd_sc_hd__nand2_1_0.B.t5 sky130_fd_sc_hd__nand2_1_1.A.t0 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X14 a_893_1460.t1 INN.t2 sky130_fd_sc_hd__nand2_1_1.A.t1 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X15 OUTN.t0 sky130_fd_sc_hd__nand2_1_1.A.t6 a_473_691.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_473_691.t1 OUT.t4 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_15_691.t0 sky130_fd_sc_hd__nand2_1_0.B.t6 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 OUTN.n1 OUTN.t4 230.155
R1 OUTN.n3 OUTN.n0 193.548
R2 OUTN.n1 OUTN.t3 157.856
R3 OUTN.n2 OUTN.n1 152
R4 OUTN.n4 OUTN.t0 135.958
R5 OUTN OUTN.n3 44.0308
R6 OUTN.n0 OUTN.t1 26.5955
R7 OUTN.n0 OUTN.t2 26.5955
R8 OUTN.n3 OUTN.n2 23.8989
R9 OUTN.n5 OUTN 16.5652
R10 OUTN.n4 OUTN 14.2478
R11 OUTN.n5 OUTN 9.03579
R12 OUTN.n5 OUTN.n4 4.57193
R13 OUTN.n2 OUTN 2.10199
R14 OUTN OUTN.n5 1.72748
R15 a_15_691.t0 a_15_691.t1 49.8467
R16 OUT OUT.n1 237.577
R17 OUT.n0 OUT.t3 229.369
R18 OUT.n0 OUT.t4 157.07
R19 OUT.n5 OUT.n0 152
R20 OUT.n3 OUT.t0 131.691
R21 OUT.n1 OUT.t1 26.5955
R22 OUT.n1 OUT.t2 26.5955
R23 OUT.n2 OUT 16.5652
R24 OUT.n5 OUT.n4 10.0773
R25 OUT.n4 OUT.n3 9.3005
R26 OUT.n2 OUT 9.03579
R27 OUT.n3 OUT.n2 8.8386
R28 OUT OUT.n5 5.92643
R29 OUT.n4 OUT 5.41118
R30 OUT.n2 OUT 1.72748
R31 VSS.t0 VSS.n29 3609.23
R32 VSS.n31 VSS 3208.68
R33 VSS.n30 VSS.n2 2306.06
R34 VSS.n38 VSS.n2 2306.06
R35 VSS.n32 VSS.n5 2306.06
R36 VSS.n36 VSS.n5 2306.06
R37 VSS.n23 VSS.n10 2306.06
R38 VSS.n23 VSS.n22 2306.06
R39 VSS.n20 VSS.n11 2306.06
R40 VSS.n28 VSS.n11 2306.06
R41 VSS.t5 VSS 1844.97
R42 VSS.n31 VSS.t1 1532.25
R43 VSS.n37 VSS.t1 1532.25
R44 VSS.n21 VSS.t8 1532.25
R45 VSS.n29 VSS.t8 1532.25
R46 VSS.n9 VSS.n8 1489.09
R47 VSS.n8 VSS.n4 1489.09
R48 VSS.n17 VSS.n16 1489.09
R49 VSS.n16 VSS.n12 1489.09
R50 VSS.n30 VSS.n9 816.971
R51 VSS.n32 VSS.n9 816.971
R52 VSS.n36 VSS.n4 816.971
R53 VSS.n38 VSS.n4 816.971
R54 VSS.n12 VSS.n10 816.971
R55 VSS.n20 VSS.n17 816.971
R56 VSS.n22 VSS.n17 816.971
R57 VSS.n28 VSS.n12 816.971
R58 VSS.t6 VSS.t0 509.793
R59 VSS.t2 VSS.t5 509.793
R60 VSS VSS.t6 424.829
R61 VSS VSS.t2 424.829
R62 VSS.n36 VSS.n35 292.5
R63 VSS.n37 VSS.n36 292.5
R64 VSS.n39 VSS.n38 292.5
R65 VSS.n38 VSS.n37 292.5
R66 VSS.n30 VSS.n1 292.5
R67 VSS.n31 VSS.n30 292.5
R68 VSS.n33 VSS.n32 292.5
R69 VSS.n32 VSS.n31 292.5
R70 VSS.n28 VSS.n27 292.5
R71 VSS.n29 VSS.n28 292.5
R72 VSS.n20 VSS.n19 292.5
R73 VSS.n21 VSS.n20 292.5
R74 VSS.n22 VSS.n15 292.5
R75 VSS.n22 VSS.n21 292.5
R76 VSS.n25 VSS.n10 292.5
R77 VSS.n29 VSS.n10 292.5
R78 VSS.n44 VSS.t3 157.988
R79 VSS.n43 VSS.t7 157.988
R80 VSS.n40 VSS.n1 149.835
R81 VSS.n40 VSS.n39 149.835
R82 VSS.n34 VSS.n33 149.835
R83 VSS.n35 VSS.n34 149.835
R84 VSS.n27 VSS.n13 149.835
R85 VSS.n19 VSS.n13 149.835
R86 VSS.n24 VSS.n15 149.835
R87 VSS.n25 VSS.n24 149.835
R88 VSS.n8 VSS.n7 117.001
R89 VSS.n8 VSS.t1 117.001
R90 VSS.n40 VSS.n2 117.001
R91 VSS.t1 VSS.n2 117.001
R92 VSS.n34 VSS.n5 117.001
R93 VSS.n5 VSS.t1 117.001
R94 VSS.n13 VSS.n11 117.001
R95 VSS.n11 VSS.t8 117.001
R96 VSS.n16 VSS.n14 117.001
R97 VSS.n16 VSS.t8 117.001
R98 VSS.n24 VSS.n23 117.001
R99 VSS.n23 VSS.t8 117.001
R100 VSS.n7 VSS.n6 96.7534
R101 VSS.n7 VSS.n3 96.7534
R102 VSS.n18 VSS.n14 96.7534
R103 VSS.n26 VSS.n14 96.7534
R104 VSS.n0 VSS.t9 84.028
R105 VSS.n41 VSS.t4 84.028
R106 VSS.n6 VSS.n1 53.0829
R107 VSS.n33 VSS.n6 53.0829
R108 VSS.n35 VSS.n3 53.0829
R109 VSS.n39 VSS.n3 53.0829
R110 VSS.n27 VSS.n26 53.0829
R111 VSS.n19 VSS.n18 53.0829
R112 VSS.n18 VSS.n15 53.0829
R113 VSS.n26 VSS.n25 53.0829
R114 VSS.n24 VSS.n0 1.95715
R115 VSS.n41 VSS.n40 1.95715
R116 VSS VSS.n41 1.34199
R117 VSS.n42 VSS.n0 0.932201
R118 VSS.n43 VSS.n42 0.858576
R119 VSS VSS.n44 0.504285
R120 VSS.n42 VSS 0.454108
R121 VSS VSS.n43 0.0578348
R122 VSS.n44 VSS 0.0578348
R123 INP.t1 INP.t2 1458.02
R124 INP INP.t1 721.894
R125 INP INP.t0 397.69
R126 a_n964_406.t0 a_n964_406.t1 168.275
R127 INN.t0 INN.t2 1455.17
R128 INN.t2 INN.t1 1119.58
R129 INN INN.t0 721.894
R130 a_n955_1460.t0 a_n955_1460.t1 169.548
R131 VDD.n58 VDD.n9 2142.35
R132 VDD.n54 VDD.n9 2142.35
R133 VDD.n52 VDD.n4 2142.35
R134 VDD.n60 VDD.n4 2142.35
R135 VDD.n36 VDD.n27 2142.35
R136 VDD.n27 VDD.n17 2142.35
R137 VDD.n24 VDD.n18 2142.35
R138 VDD.n44 VDD.n18 2142.35
R139 VDD.n15 VDD.n14 1644.71
R140 VDD.n14 VDD.n8 1644.71
R141 VDD.n51 VDD.n50 1644.71
R142 VDD.n50 VDD.n6 1644.71
R143 VDD.n30 VDD.n25 1644.71
R144 VDD.n30 VDD.n29 1644.71
R145 VDD.n40 VDD.n39 1644.71
R146 VDD.n40 VDD.n19 1644.71
R147 VDD.n58 VDD.n8 497.647
R148 VDD.n51 VDD.n46 497.647
R149 VDD.n46 VDD.n15 497.647
R150 VDD.n54 VDD.n15 497.647
R151 VDD.n52 VDD.n51 497.647
R152 VDD.n60 VDD.n6 497.647
R153 VDD.n7 VDD.n6 497.647
R154 VDD.n8 VDD.n7 497.647
R155 VDD.n36 VDD.n25 497.647
R156 VDD.n19 VDD.n16 497.647
R157 VDD.n29 VDD.n16 497.647
R158 VDD.n29 VDD.n17 497.647
R159 VDD.n39 VDD.n24 497.647
R160 VDD.n39 VDD.n38 497.647
R161 VDD.n38 VDD.n25 497.647
R162 VDD.n44 VDD.n19 497.647
R163 VDD.n37 VDD.t2 426.493
R164 VDD.n45 VDD.t2 426.493
R165 VDD.n53 VDD.t7 426.493
R166 VDD.n59 VDD.t7 426.493
R167 VDD.t4 VDD 278.228
R168 VDD.n75 VDD.t5 249.363
R169 VDD.n69 VDD.t1 249.363
R170 VDD.n77 VDD.t12 247.394
R171 VDD.n67 VDD.t9 247.394
R172 VDD.n57 VDD.n56 228.518
R173 VDD.n56 VDD.n55 228.518
R174 VDD.n62 VDD.n3 228.518
R175 VDD.n62 VDD.n61 228.518
R176 VDD.n34 VDD.n33 228.518
R177 VDD.n35 VDD.n34 228.518
R178 VDD.n43 VDD.n20 228.518
R179 VDD.n23 VDD.n20 228.518
R180 VDD.n13 VDD.n12 175.435
R181 VDD.n13 VDD.n11 175.435
R182 VDD.n49 VDD.n48 175.435
R183 VDD.n49 VDD.n5 175.435
R184 VDD.n31 VDD.n28 175.435
R185 VDD.n32 VDD.n31 175.435
R186 VDD.n41 VDD.n22 175.435
R187 VDD.n42 VDD.n41 175.435
R188 VDD.t0 VDD.n45 169.316
R189 VDD.n53 VDD 108.912
R190 VDD.n61 VDD.n60 92.5005
R191 VDD.n60 VDD.n59 92.5005
R192 VDD.n10 VDD.n7 92.5005
R193 VDD.n59 VDD.n7 92.5005
R194 VDD.n58 VDD.n57 92.5005
R195 VDD.n59 VDD.n58 92.5005
R196 VDD.n55 VDD.n54 92.5005
R197 VDD.n54 VDD.n53 92.5005
R198 VDD.n47 VDD.n46 92.5005
R199 VDD.n53 VDD.n46 92.5005
R200 VDD.n52 VDD.n3 92.5005
R201 VDD.n53 VDD.n52 92.5005
R202 VDD.n36 VDD.n35 92.5005
R203 VDD.n37 VDD.n36 92.5005
R204 VDD.n33 VDD.n17 92.5005
R205 VDD.n45 VDD.n17 92.5005
R206 VDD.n38 VDD.n26 92.5005
R207 VDD.n38 VDD.n37 92.5005
R208 VDD.n44 VDD.n43 92.5005
R209 VDD.n45 VDD.n44 92.5005
R210 VDD.n21 VDD.n16 92.5005
R211 VDD.n45 VDD.n16 92.5005
R212 VDD.n24 VDD.n23 92.5005
R213 VDD.n37 VDD.n24 92.5005
R214 VDD.n80 VDD.t13 89.8482
R215 VDD.n72 VDD.t3 89.8122
R216 VDD.n63 VDD.t10 84.664
R217 VDD.n2 VDD.t6 84.664
R218 VDD.t8 VDD.t0 76.8791
R219 VDD.t11 VDD.t4 76.8791
R220 VDD VDD.t8 64.066
R221 VDD VDD.t11 64.066
R222 VDD.n57 VDD.n11 53.0829
R223 VDD.n48 VDD.n47 53.0829
R224 VDD.n47 VDD.n12 53.0829
R225 VDD.n55 VDD.n12 53.0829
R226 VDD.n48 VDD.n3 53.0829
R227 VDD.n61 VDD.n5 53.0829
R228 VDD.n10 VDD.n5 53.0829
R229 VDD.n11 VDD.n10 53.0829
R230 VDD.n26 VDD.n22 53.0829
R231 VDD.n28 VDD.n26 53.0829
R232 VDD.n33 VDD.n32 53.0829
R233 VDD.n35 VDD.n28 53.0829
R234 VDD.n43 VDD.n42 53.0829
R235 VDD.n42 VDD.n21 53.0829
R236 VDD.n32 VDD.n21 53.0829
R237 VDD.n23 VDD.n22 53.0829
R238 VDD.n76 VDD.n75 25.977
R239 VDD.n69 VDD.n68 25.977
R240 VDD.n77 VDD.n76 24.4711
R241 VDD.n68 VDD.n67 24.4711
R242 VDD.n50 VDD.n49 16.8187
R243 VDD.n50 VDD.t7 16.8187
R244 VDD.n14 VDD.n13 16.8187
R245 VDD.n14 VDD.t7 16.8187
R246 VDD.n56 VDD.n9 16.8187
R247 VDD.n9 VDD.t7 16.8187
R248 VDD.n62 VDD.n4 16.8187
R249 VDD.t7 VDD.n4 16.8187
R250 VDD.n34 VDD.n27 16.8187
R251 VDD.n27 VDD.t2 16.8187
R252 VDD.n31 VDD.n30 16.8187
R253 VDD.n30 VDD.t2 16.8187
R254 VDD.n41 VDD.n40 16.8187
R255 VDD.n40 VDD.t2 16.8187
R256 VDD.n20 VDD.n18 16.8187
R257 VDD.n18 VDD.t2 16.8187
R258 VDD.n70 VDD.n69 9.3005
R259 VDD.n68 VDD.n65 9.3005
R260 VDD.n67 VDD.n66 9.3005
R261 VDD.n75 VDD.n0 9.3005
R262 VDD.n76 VDD.n74 9.3005
R263 VDD.n78 VDD.n77 9.3005
R264 VDD.n73 VDD.n1 4.51973
R265 VDD.n82 VDD.n81 4.51973
R266 VDD.n80 VDD.n79 4.51973
R267 VDD.n72 VDD.n71 4.51973
R268 VDD.n71 VDD.n64 1.27487
R269 VDD.n20 VDD.n2 1.20034
R270 VDD.n63 VDD.n62 1.20034
R271 VDD VDD.n63 0.795603
R272 VDD.n81 VDD.n73 0.663962
R273 VDD.n64 VDD 0.473438
R274 VDD.n81 VDD.n80 0.445212
R275 VDD.n73 VDD.n72 0.442808
R276 VDD.n64 VDD.n2 0.405139
R277 VDD VDD.n82 0.28826
R278 VDD.n70 VDD.n65 0.120292
R279 VDD.n74 VDD.n0 0.120292
R280 VDD.n79 VDD.n74 0.112479
R281 VDD.n65 VDD.n1 0.108573
R282 VDD.n66 VDD 0.0239375
R283 VDD.n78 VDD 0.0239375
R284 VDD.n71 VDD.n70 0.0122188
R285 VDD.n66 VDD.n1 0.0122188
R286 VDD.n82 VDD.n0 0.00961458
R287 VDD.n79 VDD.n78 0.0083125
R288 sky130_fd_sc_hd__nand2_1_1.A.n3 sky130_fd_sc_hd__nand2_1_1.A.t3 717.817
R289 sky130_fd_sc_hd__nand2_1_1.A.n3 sky130_fd_sc_hd__nand2_1_1.A.t5 381.747
R290 sky130_fd_sc_hd__nand2_1_1.A.n1 sky130_fd_sc_hd__nand2_1_1.A.t4 230.155
R291 sky130_fd_sc_hd__nand2_1_1.A.n1 sky130_fd_sc_hd__nand2_1_1.A.t6 157.856
R292 sky130_fd_sc_hd__nand2_1_1.A.n4 sky130_fd_sc_hd__nand2_1_1.A.n1 152
R293 sky130_fd_sc_hd__nand2_1_1.A.n0 sky130_fd_sc_hd__nand2_1_1.A.t1 99.744
R294 sky130_fd_sc_hd__nand2_1_1.A.n2 sky130_fd_sc_hd__nand2_1_1.A.t0 84.6561
R295 sky130_fd_sc_hd__nand2_1_1.A.n2 sky130_fd_sc_hd__nand2_1_1.A.t2 84.0933
R296 sky130_fd_sc_hd__nand2_1_1.A.n4 sky130_fd_sc_hd__nand2_1_1.A.n0 13.8005
R297 sky130_fd_sc_hd__nand2_1_1.A.n0 sky130_fd_sc_hd__nand2_1_1.A.n3 8.307
R298 sky130_fd_sc_hd__nand2_1_1.A.n0 sky130_fd_sc_hd__nand2_1_1.A.n2 6.23388
R299 sky130_fd_sc_hd__nand2_1_1.A sky130_fd_sc_hd__nand2_1_1.A.n4 2.10199
R300 sky130_fd_sc_hd__nand2_1_0.B.n2 sky130_fd_sc_hd__nand2_1_0.B.t5 717.539
R301 sky130_fd_sc_hd__nand2_1_0.B.n2 sky130_fd_sc_hd__nand2_1_0.B.t4 382.024
R302 sky130_fd_sc_hd__nand2_1_0.B.n1 sky130_fd_sc_hd__nand2_1_0.B.t3 229.369
R303 sky130_fd_sc_hd__nand2_1_0.B.n1 sky130_fd_sc_hd__nand2_1_0.B.t6 157.07
R304 sky130_fd_sc_hd__nand2_1_0.B.n4 sky130_fd_sc_hd__nand2_1_0.B.n1 152
R305 sky130_fd_sc_hd__nand2_1_0.B.n0 sky130_fd_sc_hd__nand2_1_0.B.t2 99.4459
R306 sky130_fd_sc_hd__nand2_1_0.B.n3 sky130_fd_sc_hd__nand2_1_0.B.t0 84.4033
R307 sky130_fd_sc_hd__nand2_1_0.B.n3 sky130_fd_sc_hd__nand2_1_0.B.t1 84.3461
R308 sky130_fd_sc_hd__nand2_1_0.B.n4 sky130_fd_sc_hd__nand2_1_0.B.n0 13.9367
R309 sky130_fd_sc_hd__nand2_1_0.B.n0 sky130_fd_sc_hd__nand2_1_0.B.n2 8.31548
R310 sky130_fd_sc_hd__nand2_1_0.B.n0 sky130_fd_sc_hd__nand2_1_0.B.n3 6.2204
R311 sky130_fd_sc_hd__nand2_1_0.B sky130_fd_sc_hd__nand2_1_0.B.n4 5.92643
R312 a_1302_406.t0 a_1302_406.t1 168.275
R313 a_893_1460.t0 a_893_1460.t1 169.548
R314 a_473_691.t0 a_473_691.t1 49.8467
C0 sky130_fd_sc_hd__nand2_1_0.B INN 0.260361f
C1 VDD OUTN 0.68162f
C2 sky130_fd_sc_hd__nand2_1_1.A OUTN 0.348394f
C3 INP INN 0.316567f
C4 VDD sky130_fd_sc_hd__nand2_1_0.B 2.55121f
C5 sky130_fd_sc_hd__nand2_1_0.B sky130_fd_sc_hd__nand2_1_1.A 1.56027f
C6 OUT VDD 0.336255f
C7 INP VDD 1.07005f
C8 OUT sky130_fd_sc_hd__nand2_1_1.A 0.386287f
C9 INP sky130_fd_sc_hd__nand2_1_1.A 0.26762f
C10 sky130_fd_sc_hd__nand2_1_0.B OUTN 0.295843f
C11 VDD INN 1.49464f
C12 sky130_fd_sc_hd__nand2_1_1.A INN 0.147982f
C13 OUT OUTN 0.34321f
C14 VDD sky130_fd_sc_hd__nand2_1_1.A 2.0435f
C15 OUT sky130_fd_sc_hd__nand2_1_0.B 0.110433f
C16 INP sky130_fd_sc_hd__nand2_1_0.B 0.150243f
C17 OUT VSS 0.693673f
C18 OUTN VSS 0.484651f
C19 INP VSS 1.45184f
C20 INN VSS 1.26224f
C21 VDD VSS 12.108155f
C22 sky130_fd_sc_hd__nand2_1_1.A VSS 1.281186f
C23 sky130_fd_sc_hd__nand2_1_0.B VSS 1.034938f
C24 sky130_fd_sc_hd__nand2_1_0.B.n0 VSS 1.05323f
C25 sky130_fd_sc_hd__nand2_1_0.B.t3 VSS 0.024984f
C26 sky130_fd_sc_hd__nand2_1_0.B.t6 VSS 0.015592f
C27 sky130_fd_sc_hd__nand2_1_0.B.n1 VSS 0.049158f
C28 sky130_fd_sc_hd__nand2_1_0.B.t5 VSS 0.112699f
C29 sky130_fd_sc_hd__nand2_1_0.B.t4 VSS 0.063098f
C30 sky130_fd_sc_hd__nand2_1_0.B.n2 VSS 0.3435f
C31 sky130_fd_sc_hd__nand2_1_0.B.t1 VSS 0.181196f
C32 sky130_fd_sc_hd__nand2_1_0.B.t0 VSS 0.057939f
C33 sky130_fd_sc_hd__nand2_1_0.B.n3 VSS 0.423038f
C34 sky130_fd_sc_hd__nand2_1_0.B.t2 VSS 0.242161f
C35 sky130_fd_sc_hd__nand2_1_0.B.n4 VSS 0.026911f
C36 sky130_fd_sc_hd__nand2_1_1.A.n0 VSS 0.822986f
C37 sky130_fd_sc_hd__nand2_1_1.A.t4 VSS 0.019075f
C38 sky130_fd_sc_hd__nand2_1_1.A.t6 VSS 0.01191f
C39 sky130_fd_sc_hd__nand2_1_1.A.n1 VSS 0.036309f
C40 sky130_fd_sc_hd__nand2_1_1.A.t0 VSS 0.138855f
C41 sky130_fd_sc_hd__nand2_1_1.A.t2 VSS 0.043796f
C42 sky130_fd_sc_hd__nand2_1_1.A.n2 VSS 0.322247f
C43 sky130_fd_sc_hd__nand2_1_1.A.t1 VSS 0.186869f
C44 sky130_fd_sc_hd__nand2_1_1.A.t3 VSS 0.085969f
C45 sky130_fd_sc_hd__nand2_1_1.A.t5 VSS 0.048052f
C46 sky130_fd_sc_hd__nand2_1_1.A.n3 VSS 0.261649f
C47 sky130_fd_sc_hd__nand2_1_1.A.n4 VSS 0.018997f
C48 VDD.t3 VSS 0.035442f
C49 VDD.t6 VSS 0.032436f
C50 VDD.n2 VSS 0.125759f
C51 VDD.t10 VSS 0.032436f
C52 VDD.n3 VSS 0.013105f
C53 VDD.n4 VSS 0.020819f
C54 VDD.n5 VSS 0.013238f
C55 VDD.n6 VSS 0.013238f
C56 VDD.t7 VSS 0.465145f
C57 VDD.n8 VSS 0.013238f
C58 VDD.n9 VSS 0.020819f
C59 VDD.n11 VSS 0.013238f
C60 VDD.n12 VSS 0.013238f
C61 VDD.n13 VSS 0.015778f
C62 VDD.n14 VSS 0.015778f
C63 VDD.n15 VSS 0.013238f
C64 VDD.t2 VSS 0.465145f
C65 VDD.n17 VSS 0.013105f
C66 VDD.n18 VSS 0.020819f
C67 VDD.n19 VSS 0.013238f
C68 VDD.n20 VSS 0.039549f
C69 VDD.n22 VSS 0.013238f
C70 VDD.n23 VSS 0.013105f
C71 VDD.n24 VSS 0.013105f
C72 VDD.n25 VSS 0.013238f
C73 VDD.n27 VSS 0.020819f
C74 VDD.n28 VSS 0.013238f
C75 VDD.n29 VSS 0.013238f
C76 VDD.n30 VSS 0.015778f
C77 VDD.n31 VSS 0.015778f
C78 VDD.n32 VSS 0.013238f
C79 VDD.n33 VSS 0.013105f
C80 VDD.n34 VSS 0.020819f
C81 VDD.n35 VSS 0.013105f
C82 VDD.n36 VSS 0.013105f
C83 VDD.n37 VSS 0.295625f
C84 VDD.n39 VSS 0.013238f
C85 VDD.n40 VSS 0.015778f
C86 VDD.n41 VSS 0.015778f
C87 VDD.n42 VSS 0.013238f
C88 VDD.n43 VSS 0.013105f
C89 VDD.n44 VSS 0.013105f
C90 VDD.n45 VSS 0.336455f
C91 VDD.t0 VSS 0.139027f
C92 VDD.t8 VSS 0.079591f
C93 VDD.t4 VSS 0.196424f
C94 VDD.t11 VSS 0.079591f
C95 VDD.n48 VSS 0.013238f
C96 VDD.n49 VSS 0.015778f
C97 VDD.n50 VSS 0.015778f
C98 VDD.n51 VSS 0.013238f
C99 VDD.n52 VSS 0.013105f
C100 VDD.n53 VSS 0.302344f
C101 VDD.n54 VSS 0.013105f
C102 VDD.n55 VSS 0.013105f
C103 VDD.n56 VSS 0.020819f
C104 VDD.n57 VSS 0.013105f
C105 VDD.n58 VSS 0.013105f
C106 VDD.n59 VSS 0.295625f
C107 VDD.n60 VSS 0.013105f
C108 VDD.n61 VSS 0.013105f
C109 VDD.n62 VSS 0.039549f
C110 VDD.n63 VSS 0.140392f
C111 VDD.n64 VSS 0.053053f
C112 VDD.t9 VSS 0.010727f
C113 VDD.n67 VSS 0.014765f
C114 VDD.t1 VSS 0.010723f
C115 VDD.n69 VSS 0.013793f
C116 VDD.n71 VSS 0.023901f
C117 VDD.n72 VSS 0.072085f
C118 VDD.n73 VSS 0.014179f
C119 VDD.t12 VSS 0.010727f
C120 VDD.t5 VSS 0.010723f
C121 VDD.n75 VSS 0.013793f
C122 VDD.n77 VSS 0.014765f
C123 VDD.t13 VSS 0.035469f
C124 VDD.n80 VSS 0.072861f
C125 VDD.n81 VSS 0.014205f
C126 VDD.n82 VSS 0.010907f
.ends

