magic
tech sky130A
magscale 1 2
timestamp 1730868527
<< metal1 >>
rect 2801 -4034 3281 -3938
rect 2801 -4158 3281 -4062
rect 61 -4244 3281 -4186
<< via1 >>
rect 767 -4034 863 -3944
rect 330 -4158 426 -4068
<< metal2 >>
rect 1543 -946 1599 -937
rect 472 -1074 528 -1065
rect 330 -4068 426 -4062
rect 330 -4368 426 -4158
rect 472 -4328 528 -1130
rect 1543 -2447 1599 -1002
rect 665 -4328 721 -3755
rect 767 -3944 863 -3938
rect 767 -4368 863 -4034
rect 1157 -4328 1213 -3755
rect 2035 -4328 2091 -3755
rect 2527 -4328 2583 -3755
<< via2 >>
rect 749 -874 805 -818
rect 2119 -874 2175 -818
rect 1543 -1002 1599 -946
rect 472 -1130 528 -1074
<< metal3 >>
rect 744 -818 3281 -812
rect 744 -874 749 -818
rect 805 -874 2119 -818
rect 2175 -874 3281 -818
rect 744 -880 3281 -874
rect 1538 -946 3281 -940
rect 1538 -1002 1543 -946
rect 1599 -1002 3281 -946
rect 1538 -1008 3281 -1002
rect 467 -1074 3281 -1068
rect 467 -1130 472 -1074
rect 528 -1130 3281 -1074
rect 467 -1136 3281 -1130
use nooverlap_clk  x1
timestamp 1730868527
transform 1 0 585 0 1 -4673
box -562 -783 2734 401
use tg_sw_8  x2
timestamp 1730624594
transform 1 0 1748 0 1 -1986
box 69 -2258 1053 2538
use dac_sw_8  x3
timestamp 1730624594
transform 1 0 -181 0 1 -1797
box 242 -2361 1998 2349
<< labels >>
flabel metal1 3185 -4034 3281 -3938 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel metal1 3185 -4158 3281 -4062 0 FreeSans 320 0 0 0 vssa
port 5 nsew
flabel metal1 3223 -4244 3281 -4186 0 FreeSans 320 0 0 0 vcm
port 4 nsew
flabel metal3 3213 -1136 3281 -1068 0 FreeSans 320 0 0 0 cki
port 2 nsew
flabel metal3 3213 -1008 3281 -940 0 FreeSans 320 0 0 0 bi
port 3 nsew
flabel metal3 3213 -880 3281 -812 0 FreeSans 320 0 0 0 dac_out
port 6 nsew
<< end >>
