magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect -606 -2116 -572 -2040
rect -606 -2206 -572 -2200
rect -220 -2116 -186 -2040
rect -220 -2206 -186 -2200
rect 166 -2116 200 -2040
rect 166 -2206 200 -2200
rect 272 -2240 306 -2040
rect 272 -2330 306 -2324
rect 658 -2240 692 -2040
rect 658 -2330 692 -2324
rect 1044 -2240 1078 -2040
rect 1044 -2330 1078 -2324
<< viali >>
rect -606 -2200 -572 -2116
rect -220 -2200 -186 -2116
rect 166 -2200 200 -2116
rect 272 -2324 306 -2240
rect 658 -2324 692 -2240
rect 1044 -2324 1078 -2240
<< metal1 >>
rect -442 6487 -422 6539
rect -370 6487 -350 6539
rect -56 6487 -36 6539
rect 16 6487 36 6539
rect -512 6397 -506 6449
rect -454 6397 -448 6449
rect -512 6325 -448 6397
rect -512 6273 -506 6325
rect -454 6273 -448 6325
rect -512 6201 -448 6273
rect -512 6149 -506 6201
rect -454 6149 -448 6201
rect -344 6397 -338 6449
rect -286 6397 -120 6449
rect -68 6397 -62 6449
rect -344 6325 -62 6397
rect -344 6273 -338 6325
rect -286 6273 -120 6325
rect -68 6273 -62 6325
rect -344 6201 -62 6273
rect -344 6149 -338 6201
rect -286 6149 -120 6201
rect -68 6149 -62 6201
rect 42 6397 48 6449
rect 100 6397 106 6449
rect 42 6325 106 6397
rect 42 6273 48 6325
rect 100 6273 106 6325
rect 42 6201 106 6273
rect 42 6149 48 6201
rect 100 6149 106 6201
rect -442 6059 -422 6111
rect -370 6059 -350 6111
rect -56 6059 -36 6111
rect 16 6059 36 6111
rect -442 5951 -422 6003
rect -370 5951 -350 6003
rect -56 5951 -36 6003
rect 16 5951 36 6003
rect -512 5861 -506 5913
rect -454 5861 -448 5913
rect -512 5789 -448 5861
rect -512 5737 -506 5789
rect -454 5737 -448 5789
rect -512 5665 -448 5737
rect -512 5613 -506 5665
rect -454 5613 -448 5665
rect -344 5861 -338 5913
rect -286 5861 -120 5913
rect -68 5861 -62 5913
rect -344 5789 -62 5861
rect -344 5737 -338 5789
rect -286 5737 -120 5789
rect -68 5737 -62 5789
rect -344 5665 -62 5737
rect -344 5613 -338 5665
rect -286 5613 -120 5665
rect -68 5613 -62 5665
rect 42 5861 48 5913
rect 100 5861 106 5913
rect 42 5789 106 5861
rect 42 5737 48 5789
rect 100 5737 106 5789
rect 42 5665 106 5737
rect 42 5613 48 5665
rect 100 5613 106 5665
rect -442 5523 -422 5575
rect -370 5523 -350 5575
rect -56 5523 -36 5575
rect 16 5523 36 5575
rect -442 5415 -422 5467
rect -370 5415 -350 5467
rect -56 5415 -36 5467
rect 16 5415 36 5467
rect -512 5325 -506 5377
rect -454 5325 -448 5377
rect -512 5253 -448 5325
rect -512 5201 -506 5253
rect -454 5201 -448 5253
rect -512 5129 -448 5201
rect -512 5077 -506 5129
rect -454 5077 -448 5129
rect -344 5325 -338 5377
rect -286 5325 -120 5377
rect -68 5325 -62 5377
rect -344 5253 -62 5325
rect -344 5201 -338 5253
rect -286 5201 -120 5253
rect -68 5201 -62 5253
rect -344 5129 -62 5201
rect -344 5077 -338 5129
rect -286 5077 -120 5129
rect -68 5077 -62 5129
rect 42 5325 48 5377
rect 100 5325 106 5377
rect 42 5253 106 5325
rect 42 5201 48 5253
rect 100 5201 106 5253
rect 42 5129 106 5201
rect 42 5077 48 5129
rect 100 5077 106 5129
rect -442 4987 -422 5039
rect -370 4987 -350 5039
rect -56 4987 -36 5039
rect 16 4987 36 5039
rect -442 4879 -422 4931
rect -370 4879 -350 4931
rect -56 4879 -36 4931
rect 16 4879 36 4931
rect -512 4789 -506 4841
rect -454 4789 -448 4841
rect -512 4717 -448 4789
rect -512 4665 -506 4717
rect -454 4665 -448 4717
rect -512 4593 -448 4665
rect -512 4541 -506 4593
rect -454 4541 -448 4593
rect -344 4789 -338 4841
rect -286 4789 -120 4841
rect -68 4789 -62 4841
rect -344 4717 -62 4789
rect -344 4665 -338 4717
rect -286 4665 -120 4717
rect -68 4665 -62 4717
rect -344 4593 -62 4665
rect -344 4541 -338 4593
rect -286 4541 -120 4593
rect -68 4541 -62 4593
rect 42 4789 48 4841
rect 100 4789 106 4841
rect 42 4717 106 4789
rect 42 4665 48 4717
rect 100 4665 106 4717
rect 42 4593 106 4665
rect 42 4541 48 4593
rect 100 4541 106 4593
rect -442 4451 -422 4503
rect -370 4451 -350 4503
rect -56 4451 -36 4503
rect 16 4451 36 4503
rect -442 4343 -422 4395
rect -370 4343 -350 4395
rect -56 4343 -36 4395
rect 16 4343 36 4395
rect -512 4253 -506 4305
rect -454 4253 -448 4305
rect -512 4181 -448 4253
rect -512 4129 -506 4181
rect -454 4129 -448 4181
rect -512 4057 -448 4129
rect -512 4005 -506 4057
rect -454 4005 -448 4057
rect -344 4253 -338 4305
rect -286 4253 -120 4305
rect -68 4253 -62 4305
rect -344 4181 -62 4253
rect -344 4129 -338 4181
rect -286 4129 -120 4181
rect -68 4129 -62 4181
rect -344 4057 -62 4129
rect -344 4005 -338 4057
rect -286 4005 -120 4057
rect -68 4005 -62 4057
rect 42 4253 48 4305
rect 100 4253 106 4305
rect 42 4181 106 4253
rect 42 4129 48 4181
rect 100 4129 106 4181
rect 42 4057 106 4129
rect 42 4005 48 4057
rect 100 4005 106 4057
rect -442 3915 -422 3967
rect -370 3915 -350 3967
rect -56 3915 -36 3967
rect 16 3915 36 3967
rect -442 3807 -422 3859
rect -370 3807 -350 3859
rect -56 3807 -36 3859
rect 16 3807 36 3859
rect -512 3717 -506 3769
rect -454 3717 -448 3769
rect -512 3645 -448 3717
rect -512 3593 -506 3645
rect -454 3593 -448 3645
rect -512 3521 -448 3593
rect -512 3469 -506 3521
rect -454 3469 -448 3521
rect -344 3717 -338 3769
rect -286 3717 -120 3769
rect -68 3717 -62 3769
rect -344 3645 -62 3717
rect -344 3593 -338 3645
rect -286 3593 -120 3645
rect -68 3593 -62 3645
rect -344 3521 -62 3593
rect -344 3469 -338 3521
rect -286 3469 -120 3521
rect -68 3469 -62 3521
rect 42 3717 48 3769
rect 100 3717 106 3769
rect 42 3645 106 3717
rect 42 3593 48 3645
rect 100 3593 106 3645
rect 42 3521 106 3593
rect 42 3469 48 3521
rect 100 3469 106 3521
rect -442 3379 -422 3431
rect -370 3379 -350 3431
rect -56 3379 -36 3431
rect 16 3379 36 3431
rect -442 3271 -422 3323
rect -370 3271 -350 3323
rect -56 3271 -36 3323
rect 16 3271 36 3323
rect -512 3181 -506 3233
rect -454 3181 -448 3233
rect -512 3109 -448 3181
rect -512 3057 -506 3109
rect -454 3057 -448 3109
rect -512 2985 -448 3057
rect -512 2933 -506 2985
rect -454 2933 -448 2985
rect -344 3181 -338 3233
rect -286 3181 -120 3233
rect -68 3181 -62 3233
rect -344 3109 -62 3181
rect -344 3057 -338 3109
rect -286 3057 -120 3109
rect -68 3057 -62 3109
rect -344 2985 -62 3057
rect -344 2933 -338 2985
rect -286 2933 -120 2985
rect -68 2933 -62 2985
rect 42 3181 48 3233
rect 100 3181 106 3233
rect 42 3109 106 3181
rect 42 3057 48 3109
rect 100 3057 106 3109
rect 42 2985 106 3057
rect 436 2999 456 3051
rect 508 2999 528 3051
rect 822 2999 842 3051
rect 894 2999 914 3051
rect 42 2933 48 2985
rect 100 2933 106 2985
rect 366 2922 430 2970
rect -442 2843 -422 2895
rect -370 2843 -350 2895
rect -56 2843 -36 2895
rect 16 2843 36 2895
rect 366 2870 372 2922
rect 424 2870 430 2922
rect 534 2922 816 2970
rect 534 2870 540 2922
rect 592 2870 758 2922
rect 810 2870 816 2922
rect 920 2922 984 2970
rect 920 2870 926 2922
rect 978 2870 984 2922
rect 436 2789 456 2841
rect 508 2789 528 2841
rect 822 2789 842 2841
rect 894 2789 914 2841
rect -442 2735 -422 2787
rect -370 2735 -350 2787
rect -56 2735 -36 2787
rect 16 2735 36 2787
rect -512 2645 -506 2697
rect -454 2645 -448 2697
rect -512 2573 -448 2645
rect -512 2521 -506 2573
rect -454 2521 -448 2573
rect -512 2449 -448 2521
rect -512 2397 -506 2449
rect -454 2397 -448 2449
rect -344 2645 -338 2697
rect -286 2645 -120 2697
rect -68 2645 -62 2697
rect -344 2573 -62 2645
rect -344 2521 -338 2573
rect -286 2521 -120 2573
rect -68 2521 -62 2573
rect -344 2449 -62 2521
rect -344 2397 -338 2449
rect -286 2397 -120 2449
rect -68 2397 -62 2449
rect 42 2645 48 2697
rect 100 2652 106 2697
rect 436 2681 456 2733
rect 508 2681 528 2733
rect 822 2681 842 2733
rect 894 2681 914 2733
rect 100 2645 430 2652
rect 42 2604 430 2645
rect 42 2573 372 2604
rect 42 2521 48 2573
rect 100 2552 372 2573
rect 424 2552 430 2604
rect 534 2604 816 2652
rect 534 2552 540 2604
rect 592 2552 758 2604
rect 810 2552 816 2604
rect 920 2604 984 2652
rect 920 2552 926 2604
rect 978 2552 984 2604
rect 100 2521 106 2552
rect 42 2449 106 2521
rect 436 2471 456 2523
rect 508 2471 528 2523
rect 822 2471 842 2523
rect 894 2471 914 2523
rect 42 2397 48 2449
rect 100 2397 106 2449
rect 42 2388 106 2397
rect 437 2363 456 2415
rect 508 2363 529 2415
rect 822 2363 842 2415
rect 894 2363 914 2415
rect -442 2307 -422 2359
rect -370 2307 -350 2359
rect -56 2307 -36 2359
rect 16 2307 36 2359
rect 366 2286 430 2334
rect -442 2199 -422 2251
rect -370 2199 -350 2251
rect -56 2199 -36 2251
rect 16 2199 36 2251
rect 366 2234 372 2286
rect 424 2234 430 2286
rect 534 2286 816 2334
rect 534 2234 540 2286
rect 592 2234 758 2286
rect 810 2234 816 2286
rect 920 2286 984 2334
rect 920 2234 926 2286
rect 978 2234 984 2286
rect -512 2109 -506 2161
rect -454 2109 -448 2161
rect -512 2037 -448 2109
rect -512 1985 -506 2037
rect -454 1985 -448 2037
rect -512 1913 -448 1985
rect -512 1861 -506 1913
rect -454 1861 -448 1913
rect -344 2109 -338 2161
rect -286 2109 -120 2161
rect -68 2109 -62 2161
rect -344 2037 -62 2109
rect -344 1985 -338 2037
rect -286 1985 -120 2037
rect -68 1985 -62 2037
rect -344 1913 -62 1985
rect -344 1861 -338 1913
rect -286 1861 -120 1913
rect -68 1861 -62 1913
rect 42 2109 48 2161
rect 100 2109 106 2161
rect 436 2153 456 2205
rect 508 2153 528 2205
rect 822 2153 842 2205
rect 894 2153 914 2205
rect 42 2037 106 2109
rect 436 2045 456 2097
rect 508 2045 528 2097
rect 821 2045 842 2097
rect 894 2045 913 2097
rect 42 1985 48 2037
rect 100 2017 106 2037
rect 100 1985 430 2017
rect 42 1968 430 1985
rect 42 1917 372 1968
rect 42 1913 106 1917
rect 366 1916 372 1917
rect 424 1916 430 1968
rect 534 1968 816 2016
rect 534 1916 540 1968
rect 592 1916 758 1968
rect 810 1916 816 1968
rect 920 1968 984 2016
rect 920 1916 926 1968
rect 978 1916 984 1968
rect 42 1861 48 1913
rect 100 1861 106 1913
rect 436 1835 456 1887
rect 508 1835 528 1887
rect 822 1835 842 1887
rect 894 1835 914 1887
rect -442 1771 -422 1823
rect -370 1771 -350 1823
rect -56 1771 -36 1823
rect 16 1771 36 1823
rect 436 1727 456 1779
rect 508 1727 528 1779
rect 822 1727 842 1779
rect 894 1727 914 1779
rect -442 1663 -422 1715
rect -370 1663 -350 1715
rect -56 1663 -36 1715
rect 16 1663 36 1715
rect 366 1650 430 1698
rect -512 1573 -506 1625
rect -454 1573 -448 1625
rect -512 1501 -448 1573
rect -512 1449 -506 1501
rect -454 1449 -448 1501
rect -512 1377 -448 1449
rect -512 1325 -506 1377
rect -454 1325 -448 1377
rect -344 1573 -338 1625
rect -286 1573 -120 1625
rect -68 1573 -62 1625
rect -344 1501 -62 1573
rect -344 1449 -338 1501
rect -286 1449 -120 1501
rect -68 1449 -62 1501
rect -344 1377 -62 1449
rect -344 1325 -338 1377
rect -286 1325 -120 1377
rect -68 1325 -62 1377
rect 42 1573 48 1625
rect 100 1573 106 1625
rect 366 1598 372 1650
rect 424 1598 430 1650
rect 534 1650 816 1698
rect 534 1598 540 1650
rect 592 1598 758 1650
rect 810 1598 816 1650
rect 920 1650 984 1698
rect 920 1598 926 1650
rect 978 1598 984 1650
rect 42 1501 106 1573
rect 436 1517 456 1569
rect 508 1517 528 1569
rect 822 1517 842 1569
rect 894 1517 914 1569
rect 42 1449 48 1501
rect 100 1449 106 1501
rect 42 1377 106 1449
rect 436 1409 456 1461
rect 508 1409 528 1461
rect 822 1409 842 1461
rect 894 1409 914 1461
rect 42 1325 48 1377
rect 100 1325 106 1377
rect 366 1332 430 1380
rect -442 1235 -422 1287
rect -370 1235 -350 1287
rect -56 1235 -36 1287
rect 16 1235 36 1287
rect 366 1280 372 1332
rect 424 1280 430 1332
rect 534 1332 816 1380
rect 534 1280 540 1332
rect 592 1280 758 1332
rect 810 1280 816 1332
rect 920 1332 984 1380
rect 920 1280 926 1332
rect 978 1280 984 1332
rect 436 1199 456 1251
rect 508 1199 528 1251
rect 822 1199 842 1251
rect 894 1199 914 1251
rect -442 1127 -422 1179
rect -370 1127 -350 1179
rect -56 1127 -36 1179
rect 16 1127 36 1179
rect 437 1091 456 1143
rect 508 1091 529 1143
rect 822 1091 842 1143
rect 894 1091 914 1143
rect -512 1037 -506 1089
rect -454 1037 -448 1089
rect -512 965 -448 1037
rect -512 913 -506 965
rect -454 913 -448 965
rect -512 841 -448 913
rect -512 789 -506 841
rect -454 789 -448 841
rect -344 1037 -338 1089
rect -286 1037 -120 1089
rect -68 1037 -62 1089
rect -344 965 -62 1037
rect -344 913 -338 965
rect -286 913 -120 965
rect -68 913 -62 965
rect -344 841 -62 913
rect -344 789 -338 841
rect -286 789 -120 841
rect -68 789 -62 841
rect 42 1037 48 1089
rect 100 1062 106 1089
rect 100 1037 430 1062
rect 42 1014 430 1037
rect 42 965 372 1014
rect 42 913 48 965
rect 100 962 372 965
rect 424 962 430 1014
rect 534 1014 816 1062
rect 534 962 540 1014
rect 592 962 758 1014
rect 810 962 816 1014
rect 920 1014 984 1062
rect 920 962 926 1014
rect 978 962 984 1014
rect 100 913 106 962
rect 42 841 106 913
rect 436 881 456 933
rect 508 881 528 933
rect 822 881 842 933
rect 894 881 914 933
rect 42 789 48 841
rect 100 789 106 841
rect 436 773 456 825
rect 508 773 528 825
rect 821 773 842 825
rect 894 773 913 825
rect -442 699 -422 751
rect -370 699 -350 751
rect -56 699 -36 751
rect 16 699 36 751
rect 366 696 430 744
rect 366 644 372 696
rect 424 644 430 696
rect 534 696 816 744
rect 534 644 540 696
rect 592 644 758 696
rect 810 644 816 696
rect 920 696 984 744
rect 920 644 926 696
rect 978 644 984 696
rect -442 591 -422 643
rect -370 591 -350 643
rect -56 591 -36 643
rect 16 591 36 643
rect 436 563 456 615
rect 508 563 528 615
rect 822 563 842 615
rect 894 563 914 615
rect -512 501 -506 553
rect -454 501 -448 553
rect -512 429 -448 501
rect -512 377 -506 429
rect -454 377 -448 429
rect -512 305 -448 377
rect -512 253 -506 305
rect -454 253 -448 305
rect -344 501 -338 553
rect -286 501 -120 553
rect -68 501 -62 553
rect -344 429 -62 501
rect -344 377 -338 429
rect -286 377 -120 429
rect -68 377 -62 429
rect -344 305 -62 377
rect -344 253 -338 305
rect -286 253 -120 305
rect -68 253 -62 305
rect 42 501 48 553
rect 100 501 106 553
rect 42 429 106 501
rect 436 455 456 507
rect 508 455 528 507
rect 822 455 842 507
rect 894 455 914 507
rect 42 377 48 429
rect 100 426 106 429
rect 100 378 430 426
rect 100 377 372 378
rect 42 326 372 377
rect 424 326 430 378
rect 534 378 816 426
rect 534 326 540 378
rect 592 326 758 378
rect 810 326 816 378
rect 920 378 984 426
rect 920 326 926 378
rect 978 326 984 378
rect 42 305 106 326
rect 42 253 48 305
rect 100 253 106 305
rect 436 245 456 297
rect 508 245 528 297
rect 822 245 842 297
rect 894 245 914 297
rect -442 163 -422 215
rect -370 163 -350 215
rect -56 163 -36 215
rect 16 163 36 215
rect 436 137 456 189
rect 508 137 528 189
rect 822 137 842 189
rect 894 137 914 189
rect -442 55 -422 107
rect -370 55 -350 107
rect -56 55 -36 107
rect 16 55 36 107
rect 366 60 430 108
rect -512 -35 -506 17
rect -454 -35 -448 17
rect -512 -107 -448 -35
rect -512 -159 -506 -107
rect -454 -159 -448 -107
rect -512 -231 -448 -159
rect -512 -283 -506 -231
rect -454 -283 -448 -231
rect -344 -35 -338 17
rect -286 -35 -120 17
rect -68 -35 -62 17
rect -344 -107 -62 -35
rect -344 -159 -338 -107
rect -286 -159 -120 -107
rect -68 -159 -62 -107
rect -344 -231 -62 -159
rect -344 -283 -338 -231
rect -286 -283 -120 -231
rect -68 -283 -62 -231
rect 42 -35 48 17
rect 100 -35 106 17
rect 366 8 372 60
rect 424 8 430 60
rect 534 60 816 108
rect 534 8 540 60
rect 592 8 758 60
rect 810 8 816 60
rect 920 60 984 108
rect 920 8 926 60
rect 978 8 984 60
rect 42 -107 106 -35
rect 436 -73 456 -21
rect 508 -73 528 -21
rect 822 -73 842 -21
rect 894 -73 914 -21
rect 42 -159 48 -107
rect 100 -159 106 -107
rect 42 -231 106 -159
rect 437 -181 456 -129
rect 508 -181 529 -129
rect 822 -181 842 -129
rect 894 -181 914 -129
rect 42 -283 48 -231
rect 100 -283 106 -231
rect 366 -258 430 -210
rect 366 -310 372 -258
rect 424 -310 430 -258
rect 534 -258 816 -210
rect 534 -310 540 -258
rect 592 -310 758 -258
rect 810 -310 816 -258
rect 920 -258 984 -210
rect 920 -310 926 -258
rect 978 -310 984 -258
rect -442 -373 -422 -321
rect -370 -373 -350 -321
rect -56 -373 -36 -321
rect 16 -373 36 -321
rect 436 -391 456 -339
rect 508 -391 528 -339
rect 822 -391 842 -339
rect 894 -391 914 -339
rect -442 -481 -422 -429
rect -370 -481 -350 -429
rect -56 -481 -36 -429
rect 16 -481 36 -429
rect 436 -499 456 -447
rect 508 -499 528 -447
rect 821 -499 842 -447
rect 894 -499 913 -447
rect -512 -571 -506 -519
rect -454 -571 -448 -519
rect -512 -643 -448 -571
rect -512 -695 -506 -643
rect -454 -695 -448 -643
rect -512 -767 -448 -695
rect -512 -819 -506 -767
rect -454 -819 -448 -767
rect -344 -571 -338 -519
rect -286 -571 -120 -519
rect -68 -571 -62 -519
rect -344 -643 -62 -571
rect -344 -695 -338 -643
rect -286 -695 -120 -643
rect -68 -695 -62 -643
rect -344 -767 -62 -695
rect -344 -819 -338 -767
rect -286 -819 -120 -767
rect -68 -819 -62 -767
rect 42 -571 48 -519
rect 100 -528 106 -519
rect 100 -571 430 -528
rect 42 -576 430 -571
rect 42 -628 372 -576
rect 424 -628 430 -576
rect 534 -576 816 -528
rect 534 -628 540 -576
rect 592 -628 758 -576
rect 810 -628 816 -576
rect 920 -576 984 -528
rect 920 -628 926 -576
rect 978 -628 984 -576
rect 42 -643 106 -628
rect 42 -695 48 -643
rect 100 -695 106 -643
rect 42 -767 106 -695
rect 436 -709 456 -657
rect 508 -709 528 -657
rect 822 -709 842 -657
rect 894 -709 914 -657
rect 42 -819 48 -767
rect 100 -819 106 -767
rect 436 -817 456 -765
rect 508 -817 528 -765
rect 822 -817 842 -765
rect 894 -817 914 -765
rect -442 -909 -422 -857
rect -370 -909 -350 -857
rect -56 -909 -36 -857
rect 16 -909 36 -857
rect 366 -894 430 -846
rect 366 -946 372 -894
rect 424 -946 430 -894
rect 534 -894 816 -846
rect 534 -946 540 -894
rect 592 -946 758 -894
rect 810 -946 816 -894
rect 920 -894 984 -846
rect 920 -946 926 -894
rect 978 -946 984 -894
rect -442 -1017 -422 -965
rect -370 -1017 -350 -965
rect -56 -1017 -36 -965
rect 16 -1017 36 -965
rect 436 -1027 456 -975
rect 508 -1027 528 -975
rect 822 -1027 842 -975
rect 894 -1027 914 -975
rect -512 -1107 -506 -1055
rect -454 -1107 -448 -1055
rect -512 -1179 -448 -1107
rect -512 -1231 -506 -1179
rect -454 -1231 -448 -1179
rect -512 -1303 -448 -1231
rect -512 -1355 -506 -1303
rect -454 -1355 -448 -1303
rect -344 -1107 -338 -1055
rect -286 -1107 -120 -1055
rect -68 -1107 -62 -1055
rect -344 -1179 -62 -1107
rect -344 -1231 -338 -1179
rect -286 -1231 -120 -1179
rect -68 -1231 -62 -1179
rect -344 -1303 -62 -1231
rect -344 -1355 -338 -1303
rect -286 -1355 -120 -1303
rect -68 -1355 -62 -1303
rect 42 -1107 48 -1055
rect 100 -1107 106 -1055
rect 42 -1164 106 -1107
rect 436 -1135 456 -1083
rect 508 -1135 528 -1083
rect 822 -1135 842 -1083
rect 894 -1135 914 -1083
rect 42 -1179 430 -1164
rect 42 -1231 48 -1179
rect 100 -1212 430 -1179
rect 100 -1231 372 -1212
rect 42 -1264 372 -1231
rect 424 -1264 430 -1212
rect 534 -1212 816 -1164
rect 534 -1264 540 -1212
rect 592 -1264 758 -1212
rect 810 -1264 816 -1212
rect 920 -1212 984 -1164
rect 920 -1264 926 -1212
rect 978 -1264 984 -1212
rect 42 -1303 106 -1264
rect 42 -1355 48 -1303
rect 100 -1355 106 -1303
rect 436 -1345 456 -1293
rect 508 -1345 528 -1293
rect 822 -1345 842 -1293
rect 894 -1345 914 -1293
rect -442 -1445 -422 -1393
rect -370 -1445 -350 -1393
rect -56 -1445 -36 -1393
rect 16 -1445 36 -1393
rect 437 -1453 456 -1401
rect 508 -1453 529 -1401
rect 822 -1453 842 -1401
rect 894 -1453 914 -1401
rect -442 -1553 -422 -1501
rect -370 -1553 -350 -1501
rect -56 -1553 -36 -1501
rect 16 -1553 36 -1501
rect 366 -1530 430 -1482
rect 366 -1582 372 -1530
rect 424 -1582 430 -1530
rect 534 -1530 816 -1482
rect 534 -1582 540 -1530
rect 592 -1582 758 -1530
rect 810 -1582 816 -1530
rect 920 -1530 984 -1482
rect 920 -1582 926 -1530
rect 978 -1582 984 -1530
rect -512 -1643 -506 -1591
rect -454 -1643 -448 -1591
rect -512 -1715 -448 -1643
rect -512 -1767 -506 -1715
rect -454 -1767 -448 -1715
rect -512 -1839 -448 -1767
rect -512 -1891 -506 -1839
rect -454 -1891 -448 -1839
rect -344 -1643 -338 -1591
rect -286 -1643 -120 -1591
rect -68 -1643 -62 -1591
rect -344 -1715 -62 -1643
rect -344 -1767 -338 -1715
rect -286 -1767 -120 -1715
rect -68 -1767 -62 -1715
rect -344 -1839 -62 -1767
rect -344 -1891 -338 -1839
rect -286 -1891 -120 -1839
rect -68 -1891 -62 -1839
rect 42 -1643 48 -1591
rect 100 -1643 106 -1591
rect 42 -1715 106 -1643
rect 436 -1663 456 -1611
rect 508 -1663 528 -1611
rect 822 -1663 842 -1611
rect 894 -1663 914 -1611
rect 42 -1767 48 -1715
rect 100 -1767 106 -1715
rect 42 -1800 106 -1767
rect 436 -1771 456 -1719
rect 508 -1771 528 -1719
rect 821 -1771 842 -1719
rect 894 -1771 913 -1719
rect 42 -1839 430 -1800
rect 42 -1891 48 -1839
rect 100 -1848 430 -1839
rect 100 -1891 372 -1848
rect 42 -1900 372 -1891
rect 424 -1900 430 -1848
rect 534 -1848 816 -1800
rect 534 -1900 540 -1848
rect 592 -1900 758 -1848
rect 810 -1900 816 -1848
rect 920 -1848 984 -1800
rect 920 -1900 926 -1848
rect 978 -1900 984 -1848
rect -442 -1981 -422 -1929
rect -370 -1981 -350 -1929
rect -56 -1981 -36 -1929
rect 16 -1981 36 -1929
rect 436 -1981 456 -1929
rect 508 -1981 528 -1929
rect 822 -1981 842 -1929
rect 894 -1981 914 -1929
rect -428 -2061 -422 -2009
rect -370 -2061 842 -2009
rect 894 -2061 900 -2009
rect -642 -2116 -506 -2110
rect -642 -2200 -606 -2116
rect -572 -2200 -506 -2116
rect -454 -2116 1114 -2110
rect -454 -2200 -220 -2116
rect -186 -2200 166 -2116
rect 200 -2200 1114 -2116
rect -642 -2206 1114 -2200
rect -642 -2240 926 -2234
rect -642 -2324 272 -2240
rect 306 -2324 658 -2240
rect 692 -2324 926 -2240
rect 978 -2240 1114 -2234
rect 978 -2324 1044 -2240
rect 1078 -2324 1114 -2240
rect -642 -2330 1114 -2324
<< via1 >>
rect -422 6487 -370 6539
rect -36 6487 16 6539
rect -506 6397 -454 6449
rect -506 6273 -454 6325
rect -506 6149 -454 6201
rect -338 6397 -286 6449
rect -120 6397 -68 6449
rect -338 6273 -286 6325
rect -120 6273 -68 6325
rect -338 6149 -286 6201
rect -120 6149 -68 6201
rect 48 6397 100 6449
rect 48 6273 100 6325
rect 48 6149 100 6201
rect -422 6059 -370 6111
rect -36 6059 16 6111
rect -422 5951 -370 6003
rect -36 5951 16 6003
rect -506 5861 -454 5913
rect -506 5737 -454 5789
rect -506 5613 -454 5665
rect -338 5861 -286 5913
rect -120 5861 -68 5913
rect -338 5737 -286 5789
rect -120 5737 -68 5789
rect -338 5613 -286 5665
rect -120 5613 -68 5665
rect 48 5861 100 5913
rect 48 5737 100 5789
rect 48 5613 100 5665
rect -422 5523 -370 5575
rect -36 5523 16 5575
rect -422 5415 -370 5467
rect -36 5415 16 5467
rect -506 5325 -454 5377
rect -506 5201 -454 5253
rect -506 5077 -454 5129
rect -338 5325 -286 5377
rect -120 5325 -68 5377
rect -338 5201 -286 5253
rect -120 5201 -68 5253
rect -338 5077 -286 5129
rect -120 5077 -68 5129
rect 48 5325 100 5377
rect 48 5201 100 5253
rect 48 5077 100 5129
rect -422 4987 -370 5039
rect -36 4987 16 5039
rect -422 4879 -370 4931
rect -36 4879 16 4931
rect -506 4789 -454 4841
rect -506 4665 -454 4717
rect -506 4541 -454 4593
rect -338 4789 -286 4841
rect -120 4789 -68 4841
rect -338 4665 -286 4717
rect -120 4665 -68 4717
rect -338 4541 -286 4593
rect -120 4541 -68 4593
rect 48 4789 100 4841
rect 48 4665 100 4717
rect 48 4541 100 4593
rect -422 4451 -370 4503
rect -36 4451 16 4503
rect -422 4343 -370 4395
rect -36 4343 16 4395
rect -506 4253 -454 4305
rect -506 4129 -454 4181
rect -506 4005 -454 4057
rect -338 4253 -286 4305
rect -120 4253 -68 4305
rect -338 4129 -286 4181
rect -120 4129 -68 4181
rect -338 4005 -286 4057
rect -120 4005 -68 4057
rect 48 4253 100 4305
rect 48 4129 100 4181
rect 48 4005 100 4057
rect -422 3915 -370 3967
rect -36 3915 16 3967
rect -422 3807 -370 3859
rect -36 3807 16 3859
rect -506 3717 -454 3769
rect -506 3593 -454 3645
rect -506 3469 -454 3521
rect -338 3717 -286 3769
rect -120 3717 -68 3769
rect -338 3593 -286 3645
rect -120 3593 -68 3645
rect -338 3469 -286 3521
rect -120 3469 -68 3521
rect 48 3717 100 3769
rect 48 3593 100 3645
rect 48 3469 100 3521
rect -422 3379 -370 3431
rect -36 3379 16 3431
rect -422 3271 -370 3323
rect -36 3271 16 3323
rect -506 3181 -454 3233
rect -506 3057 -454 3109
rect -506 2933 -454 2985
rect -338 3181 -286 3233
rect -120 3181 -68 3233
rect -338 3057 -286 3109
rect -120 3057 -68 3109
rect -338 2933 -286 2985
rect -120 2933 -68 2985
rect 48 3181 100 3233
rect 48 3057 100 3109
rect 456 2999 508 3051
rect 842 2999 894 3051
rect 48 2933 100 2985
rect -422 2843 -370 2895
rect -36 2843 16 2895
rect 372 2870 424 2922
rect 540 2870 592 2922
rect 758 2870 810 2922
rect 926 2870 978 2922
rect 456 2789 508 2841
rect 842 2789 894 2841
rect -422 2735 -370 2787
rect -36 2735 16 2787
rect -506 2645 -454 2697
rect -506 2521 -454 2573
rect -506 2397 -454 2449
rect -338 2645 -286 2697
rect -120 2645 -68 2697
rect -338 2521 -286 2573
rect -120 2521 -68 2573
rect -338 2397 -286 2449
rect -120 2397 -68 2449
rect 48 2645 100 2697
rect 456 2681 508 2733
rect 842 2681 894 2733
rect 48 2521 100 2573
rect 372 2552 424 2604
rect 540 2552 592 2604
rect 758 2552 810 2604
rect 926 2552 978 2604
rect 456 2471 508 2523
rect 842 2471 894 2523
rect 48 2397 100 2449
rect 456 2363 508 2415
rect 842 2363 894 2415
rect -422 2307 -370 2359
rect -36 2307 16 2359
rect -422 2199 -370 2251
rect -36 2199 16 2251
rect 372 2234 424 2286
rect 540 2234 592 2286
rect 758 2234 810 2286
rect 926 2234 978 2286
rect -506 2109 -454 2161
rect -506 1985 -454 2037
rect -506 1861 -454 1913
rect -338 2109 -286 2161
rect -120 2109 -68 2161
rect -338 1985 -286 2037
rect -120 1985 -68 2037
rect -338 1861 -286 1913
rect -120 1861 -68 1913
rect 48 2109 100 2161
rect 456 2153 508 2205
rect 842 2153 894 2205
rect 456 2045 508 2097
rect 842 2045 894 2097
rect 48 1985 100 2037
rect 372 1916 424 1968
rect 540 1916 592 1968
rect 758 1916 810 1968
rect 926 1916 978 1968
rect 48 1861 100 1913
rect 456 1835 508 1887
rect 842 1835 894 1887
rect -422 1771 -370 1823
rect -36 1771 16 1823
rect 456 1727 508 1779
rect 842 1727 894 1779
rect -422 1663 -370 1715
rect -36 1663 16 1715
rect -506 1573 -454 1625
rect -506 1449 -454 1501
rect -506 1325 -454 1377
rect -338 1573 -286 1625
rect -120 1573 -68 1625
rect -338 1449 -286 1501
rect -120 1449 -68 1501
rect -338 1325 -286 1377
rect -120 1325 -68 1377
rect 48 1573 100 1625
rect 372 1598 424 1650
rect 540 1598 592 1650
rect 758 1598 810 1650
rect 926 1598 978 1650
rect 456 1517 508 1569
rect 842 1517 894 1569
rect 48 1449 100 1501
rect 456 1409 508 1461
rect 842 1409 894 1461
rect 48 1325 100 1377
rect -422 1235 -370 1287
rect -36 1235 16 1287
rect 372 1280 424 1332
rect 540 1280 592 1332
rect 758 1280 810 1332
rect 926 1280 978 1332
rect 456 1199 508 1251
rect 842 1199 894 1251
rect -422 1127 -370 1179
rect -36 1127 16 1179
rect 456 1091 508 1143
rect 842 1091 894 1143
rect -506 1037 -454 1089
rect -506 913 -454 965
rect -506 789 -454 841
rect -338 1037 -286 1089
rect -120 1037 -68 1089
rect -338 913 -286 965
rect -120 913 -68 965
rect -338 789 -286 841
rect -120 789 -68 841
rect 48 1037 100 1089
rect 48 913 100 965
rect 372 962 424 1014
rect 540 962 592 1014
rect 758 962 810 1014
rect 926 962 978 1014
rect 456 881 508 933
rect 842 881 894 933
rect 48 789 100 841
rect 456 773 508 825
rect 842 773 894 825
rect -422 699 -370 751
rect -36 699 16 751
rect 372 644 424 696
rect 540 644 592 696
rect 758 644 810 696
rect 926 644 978 696
rect -422 591 -370 643
rect -36 591 16 643
rect 456 563 508 615
rect 842 563 894 615
rect -506 501 -454 553
rect -506 377 -454 429
rect -506 253 -454 305
rect -338 501 -286 553
rect -120 501 -68 553
rect -338 377 -286 429
rect -120 377 -68 429
rect -338 253 -286 305
rect -120 253 -68 305
rect 48 501 100 553
rect 456 455 508 507
rect 842 455 894 507
rect 48 377 100 429
rect 372 326 424 378
rect 540 326 592 378
rect 758 326 810 378
rect 926 326 978 378
rect 48 253 100 305
rect 456 245 508 297
rect 842 245 894 297
rect -422 163 -370 215
rect -36 163 16 215
rect 456 137 508 189
rect 842 137 894 189
rect -422 55 -370 107
rect -36 55 16 107
rect -506 -35 -454 17
rect -506 -159 -454 -107
rect -506 -283 -454 -231
rect -338 -35 -286 17
rect -120 -35 -68 17
rect -338 -159 -286 -107
rect -120 -159 -68 -107
rect -338 -283 -286 -231
rect -120 -283 -68 -231
rect 48 -35 100 17
rect 372 8 424 60
rect 540 8 592 60
rect 758 8 810 60
rect 926 8 978 60
rect 456 -73 508 -21
rect 842 -73 894 -21
rect 48 -159 100 -107
rect 456 -181 508 -129
rect 842 -181 894 -129
rect 48 -283 100 -231
rect 372 -310 424 -258
rect 540 -310 592 -258
rect 758 -310 810 -258
rect 926 -310 978 -258
rect -422 -373 -370 -321
rect -36 -373 16 -321
rect 456 -391 508 -339
rect 842 -391 894 -339
rect -422 -481 -370 -429
rect -36 -481 16 -429
rect 456 -499 508 -447
rect 842 -499 894 -447
rect -506 -571 -454 -519
rect -506 -695 -454 -643
rect -506 -819 -454 -767
rect -338 -571 -286 -519
rect -120 -571 -68 -519
rect -338 -695 -286 -643
rect -120 -695 -68 -643
rect -338 -819 -286 -767
rect -120 -819 -68 -767
rect 48 -571 100 -519
rect 372 -628 424 -576
rect 540 -628 592 -576
rect 758 -628 810 -576
rect 926 -628 978 -576
rect 48 -695 100 -643
rect 456 -709 508 -657
rect 842 -709 894 -657
rect 48 -819 100 -767
rect 456 -817 508 -765
rect 842 -817 894 -765
rect -422 -909 -370 -857
rect -36 -909 16 -857
rect 372 -946 424 -894
rect 540 -946 592 -894
rect 758 -946 810 -894
rect 926 -946 978 -894
rect -422 -1017 -370 -965
rect -36 -1017 16 -965
rect 456 -1027 508 -975
rect 842 -1027 894 -975
rect -506 -1107 -454 -1055
rect -506 -1231 -454 -1179
rect -506 -1355 -454 -1303
rect -338 -1107 -286 -1055
rect -120 -1107 -68 -1055
rect -338 -1231 -286 -1179
rect -120 -1231 -68 -1179
rect -338 -1355 -286 -1303
rect -120 -1355 -68 -1303
rect 48 -1107 100 -1055
rect 456 -1135 508 -1083
rect 842 -1135 894 -1083
rect 48 -1231 100 -1179
rect 372 -1264 424 -1212
rect 540 -1264 592 -1212
rect 758 -1264 810 -1212
rect 926 -1264 978 -1212
rect 48 -1355 100 -1303
rect 456 -1345 508 -1293
rect 842 -1345 894 -1293
rect -422 -1445 -370 -1393
rect -36 -1445 16 -1393
rect 456 -1453 508 -1401
rect 842 -1453 894 -1401
rect -422 -1553 -370 -1501
rect -36 -1553 16 -1501
rect 372 -1582 424 -1530
rect 540 -1582 592 -1530
rect 758 -1582 810 -1530
rect 926 -1582 978 -1530
rect -506 -1643 -454 -1591
rect -506 -1767 -454 -1715
rect -506 -1891 -454 -1839
rect -338 -1643 -286 -1591
rect -120 -1643 -68 -1591
rect -338 -1767 -286 -1715
rect -120 -1767 -68 -1715
rect -338 -1891 -286 -1839
rect -120 -1891 -68 -1839
rect 48 -1643 100 -1591
rect 456 -1663 508 -1611
rect 842 -1663 894 -1611
rect 48 -1767 100 -1715
rect 456 -1771 508 -1719
rect 842 -1771 894 -1719
rect 48 -1891 100 -1839
rect 372 -1900 424 -1848
rect 540 -1900 592 -1848
rect 758 -1900 810 -1848
rect 926 -1900 978 -1848
rect -422 -1981 -370 -1929
rect -36 -1981 16 -1929
rect 456 -1981 508 -1929
rect 842 -1981 894 -1929
rect -422 -2061 -370 -2009
rect 842 -2061 894 -2009
rect -506 -2200 -454 -2110
rect 926 -2324 978 -2234
<< metal2 >>
rect -424 6539 -368 6545
rect -424 6487 -422 6539
rect -370 6487 -368 6539
rect -508 6449 -452 6455
rect -508 6397 -506 6449
rect -454 6397 -452 6449
rect -508 6325 -452 6397
rect -508 6273 -506 6325
rect -454 6273 -452 6325
rect -508 6201 -452 6273
rect -508 6149 -506 6201
rect -454 6149 -452 6201
rect -508 5913 -452 6149
rect -508 5861 -506 5913
rect -454 5861 -452 5913
rect -508 5789 -452 5861
rect -508 5737 -506 5789
rect -454 5737 -452 5789
rect -508 5665 -452 5737
rect -508 5613 -506 5665
rect -454 5613 -452 5665
rect -508 5377 -452 5613
rect -508 5325 -506 5377
rect -454 5325 -452 5377
rect -508 5253 -452 5325
rect -508 5201 -506 5253
rect -454 5201 -452 5253
rect -508 5129 -452 5201
rect -508 5077 -506 5129
rect -454 5077 -452 5129
rect -508 4841 -452 5077
rect -508 4789 -506 4841
rect -454 4789 -452 4841
rect -508 4717 -452 4789
rect -508 4665 -506 4717
rect -454 4665 -452 4717
rect -508 4593 -452 4665
rect -508 4541 -506 4593
rect -454 4541 -452 4593
rect -508 4305 -452 4541
rect -508 4253 -506 4305
rect -454 4253 -452 4305
rect -508 4181 -452 4253
rect -508 4129 -506 4181
rect -454 4129 -452 4181
rect -508 4057 -452 4129
rect -508 4005 -506 4057
rect -454 4005 -452 4057
rect -508 3769 -452 4005
rect -508 3717 -506 3769
rect -454 3717 -452 3769
rect -508 3645 -452 3717
rect -508 3593 -506 3645
rect -454 3593 -452 3645
rect -508 3521 -452 3593
rect -508 3469 -506 3521
rect -454 3469 -452 3521
rect -508 3233 -452 3469
rect -508 3181 -506 3233
rect -454 3181 -452 3233
rect -508 3109 -452 3181
rect -508 3057 -506 3109
rect -454 3057 -452 3109
rect -508 2985 -452 3057
rect -508 2933 -506 2985
rect -454 2933 -452 2985
rect -508 2697 -452 2933
rect -508 2645 -506 2697
rect -454 2645 -452 2697
rect -508 2573 -452 2645
rect -508 2521 -506 2573
rect -454 2521 -452 2573
rect -508 2449 -452 2521
rect -508 2397 -506 2449
rect -454 2397 -452 2449
rect -508 2161 -452 2397
rect -508 2109 -506 2161
rect -454 2109 -452 2161
rect -508 2037 -452 2109
rect -508 1985 -506 2037
rect -454 1985 -452 2037
rect -508 1913 -452 1985
rect -508 1861 -506 1913
rect -454 1861 -452 1913
rect -508 1625 -452 1861
rect -508 1573 -506 1625
rect -454 1573 -452 1625
rect -508 1501 -452 1573
rect -508 1449 -506 1501
rect -454 1449 -452 1501
rect -508 1377 -452 1449
rect -508 1325 -506 1377
rect -454 1325 -452 1377
rect -508 1089 -452 1325
rect -508 1037 -506 1089
rect -454 1037 -452 1089
rect -508 965 -452 1037
rect -508 913 -506 965
rect -454 913 -452 965
rect -508 841 -452 913
rect -508 789 -506 841
rect -454 789 -452 841
rect -508 553 -452 789
rect -508 501 -506 553
rect -454 501 -452 553
rect -508 429 -452 501
rect -508 377 -506 429
rect -454 377 -452 429
rect -508 305 -452 377
rect -508 253 -506 305
rect -454 253 -452 305
rect -508 17 -452 253
rect -508 -35 -506 17
rect -454 -35 -452 17
rect -508 -107 -452 -35
rect -508 -159 -506 -107
rect -454 -159 -452 -107
rect -508 -231 -452 -159
rect -508 -283 -506 -231
rect -454 -283 -452 -231
rect -508 -519 -452 -283
rect -508 -571 -506 -519
rect -454 -571 -452 -519
rect -508 -643 -452 -571
rect -508 -695 -506 -643
rect -454 -695 -452 -643
rect -508 -767 -452 -695
rect -508 -819 -506 -767
rect -454 -819 -452 -767
rect -508 -1055 -452 -819
rect -508 -1107 -506 -1055
rect -454 -1107 -452 -1055
rect -508 -1179 -452 -1107
rect -508 -1231 -506 -1179
rect -454 -1231 -452 -1179
rect -508 -1303 -452 -1231
rect -508 -1355 -506 -1303
rect -454 -1355 -452 -1303
rect -508 -1591 -452 -1355
rect -508 -1643 -506 -1591
rect -454 -1643 -452 -1591
rect -508 -1715 -452 -1643
rect -508 -1767 -506 -1715
rect -454 -1767 -452 -1715
rect -508 -1839 -452 -1767
rect -508 -1891 -506 -1839
rect -454 -1891 -452 -1839
rect -508 -2110 -452 -1891
rect -424 6111 -368 6487
rect -38 6539 18 6545
rect -38 6487 -36 6539
rect 16 6487 18 6539
rect -424 6059 -422 6111
rect -370 6059 -368 6111
rect -424 6003 -368 6059
rect -424 5951 -422 6003
rect -370 5951 -368 6003
rect -424 5575 -368 5951
rect -424 5523 -422 5575
rect -370 5523 -368 5575
rect -424 5467 -368 5523
rect -424 5415 -422 5467
rect -370 5415 -368 5467
rect -424 5039 -368 5415
rect -424 4987 -422 5039
rect -370 4987 -368 5039
rect -424 4931 -368 4987
rect -424 4879 -422 4931
rect -370 4879 -368 4931
rect -424 4503 -368 4879
rect -424 4451 -422 4503
rect -370 4451 -368 4503
rect -424 4395 -368 4451
rect -424 4343 -422 4395
rect -370 4343 -368 4395
rect -424 3967 -368 4343
rect -424 3915 -422 3967
rect -370 3915 -368 3967
rect -424 3859 -368 3915
rect -424 3807 -422 3859
rect -370 3807 -368 3859
rect -424 3431 -368 3807
rect -424 3379 -422 3431
rect -370 3379 -368 3431
rect -424 3323 -368 3379
rect -424 3271 -422 3323
rect -370 3271 -368 3323
rect -424 2895 -368 3271
rect -424 2843 -422 2895
rect -370 2843 -368 2895
rect -424 2787 -368 2843
rect -424 2735 -422 2787
rect -370 2735 -368 2787
rect -424 2359 -368 2735
rect -424 2307 -422 2359
rect -370 2307 -368 2359
rect -424 2251 -368 2307
rect -424 2199 -422 2251
rect -370 2199 -368 2251
rect -424 1823 -368 2199
rect -424 1771 -422 1823
rect -370 1771 -368 1823
rect -424 1715 -368 1771
rect -424 1663 -422 1715
rect -370 1663 -368 1715
rect -424 1287 -368 1663
rect -424 1235 -422 1287
rect -370 1235 -368 1287
rect -424 1179 -368 1235
rect -424 1127 -422 1179
rect -370 1127 -368 1179
rect -424 751 -368 1127
rect -424 699 -422 751
rect -370 699 -368 751
rect -424 643 -368 699
rect -424 591 -422 643
rect -370 591 -368 643
rect -424 215 -368 591
rect -424 163 -422 215
rect -370 163 -368 215
rect -424 107 -368 163
rect -424 55 -422 107
rect -370 55 -368 107
rect -424 -321 -368 55
rect -424 -373 -422 -321
rect -370 -373 -368 -321
rect -424 -429 -368 -373
rect -424 -481 -422 -429
rect -370 -481 -368 -429
rect -424 -857 -368 -481
rect -424 -909 -422 -857
rect -370 -909 -368 -857
rect -424 -965 -368 -909
rect -424 -1017 -422 -965
rect -370 -1017 -368 -965
rect -424 -1393 -368 -1017
rect -424 -1445 -422 -1393
rect -370 -1445 -368 -1393
rect -424 -1501 -368 -1445
rect -424 -1553 -422 -1501
rect -370 -1553 -368 -1501
rect -424 -1929 -368 -1553
rect -340 6449 -284 6455
rect -340 6397 -338 6449
rect -286 6397 -284 6449
rect -340 6325 -284 6397
rect -340 6273 -338 6325
rect -286 6273 -284 6325
rect -340 6201 -284 6273
rect -340 6149 -338 6201
rect -286 6149 -284 6201
rect -340 5913 -284 6149
rect -340 5861 -338 5913
rect -286 5861 -284 5913
rect -340 5789 -284 5861
rect -340 5737 -338 5789
rect -286 5737 -284 5789
rect -340 5665 -284 5737
rect -340 5613 -338 5665
rect -286 5613 -284 5665
rect -340 5377 -284 5613
rect -340 5325 -338 5377
rect -286 5325 -284 5377
rect -340 5253 -284 5325
rect -340 5201 -338 5253
rect -286 5201 -284 5253
rect -340 5129 -284 5201
rect -340 5077 -338 5129
rect -286 5077 -284 5129
rect -340 4841 -284 5077
rect -340 4789 -338 4841
rect -286 4789 -284 4841
rect -340 4717 -284 4789
rect -340 4665 -338 4717
rect -286 4665 -284 4717
rect -340 4593 -284 4665
rect -340 4541 -338 4593
rect -286 4541 -284 4593
rect -340 4305 -284 4541
rect -340 4253 -338 4305
rect -286 4253 -284 4305
rect -340 4181 -284 4253
rect -340 4129 -338 4181
rect -286 4129 -284 4181
rect -340 4057 -284 4129
rect -340 4005 -338 4057
rect -286 4005 -284 4057
rect -340 3769 -284 4005
rect -340 3717 -338 3769
rect -286 3717 -284 3769
rect -340 3645 -284 3717
rect -340 3593 -338 3645
rect -286 3593 -284 3645
rect -340 3521 -284 3593
rect -340 3469 -338 3521
rect -286 3469 -284 3521
rect -340 3233 -284 3469
rect -340 3181 -338 3233
rect -286 3181 -284 3233
rect -340 3109 -284 3181
rect -340 3057 -338 3109
rect -286 3057 -284 3109
rect -340 2985 -284 3057
rect -340 2933 -338 2985
rect -286 2933 -284 2985
rect -340 2697 -284 2933
rect -340 2645 -338 2697
rect -286 2645 -284 2697
rect -340 2573 -284 2645
rect -340 2521 -338 2573
rect -286 2521 -284 2573
rect -340 2449 -284 2521
rect -340 2397 -338 2449
rect -286 2397 -284 2449
rect -340 2161 -284 2397
rect -340 2109 -338 2161
rect -286 2109 -284 2161
rect -340 2037 -284 2109
rect -340 1985 -338 2037
rect -286 1985 -284 2037
rect -340 1913 -284 1985
rect -340 1861 -338 1913
rect -286 1861 -284 1913
rect -340 1625 -284 1861
rect -340 1573 -338 1625
rect -286 1573 -284 1625
rect -340 1501 -284 1573
rect -340 1449 -338 1501
rect -286 1449 -284 1501
rect -340 1377 -284 1449
rect -340 1325 -338 1377
rect -286 1325 -284 1377
rect -340 1089 -284 1325
rect -340 1037 -338 1089
rect -286 1037 -284 1089
rect -340 965 -284 1037
rect -340 913 -338 965
rect -286 913 -284 965
rect -340 841 -284 913
rect -340 789 -338 841
rect -286 789 -284 841
rect -340 553 -284 789
rect -340 501 -338 553
rect -286 501 -284 553
rect -340 429 -284 501
rect -340 377 -338 429
rect -286 377 -284 429
rect -340 305 -284 377
rect -340 253 -338 305
rect -286 253 -284 305
rect -340 17 -284 253
rect -340 -35 -338 17
rect -286 -35 -284 17
rect -340 -107 -284 -35
rect -340 -159 -338 -107
rect -286 -159 -284 -107
rect -340 -231 -284 -159
rect -340 -283 -338 -231
rect -286 -283 -284 -231
rect -340 -519 -284 -283
rect -340 -571 -338 -519
rect -286 -571 -284 -519
rect -340 -643 -284 -571
rect -340 -695 -338 -643
rect -286 -695 -284 -643
rect -340 -767 -284 -695
rect -340 -819 -338 -767
rect -286 -819 -284 -767
rect -340 -1055 -284 -819
rect -340 -1107 -338 -1055
rect -286 -1107 -284 -1055
rect -340 -1179 -284 -1107
rect -340 -1231 -338 -1179
rect -286 -1231 -284 -1179
rect -340 -1303 -284 -1231
rect -340 -1355 -338 -1303
rect -286 -1355 -284 -1303
rect -340 -1591 -284 -1355
rect -340 -1643 -338 -1591
rect -286 -1643 -284 -1591
rect -340 -1715 -284 -1643
rect -340 -1767 -338 -1715
rect -286 -1767 -284 -1715
rect -340 -1839 -284 -1767
rect -340 -1891 -338 -1839
rect -286 -1891 -284 -1839
rect -340 -1897 -284 -1891
rect -122 6449 -66 6455
rect -122 6397 -120 6449
rect -68 6397 -66 6449
rect -122 6325 -66 6397
rect -122 6273 -120 6325
rect -68 6273 -66 6325
rect -122 6201 -66 6273
rect -122 6149 -120 6201
rect -68 6149 -66 6201
rect -122 5913 -66 6149
rect -122 5861 -120 5913
rect -68 5861 -66 5913
rect -122 5789 -66 5861
rect -122 5737 -120 5789
rect -68 5737 -66 5789
rect -122 5665 -66 5737
rect -122 5613 -120 5665
rect -68 5613 -66 5665
rect -122 5377 -66 5613
rect -122 5325 -120 5377
rect -68 5325 -66 5377
rect -122 5253 -66 5325
rect -122 5201 -120 5253
rect -68 5201 -66 5253
rect -122 5129 -66 5201
rect -122 5077 -120 5129
rect -68 5077 -66 5129
rect -122 4841 -66 5077
rect -122 4789 -120 4841
rect -68 4789 -66 4841
rect -122 4717 -66 4789
rect -122 4665 -120 4717
rect -68 4665 -66 4717
rect -122 4593 -66 4665
rect -122 4541 -120 4593
rect -68 4541 -66 4593
rect -122 4305 -66 4541
rect -122 4253 -120 4305
rect -68 4253 -66 4305
rect -122 4181 -66 4253
rect -122 4129 -120 4181
rect -68 4129 -66 4181
rect -122 4057 -66 4129
rect -122 4005 -120 4057
rect -68 4005 -66 4057
rect -122 3769 -66 4005
rect -122 3717 -120 3769
rect -68 3717 -66 3769
rect -122 3645 -66 3717
rect -122 3593 -120 3645
rect -68 3593 -66 3645
rect -122 3521 -66 3593
rect -122 3469 -120 3521
rect -68 3469 -66 3521
rect -122 3233 -66 3469
rect -122 3181 -120 3233
rect -68 3181 -66 3233
rect -122 3109 -66 3181
rect -122 3057 -120 3109
rect -68 3057 -66 3109
rect -122 2985 -66 3057
rect -122 2933 -120 2985
rect -68 2933 -66 2985
rect -122 2697 -66 2933
rect -122 2645 -120 2697
rect -68 2645 -66 2697
rect -122 2573 -66 2645
rect -122 2521 -120 2573
rect -68 2521 -66 2573
rect -122 2449 -66 2521
rect -122 2397 -120 2449
rect -68 2397 -66 2449
rect -122 2161 -66 2397
rect -122 2109 -120 2161
rect -68 2109 -66 2161
rect -122 2037 -66 2109
rect -122 1985 -120 2037
rect -68 1985 -66 2037
rect -122 1913 -66 1985
rect -122 1861 -120 1913
rect -68 1861 -66 1913
rect -122 1625 -66 1861
rect -122 1573 -120 1625
rect -68 1573 -66 1625
rect -122 1501 -66 1573
rect -122 1449 -120 1501
rect -68 1449 -66 1501
rect -122 1377 -66 1449
rect -122 1325 -120 1377
rect -68 1325 -66 1377
rect -122 1089 -66 1325
rect -122 1037 -120 1089
rect -68 1037 -66 1089
rect -122 965 -66 1037
rect -122 913 -120 965
rect -68 913 -66 965
rect -122 841 -66 913
rect -122 789 -120 841
rect -68 789 -66 841
rect -122 553 -66 789
rect -122 501 -120 553
rect -68 501 -66 553
rect -122 429 -66 501
rect -122 377 -120 429
rect -68 377 -66 429
rect -122 305 -66 377
rect -122 253 -120 305
rect -68 253 -66 305
rect -122 17 -66 253
rect -122 -35 -120 17
rect -68 -35 -66 17
rect -122 -107 -66 -35
rect -122 -159 -120 -107
rect -68 -159 -66 -107
rect -122 -231 -66 -159
rect -122 -283 -120 -231
rect -68 -283 -66 -231
rect -122 -519 -66 -283
rect -122 -571 -120 -519
rect -68 -571 -66 -519
rect -122 -643 -66 -571
rect -122 -695 -120 -643
rect -68 -695 -66 -643
rect -122 -767 -66 -695
rect -122 -819 -120 -767
rect -68 -819 -66 -767
rect -122 -1055 -66 -819
rect -122 -1107 -120 -1055
rect -68 -1107 -66 -1055
rect -122 -1179 -66 -1107
rect -122 -1231 -120 -1179
rect -68 -1231 -66 -1179
rect -122 -1303 -66 -1231
rect -122 -1355 -120 -1303
rect -68 -1355 -66 -1303
rect -122 -1591 -66 -1355
rect -122 -1643 -120 -1591
rect -68 -1643 -66 -1591
rect -122 -1715 -66 -1643
rect -122 -1767 -120 -1715
rect -68 -1767 -66 -1715
rect -122 -1839 -66 -1767
rect -122 -1891 -120 -1839
rect -68 -1891 -66 -1839
rect -122 -1897 -66 -1891
rect -38 6111 18 6487
rect -38 6059 -36 6111
rect 16 6059 18 6111
rect -38 6003 18 6059
rect -38 5951 -36 6003
rect 16 5951 18 6003
rect -38 5575 18 5951
rect -38 5523 -36 5575
rect 16 5523 18 5575
rect -38 5467 18 5523
rect -38 5415 -36 5467
rect 16 5415 18 5467
rect -38 5039 18 5415
rect -38 4987 -36 5039
rect 16 4987 18 5039
rect -38 4931 18 4987
rect -38 4879 -36 4931
rect 16 4879 18 4931
rect -38 4503 18 4879
rect -38 4451 -36 4503
rect 16 4451 18 4503
rect -38 4395 18 4451
rect -38 4343 -36 4395
rect 16 4343 18 4395
rect -38 3967 18 4343
rect -38 3915 -36 3967
rect 16 3915 18 3967
rect -38 3859 18 3915
rect -38 3807 -36 3859
rect 16 3807 18 3859
rect -38 3431 18 3807
rect -38 3379 -36 3431
rect 16 3379 18 3431
rect -38 3323 18 3379
rect -38 3271 -36 3323
rect 16 3271 18 3323
rect -38 2895 18 3271
rect -38 2843 -36 2895
rect 16 2843 18 2895
rect -38 2787 18 2843
rect -38 2735 -36 2787
rect 16 2735 18 2787
rect -38 2359 18 2735
rect -38 2307 -36 2359
rect 16 2307 18 2359
rect -38 2251 18 2307
rect -38 2199 -36 2251
rect 16 2199 18 2251
rect -38 1823 18 2199
rect -38 1771 -36 1823
rect 16 1771 18 1823
rect -38 1715 18 1771
rect -38 1663 -36 1715
rect 16 1663 18 1715
rect -38 1287 18 1663
rect -38 1235 -36 1287
rect 16 1235 18 1287
rect -38 1179 18 1235
rect -38 1127 -36 1179
rect 16 1127 18 1179
rect -38 751 18 1127
rect -38 699 -36 751
rect 16 699 18 751
rect -38 643 18 699
rect -38 591 -36 643
rect 16 591 18 643
rect -38 215 18 591
rect -38 163 -36 215
rect 16 163 18 215
rect -38 107 18 163
rect -38 55 -36 107
rect 16 55 18 107
rect -38 -321 18 55
rect -38 -373 -36 -321
rect 16 -373 18 -321
rect -38 -429 18 -373
rect -38 -481 -36 -429
rect 16 -481 18 -429
rect -38 -857 18 -481
rect -38 -909 -36 -857
rect 16 -909 18 -857
rect -38 -965 18 -909
rect -38 -1017 -36 -965
rect 16 -1017 18 -965
rect -38 -1393 18 -1017
rect -38 -1445 -36 -1393
rect 16 -1445 18 -1393
rect -38 -1501 18 -1445
rect -38 -1553 -36 -1501
rect 16 -1553 18 -1501
rect -424 -1981 -422 -1929
rect -370 -1981 -368 -1929
rect -424 -2009 -368 -1981
rect -38 -1929 18 -1553
rect 46 6449 102 6455
rect 46 6397 48 6449
rect 100 6397 102 6449
rect 46 6325 102 6397
rect 46 6273 48 6325
rect 100 6273 102 6325
rect 46 6201 102 6273
rect 46 6149 48 6201
rect 100 6149 102 6201
rect 46 5913 102 6149
rect 46 5861 48 5913
rect 100 5861 102 5913
rect 46 5789 102 5861
rect 46 5737 48 5789
rect 100 5737 102 5789
rect 46 5665 102 5737
rect 46 5613 48 5665
rect 100 5613 102 5665
rect 46 5377 102 5613
rect 46 5325 48 5377
rect 100 5325 102 5377
rect 46 5253 102 5325
rect 46 5201 48 5253
rect 100 5201 102 5253
rect 46 5129 102 5201
rect 46 5077 48 5129
rect 100 5077 102 5129
rect 46 4841 102 5077
rect 46 4789 48 4841
rect 100 4789 102 4841
rect 46 4717 102 4789
rect 46 4665 48 4717
rect 100 4665 102 4717
rect 46 4593 102 4665
rect 46 4541 48 4593
rect 100 4541 102 4593
rect 46 4305 102 4541
rect 46 4253 48 4305
rect 100 4253 102 4305
rect 46 4181 102 4253
rect 46 4129 48 4181
rect 100 4129 102 4181
rect 46 4057 102 4129
rect 46 4005 48 4057
rect 100 4005 102 4057
rect 46 3769 102 4005
rect 46 3717 48 3769
rect 100 3717 102 3769
rect 46 3645 102 3717
rect 46 3593 48 3645
rect 100 3593 102 3645
rect 46 3521 102 3593
rect 46 3469 48 3521
rect 100 3469 102 3521
rect 46 3233 102 3469
rect 46 3181 48 3233
rect 100 3181 102 3233
rect 46 3109 102 3181
rect 46 3057 48 3109
rect 100 3057 102 3109
rect 46 2985 102 3057
rect 46 2933 48 2985
rect 100 2933 102 2985
rect 454 3051 510 3057
rect 454 2999 456 3051
rect 508 2999 510 3051
rect 46 2697 102 2933
rect 46 2645 48 2697
rect 100 2645 102 2697
rect 46 2573 102 2645
rect 46 2521 48 2573
rect 100 2521 102 2573
rect 46 2449 102 2521
rect 46 2397 48 2449
rect 100 2397 102 2449
rect 46 2161 102 2397
rect 46 2109 48 2161
rect 100 2109 102 2161
rect 46 2037 102 2109
rect 46 1985 48 2037
rect 100 1985 102 2037
rect 46 1913 102 1985
rect 46 1861 48 1913
rect 100 1861 102 1913
rect 46 1625 102 1861
rect 46 1573 48 1625
rect 100 1573 102 1625
rect 46 1501 102 1573
rect 46 1449 48 1501
rect 100 1449 102 1501
rect 46 1377 102 1449
rect 46 1325 48 1377
rect 100 1325 102 1377
rect 46 1089 102 1325
rect 46 1037 48 1089
rect 100 1037 102 1089
rect 46 965 102 1037
rect 46 913 48 965
rect 100 913 102 965
rect 46 841 102 913
rect 46 789 48 841
rect 100 789 102 841
rect 46 553 102 789
rect 46 501 48 553
rect 100 501 102 553
rect 46 429 102 501
rect 46 377 48 429
rect 100 377 102 429
rect 46 305 102 377
rect 46 253 48 305
rect 100 253 102 305
rect 46 17 102 253
rect 46 -35 48 17
rect 100 -35 102 17
rect 46 -107 102 -35
rect 46 -159 48 -107
rect 100 -159 102 -107
rect 46 -231 102 -159
rect 46 -283 48 -231
rect 100 -283 102 -231
rect 46 -519 102 -283
rect 46 -571 48 -519
rect 100 -571 102 -519
rect 46 -643 102 -571
rect 46 -695 48 -643
rect 100 -695 102 -643
rect 46 -767 102 -695
rect 46 -819 48 -767
rect 100 -819 102 -767
rect 46 -1055 102 -819
rect 46 -1107 48 -1055
rect 100 -1107 102 -1055
rect 46 -1179 102 -1107
rect 46 -1231 48 -1179
rect 100 -1231 102 -1179
rect 46 -1303 102 -1231
rect 46 -1355 48 -1303
rect 100 -1355 102 -1303
rect 46 -1591 102 -1355
rect 46 -1643 48 -1591
rect 100 -1643 102 -1591
rect 46 -1715 102 -1643
rect 46 -1767 48 -1715
rect 100 -1767 102 -1715
rect 46 -1839 102 -1767
rect 46 -1891 48 -1839
rect 100 -1891 102 -1839
rect 46 -1897 102 -1891
rect 370 2922 426 2976
rect 370 2870 372 2922
rect 424 2870 426 2922
rect 370 2604 426 2870
rect 370 2552 372 2604
rect 424 2552 426 2604
rect 370 2286 426 2552
rect 370 2234 372 2286
rect 424 2234 426 2286
rect 370 1968 426 2234
rect 370 1916 372 1968
rect 424 1916 426 1968
rect 370 1650 426 1916
rect 370 1598 372 1650
rect 424 1598 426 1650
rect 370 1332 426 1598
rect 370 1280 372 1332
rect 424 1280 426 1332
rect 370 1014 426 1280
rect 370 962 372 1014
rect 424 962 426 1014
rect 370 696 426 962
rect 370 644 372 696
rect 424 644 426 696
rect 370 378 426 644
rect 370 326 372 378
rect 424 326 426 378
rect 370 60 426 326
rect 370 8 372 60
rect 424 8 426 60
rect 370 -258 426 8
rect 370 -310 372 -258
rect 424 -310 426 -258
rect 370 -576 426 -310
rect 370 -628 372 -576
rect 424 -628 426 -576
rect 370 -894 426 -628
rect 370 -946 372 -894
rect 424 -946 426 -894
rect 370 -1212 426 -946
rect 370 -1264 372 -1212
rect 424 -1264 426 -1212
rect 370 -1530 426 -1264
rect 370 -1582 372 -1530
rect 424 -1582 426 -1530
rect 370 -1848 426 -1582
rect 370 -1900 372 -1848
rect 424 -1900 426 -1848
rect 370 -1906 426 -1900
rect 454 2841 510 2999
rect 840 3051 896 3057
rect 840 2999 842 3051
rect 894 2999 896 3051
rect 454 2789 456 2841
rect 508 2789 510 2841
rect 454 2733 510 2789
rect 454 2681 456 2733
rect 508 2681 510 2733
rect 454 2523 510 2681
rect 454 2471 456 2523
rect 508 2471 510 2523
rect 454 2415 510 2471
rect 454 2363 456 2415
rect 508 2363 510 2415
rect 454 2205 510 2363
rect 454 2153 456 2205
rect 508 2153 510 2205
rect 454 2097 510 2153
rect 454 2045 456 2097
rect 508 2045 510 2097
rect 454 1887 510 2045
rect 454 1835 456 1887
rect 508 1835 510 1887
rect 454 1779 510 1835
rect 454 1727 456 1779
rect 508 1727 510 1779
rect 454 1569 510 1727
rect 454 1517 456 1569
rect 508 1517 510 1569
rect 454 1461 510 1517
rect 454 1409 456 1461
rect 508 1409 510 1461
rect 454 1251 510 1409
rect 454 1199 456 1251
rect 508 1199 510 1251
rect 454 1143 510 1199
rect 454 1091 456 1143
rect 508 1091 510 1143
rect 454 933 510 1091
rect 454 881 456 933
rect 508 881 510 933
rect 454 825 510 881
rect 454 773 456 825
rect 508 773 510 825
rect 454 615 510 773
rect 454 563 456 615
rect 508 563 510 615
rect 454 507 510 563
rect 454 455 456 507
rect 508 455 510 507
rect 454 297 510 455
rect 454 245 456 297
rect 508 245 510 297
rect 454 189 510 245
rect 454 137 456 189
rect 508 137 510 189
rect 454 -21 510 137
rect 454 -73 456 -21
rect 508 -73 510 -21
rect 454 -129 510 -73
rect 454 -181 456 -129
rect 508 -181 510 -129
rect 454 -339 510 -181
rect 454 -391 456 -339
rect 508 -391 510 -339
rect 454 -447 510 -391
rect 454 -499 456 -447
rect 508 -499 510 -447
rect 454 -657 510 -499
rect 454 -709 456 -657
rect 508 -709 510 -657
rect 454 -765 510 -709
rect 454 -817 456 -765
rect 508 -817 510 -765
rect 454 -975 510 -817
rect 454 -1027 456 -975
rect 508 -1027 510 -975
rect 454 -1083 510 -1027
rect 454 -1135 456 -1083
rect 508 -1135 510 -1083
rect 454 -1293 510 -1135
rect 454 -1345 456 -1293
rect 508 -1345 510 -1293
rect 454 -1401 510 -1345
rect 454 -1453 456 -1401
rect 508 -1453 510 -1401
rect 454 -1611 510 -1453
rect 454 -1663 456 -1611
rect 508 -1663 510 -1611
rect 454 -1719 510 -1663
rect 454 -1771 456 -1719
rect 508 -1771 510 -1719
rect -38 -1981 -36 -1929
rect 16 -1981 18 -1929
rect -38 -1987 18 -1981
rect 454 -1929 510 -1771
rect 538 2922 594 2976
rect 538 2870 540 2922
rect 592 2870 594 2922
rect 538 2604 594 2870
rect 538 2552 540 2604
rect 592 2552 594 2604
rect 538 2286 594 2552
rect 538 2234 540 2286
rect 592 2234 594 2286
rect 538 1968 594 2234
rect 538 1916 540 1968
rect 592 1916 594 1968
rect 538 1650 594 1916
rect 538 1598 540 1650
rect 592 1598 594 1650
rect 538 1332 594 1598
rect 538 1280 540 1332
rect 592 1280 594 1332
rect 538 1014 594 1280
rect 538 962 540 1014
rect 592 962 594 1014
rect 538 696 594 962
rect 538 644 540 696
rect 592 644 594 696
rect 538 378 594 644
rect 538 326 540 378
rect 592 326 594 378
rect 538 60 594 326
rect 538 8 540 60
rect 592 8 594 60
rect 538 -258 594 8
rect 538 -310 540 -258
rect 592 -310 594 -258
rect 538 -576 594 -310
rect 538 -628 540 -576
rect 592 -628 594 -576
rect 538 -894 594 -628
rect 538 -946 540 -894
rect 592 -946 594 -894
rect 538 -1212 594 -946
rect 538 -1264 540 -1212
rect 592 -1264 594 -1212
rect 538 -1530 594 -1264
rect 538 -1582 540 -1530
rect 592 -1582 594 -1530
rect 538 -1848 594 -1582
rect 538 -1900 540 -1848
rect 592 -1900 594 -1848
rect 538 -1906 594 -1900
rect 756 2922 812 2976
rect 756 2870 758 2922
rect 810 2870 812 2922
rect 756 2604 812 2870
rect 756 2552 758 2604
rect 810 2552 812 2604
rect 756 2286 812 2552
rect 756 2234 758 2286
rect 810 2234 812 2286
rect 756 1968 812 2234
rect 756 1916 758 1968
rect 810 1916 812 1968
rect 756 1650 812 1916
rect 756 1598 758 1650
rect 810 1598 812 1650
rect 756 1332 812 1598
rect 756 1280 758 1332
rect 810 1280 812 1332
rect 756 1014 812 1280
rect 756 962 758 1014
rect 810 962 812 1014
rect 756 696 812 962
rect 756 644 758 696
rect 810 644 812 696
rect 756 378 812 644
rect 756 326 758 378
rect 810 326 812 378
rect 756 60 812 326
rect 756 8 758 60
rect 810 8 812 60
rect 756 -258 812 8
rect 756 -310 758 -258
rect 810 -310 812 -258
rect 756 -576 812 -310
rect 756 -628 758 -576
rect 810 -628 812 -576
rect 756 -894 812 -628
rect 756 -946 758 -894
rect 810 -946 812 -894
rect 756 -1212 812 -946
rect 756 -1264 758 -1212
rect 810 -1264 812 -1212
rect 756 -1530 812 -1264
rect 756 -1582 758 -1530
rect 810 -1582 812 -1530
rect 756 -1848 812 -1582
rect 756 -1900 758 -1848
rect 810 -1900 812 -1848
rect 756 -1906 812 -1900
rect 840 2841 896 2999
rect 840 2789 842 2841
rect 894 2789 896 2841
rect 840 2733 896 2789
rect 840 2681 842 2733
rect 894 2681 896 2733
rect 840 2523 896 2681
rect 840 2471 842 2523
rect 894 2471 896 2523
rect 840 2415 896 2471
rect 840 2363 842 2415
rect 894 2363 896 2415
rect 840 2205 896 2363
rect 840 2153 842 2205
rect 894 2153 896 2205
rect 840 2097 896 2153
rect 840 2045 842 2097
rect 894 2045 896 2097
rect 840 1887 896 2045
rect 840 1835 842 1887
rect 894 1835 896 1887
rect 840 1779 896 1835
rect 840 1727 842 1779
rect 894 1727 896 1779
rect 840 1569 896 1727
rect 840 1517 842 1569
rect 894 1517 896 1569
rect 840 1461 896 1517
rect 840 1409 842 1461
rect 894 1409 896 1461
rect 840 1251 896 1409
rect 840 1199 842 1251
rect 894 1199 896 1251
rect 840 1143 896 1199
rect 840 1091 842 1143
rect 894 1091 896 1143
rect 840 933 896 1091
rect 840 881 842 933
rect 894 881 896 933
rect 840 825 896 881
rect 840 773 842 825
rect 894 773 896 825
rect 840 615 896 773
rect 840 563 842 615
rect 894 563 896 615
rect 840 507 896 563
rect 840 455 842 507
rect 894 455 896 507
rect 840 297 896 455
rect 840 245 842 297
rect 894 245 896 297
rect 840 189 896 245
rect 840 137 842 189
rect 894 137 896 189
rect 840 -21 896 137
rect 840 -73 842 -21
rect 894 -73 896 -21
rect 840 -129 896 -73
rect 840 -181 842 -129
rect 894 -181 896 -129
rect 840 -339 896 -181
rect 840 -391 842 -339
rect 894 -391 896 -339
rect 840 -447 896 -391
rect 840 -499 842 -447
rect 894 -499 896 -447
rect 840 -657 896 -499
rect 840 -709 842 -657
rect 894 -709 896 -657
rect 840 -765 896 -709
rect 840 -817 842 -765
rect 894 -817 896 -765
rect 840 -975 896 -817
rect 840 -1027 842 -975
rect 894 -1027 896 -975
rect 840 -1083 896 -1027
rect 840 -1135 842 -1083
rect 894 -1135 896 -1083
rect 840 -1293 896 -1135
rect 840 -1345 842 -1293
rect 894 -1345 896 -1293
rect 840 -1401 896 -1345
rect 840 -1453 842 -1401
rect 894 -1453 896 -1401
rect 840 -1611 896 -1453
rect 840 -1663 842 -1611
rect 894 -1663 896 -1611
rect 840 -1719 896 -1663
rect 840 -1771 842 -1719
rect 894 -1771 896 -1719
rect 454 -1981 456 -1929
rect 508 -1981 510 -1929
rect 454 -1987 510 -1981
rect 840 -1929 896 -1771
rect 840 -1981 842 -1929
rect 894 -1981 896 -1929
rect -424 -2061 -422 -2009
rect -370 -2061 -368 -2009
rect -424 -2067 -368 -2061
rect 840 -2009 896 -1981
rect 840 -2061 842 -2009
rect 894 -2061 896 -2009
rect 840 -2067 896 -2061
rect 924 2922 980 2976
rect 924 2870 926 2922
rect 978 2870 980 2922
rect 924 2604 980 2870
rect 924 2552 926 2604
rect 978 2552 980 2604
rect 924 2286 980 2552
rect 924 2234 926 2286
rect 978 2234 980 2286
rect 924 1968 980 2234
rect 924 1916 926 1968
rect 978 1916 980 1968
rect 924 1650 980 1916
rect 924 1598 926 1650
rect 978 1598 980 1650
rect 924 1332 980 1598
rect 924 1280 926 1332
rect 978 1280 980 1332
rect 924 1014 980 1280
rect 924 962 926 1014
rect 978 962 980 1014
rect 924 696 980 962
rect 924 644 926 696
rect 978 644 980 696
rect 924 378 980 644
rect 924 326 926 378
rect 978 326 980 378
rect 924 60 980 326
rect 924 8 926 60
rect 978 8 980 60
rect 924 -258 980 8
rect 924 -310 926 -258
rect 978 -310 980 -258
rect 924 -576 980 -310
rect 924 -628 926 -576
rect 978 -628 980 -576
rect 924 -894 980 -628
rect 924 -946 926 -894
rect 978 -946 980 -894
rect 924 -1212 980 -946
rect 924 -1264 926 -1212
rect 978 -1264 980 -1212
rect 924 -1530 980 -1264
rect 924 -1582 926 -1530
rect 978 -1582 980 -1530
rect 924 -1848 980 -1582
rect 924 -1900 926 -1848
rect 978 -1900 980 -1848
rect -508 -2200 -506 -2110
rect -454 -2200 -452 -2110
rect -508 -2206 -452 -2200
rect 924 -2234 980 -1900
rect 924 -2324 926 -2234
rect 978 -2324 980 -2234
rect 924 -2330 980 -2324
use sky130_fd_pr__pfet_01v8_GN49S6  XM1
timestamp 1730624594
transform 1 0 -396 0 1 2279
box -246 -4389 246 4389
use sky130_fd_pr__pfet_01v8_GN49S6  XM2
timestamp 1730624594
transform 1 0 -10 0 1 2279
box -246 -4389 246 4389
use sky130_fd_pr__nfet_01v8_GPU48F  XM3
timestamp 1730624594
transform 1 0 482 0 1 535
box -246 -2645 246 2645
use sky130_fd_pr__nfet_01v8_GPU48F  XM4
timestamp 1730624594
transform 1 0 868 0 1 535
box -246 -2645 246 2645
<< labels >>
flabel metal1 -642 -2206 -546 -2110 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel metal1 -642 -2330 -546 -2234 0 FreeSans 320 0 0 0 vssa
port 5 nsew
flabel via1 -36 -1981 16 -1929 0 FreeSans 320 0 0 0 ckb
port 4 nsew
flabel via1 456 -1981 508 -1929 0 FreeSans 320 0 0 0 ck
port 3 nsew
flabel via1 842 2999 894 3051 0 FreeSans 320 0 0 0 in
port 2 nsew
flabel via1 48 6397 100 6449 0 FreeSans 320 0 0 0 out
port 6 nsew
<< end >>
