* PEX produced on Sel 05 Nov 2024 03:02:51  CST using ./iic-pex.sh with m=1 and s=1
* NGSPICE file created from cdac_10b.ext - technology: sky130A

X0 a_55274_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 a_10649_24944# single_10b_cdac_1.cdac_sw_8_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 single_10b_cdac_1.x10b_cap_array_0.SW[4] single_10b_cdac_1.cdac_sw_4_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x9.A single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 VSREF single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 single_10b_cdac_0.x8[7].dac_out single_10b_cdac_0.x8[7].x3.ck a_42394_34645# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X10 single_10b_cdac_0.x6[4].dac_out single_10b_cdac_0.x6[4].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X11 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X13 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x3.ckb a_10556_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X14 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 single_10b_cdac_0.cdac_sw_8_1.x1.x6.A single_10b_cdac_0.cdac_sw_8_1.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X18 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X19 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.cdac_sw_2_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VSREF single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.cdac_sw_4_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X25 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.cdac_sw_8_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X30 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 VSREF single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X34 a_14654_25713# single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X35 VDREF single_10b_cdac_0.x3[0].x1.x6.A single_10b_cdac_0.x3[0].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X36 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 VDREF CF[9] single_10b_cdac_1.cdac_sw_1_2.x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X38 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X40 single_10b_cdac_0.x4[2].x2.swn single_10b_cdac_0.x4[2].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X42 single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.cdac_sw_2_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X43 VDREF single_10b_cdac_0.x6[5].x1.x9.A single_10b_cdac_0.x6[5].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 VSREF single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X47 single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X49 VDREF single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X50 a_16118_33146# single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X51 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X54 single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 single_10b_cdac_1.x10[8].x3.ck single_10b_cdac_1.x10[8].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X56 single_10b_cdac_1.x8[6].x3.ck single_10b_cdac_1.x8[6].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X57 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 VDREF single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 single_10b_cdac_1.cdac_sw_16_0.x1.x6.A single_10b_cdac_1.cdac_sw_16_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X60 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 VDREF single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X63 single_10b_cdac_1.x3[0].x3.ck single_10b_cdac_1.x3[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X64 VCM single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X65 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 single_10b_cdac_1.x8[6].x2.swn single_10b_cdac_1.x8[6].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X68 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X69 single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X70 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X71 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X74 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X79 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VSREF single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X85 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X86 single_10b_cdac_1.x3[0].x1.x4.A CF[0] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X87 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X89 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 single_10b_cdac_0.cdac_sw_16_0.x1.x7.A single_10b_cdac_0.cdac_sw_16_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X91 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x9.A single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X92 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 VSREF SWN_IN[4] a_48248_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X94 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X95 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X98 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 a_57908_25713# single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[7] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X100 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 VDREF single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X102 single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X103 single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X104 VSREF single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X105 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X107 single_10b_cdac_0.cdac_sw_1_0.x1.x5.A single_10b_cdac_0.cdac_sw_1_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X108 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 single_10b_cdac_1.cdac_sw_1_2.x2.swn single_10b_cdac_1.cdac_sw_1_2.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X111 single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X112 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 a_48834_34009# SWP_IN[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X115 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X117 single_10b_cdac_0.x2[0].x1.x3.Y CF[1] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X118 single_10b_cdac_1.x8[7].dac_out single_10b_cdac_1.x8[7].x3.ck a_8800_34645# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X119 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X121 VSREF SWN_IN[5] a_17874_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X122 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X123 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X127 VSREF single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X128 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VSREF single_10b_cdac_1.x8[6].x1.x4.A single_10b_cdac_1.x8[6].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X130 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X132 VDREF single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X133 VCM single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X134 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 a_39174_34963# SWP_IN[8] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X136 VSREF single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X137 a_19338_33146# single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X138 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x2[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X140 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X141 a_18460_34009# SWP_IN[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X142 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 VSREF single_10b_cdac_0.x8[7].x1.x9.A a_43411_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X145 single_10b_cdac_1.cdac_sw_1_2.x3.ck single_10b_cdac_1.cdac_sw_1_2.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X146 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X148 VDREF single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X149 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X150 VSREF single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X151 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X153 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X155 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 VDREF single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X158 VCM single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X159 single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X160 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X161 VDREF single_10b_cdac_0.x3[1].x1.x8.A single_10b_cdac_0.x3[1].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X162 VSREF single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X163 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VCM single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X166 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 single_10b_cdac_0.x10b_cap_array_0.SW[5] single_10b_cdac_0.cdac_sw_4_0.x3.ckb a_50590_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X169 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X170 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 VDREF single_10b_cdac_1.x6[5].x1.x9.A single_10b_cdac_1.x6[5].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X172 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X174 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.cdac_sw_4_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X177 VDREF single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X178 VDREF CF[0] single_10b_cdac_1.cdac_sw_16_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X179 single_10b_cdac_1.x4[3].x3.ck single_10b_cdac_1.x4[3].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X180 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X182 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X184 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 single_10b_cdac_0.cdac_sw_4_1.x1.x9.A single_10b_cdac_0.cdac_sw_4_1.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X187 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X190 single_10b_cdac_1.cdac_sw_1_1.x2.swn single_10b_cdac_1.cdac_sw_1_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X191 VCM single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X192 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X197 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 VSREF single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X200 single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.cdac_sw_8_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X201 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X206 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X208 single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.cdac_sw_2_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X209 VSREF single_10b_cdac_1.x3[0].x1.x9.A single_10b_cdac_1.x3[0].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X210 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x4.A single_10b_cdac_1.cdac_sw_1_2.x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X213 VSREF single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X214 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 a_64348_25713# single_10b_cdac_0.cdac_sw_1_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[9] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X225 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VSREF single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X228 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x8.A single_10b_cdac_1.cdac_sw_4_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X230 single_10b_cdac_0.x8[7].x2.swn single_10b_cdac_0.x8[7].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X231 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X233 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 VSREF single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X237 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X240 VSREF single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X241 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 single_10b_cdac_0.cdac_sw_4_0.x1.x5.A single_10b_cdac_0.cdac_sw_4_0.x1.x8.A a_50683_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X244 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X246 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X248 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 single_10b_cdac_0.cdac_sw_1_1.x3.ck single_10b_cdac_0.cdac_sw_1_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X251 single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.cdac_sw_8_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X252 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X253 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.cdac_sw_16_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X257 single_10b_cdac_1.x6[5].x3.ck single_10b_cdac_1.x6[5].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X258 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 a_59372_31002# single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X260 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 VDREF single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X262 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 single_10b_cdac_0.x4[3].x1.x5.A single_10b_cdac_0.x4[3].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X266 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X267 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 VCP single_10b_cdac_0.x3[1].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VCM single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X270 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X271 single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X272 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X275 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X278 VSREF single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X279 single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 VCM single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X281 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X282 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 VSREF single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X288 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X291 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 single_10b_cdac_1.x3[1].x3.ck single_10b_cdac_1.x3[1].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X293 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X294 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X296 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X297 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x8.A single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X299 single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X300 single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X301 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.cdac_sw_4_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X304 single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X305 VSREF single_10b_cdac_1.x4[2].x1.x9.A single_10b_cdac_1.x4[2].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X306 single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X307 VDREF single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X308 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x2[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X311 VDREF single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X312 a_41808_25713# single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X313 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VDREF single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X316 single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X317 single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.cdac_sw_4_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X318 VSREF single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X319 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x3.ck a_21680_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X325 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 single_10b_cdac_1.cdac_sw_1_2.dac_out single_10b_cdac_1.cdac_sw_1_2.x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X327 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X329 single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X330 VSREF single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X331 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 VSREF single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X334 VSREF single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X335 VDREF single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X336 single_10b_cdac_0.x8[6].x2.swn single_10b_cdac_0.x8[6].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X337 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X338 a_59372_31002# single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X339 single_10b_cdac_1.cdac_sw_2_0.x1.x5.A single_10b_cdac_1.cdac_sw_2_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X340 single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X341 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X344 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X347 VSREF single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X348 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X351 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X353 single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X354 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x8.A single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X356 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 single_10b_cdac_0.cdac_sw_2_1.x1.x7.A single_10b_cdac_0.cdac_sw_2_1.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X358 single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.cdac_sw_8_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X359 single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X360 VDREF single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X361 a_44150_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X362 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X366 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X367 single_10b_cdac_1.cdac_sw_1_0.x1.x3.Y CF[9] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X368 single_10b_cdac_0.cdac_sw_4_0.x1.x4.A single_10b_cdac_0.cdac_sw_4_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X369 VSREF SWN_IN[2] a_8214_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X370 VCM single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X371 VDREF SWP_IN[3] a_22558_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X372 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 VDREF single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X374 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 VDREF single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X381 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X385 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X387 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 a_9817_36566# single_10b_cdac_1.x8[7].x1.x8.A single_10b_cdac_1.x8[7].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X389 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X390 single_10b_cdac_1.cdac_sw_1_0.x2.swn single_10b_cdac_1.cdac_sw_1_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X391 single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X392 VCM single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X393 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X396 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X398 single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X399 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X400 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 VSREF single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X403 single_10b_cdac_0.x2[0].x1.x9.A single_10b_cdac_0.x2[0].x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X404 VSREF CF[3] single_10b_cdac_1.x4[3].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X405 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 VDREF single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X409 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VSREF single_10b_cdac_0.x10[8].x1.x9.A single_10b_cdac_0.x10[8].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X412 VDREF single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X413 single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.cdac_sw_8_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X414 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X420 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x9.A single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X421 VDREF single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X422 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X425 VSREF SWN_IN[7] a_24314_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X426 single_10b_cdac_0.x8[6].dac_out single_10b_cdac_0.x8[6].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X427 VDREF single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X428 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X429 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X431 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 single_10b_cdac_1.x8[7].x2.swn single_10b_cdac_1.x8[7].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X434 single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.cdac_sw_4_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X435 VSREF single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X436 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x2[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X438 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x3.ckb a_7336_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X439 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X442 single_10b_cdac_0.x6[4].x2.swn single_10b_cdac_0.x6[4].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X443 single_10b_cdac_0.x10[8].x2.swn single_10b_cdac_0.x10[8].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X444 VDREF single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X445 single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X446 single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X447 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 VSREF single_10b_cdac_0.x8[6].x1.x8.A single_10b_cdac_0.x8[6].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X450 a_58494_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X451 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.cdac_sw_4_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X453 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 VSREF single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X456 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X458 VSREF single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X459 single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X460 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X463 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X464 VDREF single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X465 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X468 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 VDREF single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X471 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X473 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X476 single_10b_cdac_1.cdac_sw_2_0.x1.x6.A single_10b_cdac_1.cdac_sw_2_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X477 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X478 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X481 VSREF single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X482 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 single_10b_cdac_0.x10[8].x2.swn single_10b_cdac_0.x10[8].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X484 VCM single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X485 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X486 a_17874_25713# single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X487 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.cdac_sw_2_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X489 VSREF single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X490 a_2360_34963# SWP_IN[9] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X491 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 single_10b_cdac_0.cdac_sw_2_0.x1.x8.A single_10b_cdac_0.cdac_sw_2_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X494 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 a_989_24080# single_10b_cdac_1.cdac_sw_16_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X501 VSREF single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X502 VSREF single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X503 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x3.ckb a_7336_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X504 single_10b_cdac_1.cdac_sw_1_0.x3.ck single_10b_cdac_1.cdac_sw_1_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X505 single_10b_cdac_0.x10[8].x1.x5.A single_10b_cdac_0.x10[8].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X506 single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X507 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X509 single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X510 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 VDREF single_10b_cdac_1.x8[7].x1.x5.A single_10b_cdac_1.x8[7].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X512 single_10b_cdac_0.x3[1].x3.ck single_10b_cdac_0.x3[1].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X513 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x9.A single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X514 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X515 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 single_10b_cdac_1.cdac_sw_1_1.x1.x9.A single_10b_cdac_1.cdac_sw_1_1.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X519 a_9678_34218# single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X520 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X521 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 VCP single_10b_cdac_0.x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 a_10556_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X524 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 single_10b_cdac_1.x8[6].x3.ck single_10b_cdac_1.x8[6].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X527 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X528 VDREF single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X529 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X530 single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X531 a_57123_24944# single_10b_cdac_0.cdac_sw_2_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X532 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X533 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x8.A single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X535 single_10b_cdac_0.x4[3].x2.swn single_10b_cdac_0.x4[3].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X536 VDREF single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X537 single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X538 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X539 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 VSREF single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X542 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X543 VSREF single_10b_cdac_1.x6[5].x1.x7.A single_10b_cdac_1.x6[5].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X544 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X545 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X547 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X549 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X552 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X553 single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X554 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X555 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 VSREF SWN_IN[9] a_30754_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X557 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 VSREF single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X559 single_10b_cdac_1.cdac_sw_2_1.x1.x4.A CF[6] a_20309_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X560 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X561 single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X562 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X564 VDREF single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X565 VSREF single_10b_cdac_0.x6[5].x1.x5.A single_10b_cdac_0.x6[5].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X566 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X567 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X568 a_43272_34218# single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X569 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X572 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X573 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 single_10b_cdac_0.cdac_sw_1_0.x1.x3.Y CF[9] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X575 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x9.A a_36971_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X576 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VCM single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X579 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X580 VSREF single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X581 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X585 a_8214_25713# single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X586 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X587 VDREF single_10b_cdac_0.x4[3].x1.x8.A single_10b_cdac_0.x4[3].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X588 VSREF single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X589 single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X590 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 a_24900_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X593 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 single_10b_cdac_1.cdac_sw_4_1.x1.x3.Y CF[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X597 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x3.ckb a_44150_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X598 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X599 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X601 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X603 single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X604 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X605 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X606 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X609 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X611 single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.cdac_sw_2_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X612 single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X613 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X614 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X616 single_10b_cdac_0.x4[3].x3.ck single_10b_cdac_0.x4[3].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X617 VSREF single_10b_cdac_1.x4[2].x1.x9.A a_25917_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X618 single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X619 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 single_10b_cdac_1.x3[0].x2.swn single_10b_cdac_1.x3[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X622 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X623 VCM single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X624 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 VDREF SWP_IN[2] a_25778_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X626 VSREF single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X627 single_10b_cdac_1.x10b_cap_array_0.SW[9] single_10b_cdac_1.cdac_sw_1_0.x3.ckb a_29876_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X628 VSREF single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X629 single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X630 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X633 single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X634 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X635 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X637 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 VSREF single_10b_cdac_1.x4[2].x1.x9.A single_10b_cdac_1.x4[2].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X640 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X643 VDREF single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X644 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X648 VSREF single_10b_cdac_1.x4[2].x1.x6.A single_10b_cdac_1.x4[2].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X649 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X650 VDREF single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X651 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 single_10b_cdac_1.cdac_sw_8_1.x1.x7.A single_10b_cdac_1.cdac_sw_8_1.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X653 single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X654 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 single_10b_cdac_1.x4[3].x3.ck single_10b_cdac_1.x4[3].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X656 a_50590_25722# SWN_IN[5] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X657 single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X658 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X662 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X664 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 single_10b_cdac_1.cdac_sw_16_0.x1.x8.A single_10b_cdac_1.cdac_sw_16_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X667 VDREF single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X668 VSREF single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X669 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X670 single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X671 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X672 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X676 VDREF single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X677 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x9.A single_10b_cdac_1.cdac_sw_1_2.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X678 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X679 VSREF single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X680 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X681 single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X682 a_21680_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X683 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X684 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 VSREF single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X686 single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X687 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X689 single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X690 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X691 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X692 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X693 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X696 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X698 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 VDREF single_10b_cdac_1.x3[0].x1.x5.A single_10b_cdac_1.x3[0].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X700 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X701 VCM single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[7] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X702 a_36971_36566# single_10b_cdac_0.cdac_sw_1_2.x1.x8.A single_10b_cdac_0.cdac_sw_1_2.x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X703 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X704 single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X705 VDREF single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X706 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X707 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.cdac_sw_4_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X709 VDREF single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X710 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 VDREF single_10b_cdac_1.x3[0].x1.x6.A single_10b_cdac_1.x3[0].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X712 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X714 single_10b_cdac_0.cdac_sw_8_1.x1.x8.A single_10b_cdac_0.cdac_sw_8_1.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X715 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X716 single_10b_cdac_1.x4[2].x2.swn single_10b_cdac_1.x4[2].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X717 single_10b_cdac_0.cdac_sw_1_1.x1.x6.A single_10b_cdac_0.cdac_sw_1_1.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X718 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X720 single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X721 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X724 VSREF single_10b_cdac_0.x2[0].x1.x8.A single_10b_cdac_0.x2[0].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X725 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X727 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x9.A single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X729 single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X730 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 VCP single_10b_cdac_1.x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X732 single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X733 VDREF single_10b_cdac_0.x3[0].x1.x4.A single_10b_cdac_0.x3[0].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X734 VSREF single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X735 single_10b_cdac_1.x2[0].x1.x5.A single_10b_cdac_1.x2[0].x1.x8.A a_4209_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X736 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 single_10b_cdac_1.cdac_sw_4_0.x1.x9.A single_10b_cdac_1.cdac_sw_4_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X738 single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X739 single_10b_cdac_1.cdac_sw_8_0.x1.x9.A single_10b_cdac_1.cdac_sw_8_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X740 a_55274_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X741 single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X742 VSREF single_10b_cdac_1.x6[4].x1.x9.A single_10b_cdac_1.x6[4].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X743 VDREF single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X744 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x9.A single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X746 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X749 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x3.ck a_55274_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X750 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X751 single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.cdac_sw_8_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X752 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X753 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X756 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X757 VDREF single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X758 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X759 single_10b_cdac_1.x6[5].dac_out single_10b_cdac_1.x6[5].x3.ck a_15240_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X760 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 single_10b_cdac_0.cdac_sw_8_0.x1.x8.A single_10b_cdac_0.cdac_sw_8_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X762 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X763 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X765 VSREF SWN_IN[2] a_41808_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X766 VSREF single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X767 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X768 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X769 single_10b_cdac_0.x10[8].x2.swn single_10b_cdac_0.x10[8].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X770 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X771 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X773 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X774 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.cdac_sw_2_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X776 VDREF single_10b_cdac_0.x2[0].x1.x8.A single_10b_cdac_0.x2[0].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X777 single_10b_cdac_1.cdac_sw_4_0.x1.x5.A single_10b_cdac_1.cdac_sw_4_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X778 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X779 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X780 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X781 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X782 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X784 VSREF SWN_IN[4] a_14654_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X785 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X786 VDREF single_10b_cdac_0.x6[4].x1.x7.A single_10b_cdac_0.x6[4].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X787 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X788 single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X789 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X790 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X791 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X792 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X793 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X794 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X795 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X796 VSREF single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X797 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X798 a_41808_25713# single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X799 single_10b_cdac_0.cdac_sw_8_0.x1.x4.A single_10b_cdac_0.cdac_sw_8_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X800 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X801 single_10b_cdac_0.x8[7].x2.swn single_10b_cdac_0.x8[7].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X802 VDREF SWP_IN[5] a_16118_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X803 VCM single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X804 VDREF single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X805 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X806 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X807 single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x2[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X808 single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X809 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X810 single_10b_cdac_0.cdac_sw_1_1.x1.x8.A single_10b_cdac_0.cdac_sw_1_1.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X811 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X812 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X813 single_10b_cdac_1.x3[1].x2.swn single_10b_cdac_1.x3[1].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X814 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X815 single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X816 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X817 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X818 single_10b_cdac_1.x6[4].x2.swn single_10b_cdac_1.x6[4].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X819 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x8.A single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X820 VCN single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X821 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x5.A single_10b_cdac_0.cdac_sw_1_2.x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X822 single_10b_cdac_0.cdac_sw_1_0.x2.swn single_10b_cdac_0.cdac_sw_1_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X823 VSREF CF[5] single_10b_cdac_1.x6[5].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X824 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X825 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X826 a_22558_31002# single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X827 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X828 VSREF single_10b_cdac_0.x6[4].x1.x8.A single_10b_cdac_0.x6[4].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X829 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X830 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X831 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X832 a_36832_34754# single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X833 single_10b_cdac_1.cdac_sw_1_0.x1.x7.A single_10b_cdac_1.cdac_sw_1_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X834 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X835 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X836 VSREF single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X837 VDREF single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X838 single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.cdac_sw_8_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X839 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X840 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X841 a_60343_24944# single_10b_cdac_0.cdac_sw_1_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X842 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x9.A single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X843 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X844 VDREF single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X845 VSREF single_10b_cdac_1.x3[1].x1.x8.A single_10b_cdac_1.x3[1].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X846 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X847 VDREF single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X848 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X849 VSREF single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X850 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X851 VSREF single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X852 single_10b_cdac_0.x6[4].x3.ck single_10b_cdac_0.x6[4].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X853 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X854 single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X855 single_10b_cdac_1.x10[8].x2.swn single_10b_cdac_1.x10[8].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X856 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X857 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X858 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X859 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X860 VSREF single_10b_cdac_0.x6[4].x1.x5.A single_10b_cdac_0.x6[4].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X861 single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X862 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X863 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X864 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X865 VSREF single_10b_cdac_0.x10[8].x1.x8.A single_10b_cdac_0.x10[8].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X866 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X867 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X868 VDREF single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X869 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X870 single_10b_cdac_0.x10[8].dac_out single_10b_cdac_0.x10[8].x3.ck a_39174_34963# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X871 VSREF single_10b_cdac_1.x3[1].x1.x5.A single_10b_cdac_1.x3[1].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X872 VDREF SWP_IN[4] a_19338_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X873 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X874 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X875 VDREF single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X876 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X877 a_22558_31002# single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X878 VDREF SWP_IN[3] a_56152_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X879 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x8.A single_10b_cdac_0.cdac_sw_16_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X880 single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X881 a_65951_35702# CF[0] single_10b_cdac_0.x3[0].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X882 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X883 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X884 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X885 VSREF single_10b_cdac_0.x4[2].x1.x3.Y a_59511_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X886 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X887 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X888 single_10b_cdac_0.x3[1].x2.swn single_10b_cdac_0.x3[1].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X889 single_10b_cdac_1.x8[7].x2.swn single_10b_cdac_1.x8[7].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X890 single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.cdac_sw_4_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X891 single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X892 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X893 VSREF single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X894 VSREF single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X895 VCM single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X896 a_24900_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X897 VCM single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X898 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X899 a_30754_25713# single_10b_cdac_1.cdac_sw_1_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[9] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X900 a_53903_24080# single_10b_cdac_0.cdac_sw_2_1.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X901 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X902 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X903 single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.cdac_sw_2_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X904 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X905 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X906 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X907 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X908 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X909 VDREF single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X910 single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X911 single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X912 single_10b_cdac_0.x4[3].x3.ck single_10b_cdac_0.x4[3].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X913 VDREF single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X914 single_10b_cdac_0.cdac_sw_1_1.x2.swn single_10b_cdac_0.cdac_sw_1_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X915 VDREF single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X916 VDREF CF[1] single_10b_cdac_0.x2[0].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X917 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X918 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X919 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X920 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X921 VDREF single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X922 VCM single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X923 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X924 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X925 single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X926 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X927 VSREF single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X928 VDREF single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X929 single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X930 single_10b_cdac_0.x6[5].x2.swn single_10b_cdac_0.x6[5].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X931 VDREF single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X932 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X933 VSREF single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X934 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x9.A single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X935 VDREF single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X936 VDREF SWP_IN[3] a_56152_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X937 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X938 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X939 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X940 VSREF single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X941 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X942 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X943 VDREF single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X944 single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X945 single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X946 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X947 VSREF single_10b_cdac_0.x3[1].x1.x4.A single_10b_cdac_0.x3[1].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X948 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X949 single_10b_cdac_1.x10b_cap_array_0.SW[5] single_10b_cdac_1.cdac_sw_4_0.x3.ckb a_16996_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X950 VSREF single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X951 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x3.ckb a_40930_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X952 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X953 a_25778_31002# single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X954 single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.cdac_sw_8_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X955 single_10b_cdac_0.cdac_sw_2_1.x1.x4.A CF[6] a_53903_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X956 VSREF SWN_IN[9] a_64348_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X957 VDREF single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X958 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X959 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X960 single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X961 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X962 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x8.A single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X963 VSREF single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X964 VDREF single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X965 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X966 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X967 VDREF single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X968 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X969 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X970 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X971 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X972 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X973 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X974 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X975 single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X976 single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X977 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X978 VDREF single_10b_cdac_0.x3[0].x1.x9.A single_10b_cdac_0.x3[0].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X979 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X980 VCN single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X981 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X982 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X983 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X984 single_10b_cdac_1.cdac_sw_1_0.x3.ck single_10b_cdac_1.cdac_sw_1_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X985 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X986 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X987 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X988 single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.cdac_sw_4_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X989 single_10b_cdac_1.x8[6].x2.swn single_10b_cdac_1.x8[6].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X990 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X991 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X992 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X993 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X994 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X995 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X996 VDREF single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X997 single_10b_cdac_0.x6[5].x3.ck single_10b_cdac_0.x6[5].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X998 VSREF single_10b_cdac_1.x6[4].x1.x9.A a_19477_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X999 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1000 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1001 single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1002 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1003 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1004 single_10b_cdac_1.x3[1].x1.x5.A single_10b_cdac_1.x3[1].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1005 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1006 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1007 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1008 single_10b_cdac_1.cdac_sw_2_1.x1.x8.A single_10b_cdac_1.cdac_sw_2_1.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1009 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1010 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1011 VSREF single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1012 single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1013 single_10b_cdac_1.cdac_sw_2_1.x1.x7.A single_10b_cdac_1.cdac_sw_2_1.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1014 single_10b_cdac_0.x3[0].x2.swn single_10b_cdac_0.x3[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1015 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1016 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1017 single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.cdac_sw_16_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1018 VDREF SWP_IN[2] a_59372_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1019 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1020 VSREF single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1021 single_10b_cdac_0.x10b_cap_array_0.SW[9] single_10b_cdac_0.cdac_sw_1_0.x3.ckb a_63470_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1022 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1023 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x9.A single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1024 VSREF single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1025 VSREF single_10b_cdac_1.x8[6].x1.x8.A single_10b_cdac_1.x8[6].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1026 VCM single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1027 VDREF CF[4] single_10b_cdac_0.x6[4].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1028 single_10b_cdac_0.x10b_cap_array_0.SW[4] single_10b_cdac_0.cdac_sw_4_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1029 single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.cdac_sw_4_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1030 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1031 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1032 VCP single_10b_cdac_1.x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1033 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1034 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1035 single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1036 a_20309_24944# single_10b_cdac_1.cdac_sw_2_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1037 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1038 a_44150_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1039 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1040 single_10b_cdac_1.x8[7].x3.ck single_10b_cdac_1.x8[7].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1041 VSREF single_10b_cdac_0.x4[2].x1.x6.A single_10b_cdac_0.x4[2].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1042 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1043 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x8.A single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1044 single_10b_cdac_1.x10b_cap_array_0.SW[7] single_10b_cdac_1.cdac_sw_2_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1045 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1046 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1047 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x9.A single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1048 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1049 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1050 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1051 single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1052 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1053 VSREF single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1054 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1055 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1056 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1057 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1058 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1059 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1060 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1061 single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1062 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1063 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x8.A single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1064 VDREF single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1065 VSREF single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1066 VSREF single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1067 single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1068 VDREF single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1069 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1070 single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1071 VSREF single_10b_cdac_1.x8[6].x1.x5.A single_10b_cdac_1.x8[6].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1072 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1073 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1074 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1075 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1076 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1077 single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1078 VDREF single_10b_cdac_0.x4[2].x1.x9.A single_10b_cdac_0.x4[2].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1079 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1080 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1081 VSREF single_10b_cdac_0.x8[7].x1.x3.Y a_43411_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1082 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1083 single_10b_cdac_1.cdac_sw_1_2.x2.swn single_10b_cdac_1.cdac_sw_1_2.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1084 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1085 single_10b_cdac_0.x3[0].x3.ck single_10b_cdac_0.x3[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1086 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1087 VDREF single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1088 VDREF single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1089 a_25917_35702# CF[2] single_10b_cdac_1.x4[2].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1090 single_10b_cdac_0.cdac_sw_16_0.x1.x8.A single_10b_cdac_0.cdac_sw_16_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1091 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1092 single_10b_cdac_1.x6[4].x2.swn single_10b_cdac_1.x6[4].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1093 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1094 VDREF single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1095 single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1096 a_44150_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1097 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1098 single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.cdac_sw_8_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1099 VDREF single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1100 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1101 single_10b_cdac_0.cdac_sw_1_0.x2.swn single_10b_cdac_0.cdac_sw_1_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1102 single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1103 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1104 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1105 single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1106 VSREF single_10b_cdac_1.x2[0].x1.x8.A single_10b_cdac_1.x2[0].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1107 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1108 single_10b_cdac_1.cdac_sw_1_1.x1.x5.A single_10b_cdac_1.cdac_sw_1_1.x1.x8.A a_26749_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1109 VDREF single_10b_cdac_0.x4[2].x1.x4.A single_10b_cdac_0.x4[2].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1110 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1111 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1112 VSREF single_10b_cdac_1.x3[0].x1.x8.A single_10b_cdac_1.x3[0].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1113 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1114 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1115 VDREF single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1116 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1117 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1118 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1119 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1120 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1121 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1122 single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1123 VDREF single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1124 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1125 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1126 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1127 single_10b_cdac_0.x10b_cap_array_0.SW[5] single_10b_cdac_0.cdac_sw_4_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1128 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x9.A single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1129 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1130 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1131 VDREF single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1132 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1133 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1134 VSREF single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1135 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1136 VCN single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1137 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1138 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1139 single_10b_cdac_1.x4[2].x2.swn single_10b_cdac_1.x4[2].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1140 single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1141 VSREF single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1142 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x8.A single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1143 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1144 VDREF single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1145 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1146 single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1147 single_10b_cdac_1.x8[7].dac_out single_10b_cdac_1.x8[7].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1148 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1149 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1150 single_10b_cdac_1.cdac_sw_1_2.x1.x4.A CF[9] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1151 a_58494_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1152 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1153 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1154 single_10b_cdac_0.cdac_sw_4_1.x1.x3.Y CF[4] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1155 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x5.A single_10b_cdac_1.cdac_sw_1_2.x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1156 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1157 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1158 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x3.ck a_58494_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1159 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1160 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1161 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1162 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1163 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1164 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1165 VDREF single_10b_cdac_1.x10[8].x1.x3.Y single_10b_cdac_1.x10[8].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1166 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1167 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1168 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1169 single_10b_cdac_1.cdac_sw_1_1.x3.ck single_10b_cdac_1.cdac_sw_1_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1170 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1171 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1172 single_10b_cdac_1.x2[0].x1.x9.A single_10b_cdac_1.x2[0].x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1173 single_10b_cdac_1.x6[4].dac_out single_10b_cdac_1.x6[4].x3.ck a_18460_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1174 single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1175 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1176 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1177 single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1178 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1179 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1180 single_10b_cdac_0.x4[2].x3.ck single_10b_cdac_0.x4[2].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1181 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1182 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1183 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1184 VCN single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1185 single_10b_cdac_1.cdac_sw_16_0.x1.x3.Y CF[0] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1186 single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1187 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1188 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1189 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x8.A single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1190 VDREF single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1191 single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1192 single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.cdac_sw_2_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1193 single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1194 single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1195 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1196 VDREF single_10b_cdac_1.x10[8].x1.x7.A single_10b_cdac_1.x10[8].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1197 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1198 single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1199 a_4209_24080# single_10b_cdac_1.x2[0].x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1200 single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1201 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1202 VCM single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1203 single_10b_cdac_1.x8[6].x1.x5.A single_10b_cdac_1.x8[6].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1204 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1205 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1206 VDREF single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1207 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1208 single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1209 single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1210 VDREF single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1211 single_10b_cdac_0.cdac_sw_1_0.x1.x7.A single_10b_cdac_0.cdac_sw_1_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1212 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1213 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1214 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1215 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1216 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1217 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1218 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1219 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1220 VDREF SWP_IN[7] a_9678_34218# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1221 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1222 single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1223 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1224 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x3.ckb a_10556_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1225 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1226 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1227 VSREF single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1228 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1229 single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1230 single_10b_cdac_1.x3[1].x2.swn single_10b_cdac_1.x3[1].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1231 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1232 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1233 VDREF single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1234 single_10b_cdac_0.x8[6].x1.x4.A CF[6] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1235 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1236 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1237 VSREF single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1238 single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1239 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1240 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1241 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1242 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1243 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1244 VSREF single_10b_cdac_0.x8[7].x1.x6.A single_10b_cdac_0.x8[7].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1245 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1246 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1247 single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1248 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1249 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1250 single_10b_cdac_0.cdac_sw_1_0.x3.ck single_10b_cdac_0.cdac_sw_1_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1251 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1252 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1253 VDREF single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1254 single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1255 VSREF single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1256 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1257 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1258 a_16118_33146# single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1259 single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.cdac_sw_2_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1260 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1261 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1262 VDREF single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1263 VDREF single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1264 single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1265 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1266 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1267 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1268 a_40930_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1269 single_10b_cdac_1.x10[8].x3.ck single_10b_cdac_1.x10[8].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1270 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1271 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1272 VSREF single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1273 VSREF SWN_IN[2] a_8214_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1274 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1275 single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1276 VDREF single_10b_cdac_0.x8[7].x1.x9.A single_10b_cdac_0.x8[7].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1277 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1278 single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1279 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1280 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1281 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1282 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x9.A single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1283 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1284 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1285 a_24314_25713# single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[7] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1286 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1287 a_47463_24080# single_10b_cdac_0.cdac_sw_4_1.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1288 single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1289 a_16996_25722# SWN_IN[5] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1290 single_10b_cdac_0.cdac_sw_1_1.x1.x5.A single_10b_cdac_0.cdac_sw_1_1.x1.x8.A a_60343_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1291 VDREF single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1292 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1293 single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1294 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1295 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1296 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1297 VDREF single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1298 a_8800_34645# SWP_IN[7] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1299 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1300 single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1301 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1302 single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.cdac_sw_2_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1303 VCM single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1304 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1305 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1306 VDREF single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1307 single_10b_cdac_1.cdac_sw_8_0.x1.x5.A single_10b_cdac_1.cdac_sw_8_0.x1.x8.A a_10649_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1308 VDREF single_10b_cdac_0.x8[7].x1.x4.A single_10b_cdac_0.x8[7].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1309 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1310 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1311 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1312 single_10b_cdac_0.x3[1].x3.ck single_10b_cdac_0.x3[1].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1313 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1314 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1315 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1316 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1317 single_10b_cdac_0.cdac_sw_1_2.x3.ck single_10b_cdac_0.cdac_sw_1_2.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1318 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1319 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1320 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1321 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1322 VCM single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[7] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1323 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1324 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1325 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1326 VDREF single_10b_cdac_1.x10[8].x1.x9.A single_10b_cdac_1.x10[8].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1327 single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1328 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1329 VDREF single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1330 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1331 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1332 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x9.A single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1333 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1334 VSREF SWN_IN[2] a_41808_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1335 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1336 single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1337 VSREF single_10b_cdac_0.x4[3].x1.x4.A single_10b_cdac_0.x4[3].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1338 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1339 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1340 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1341 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1342 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1343 single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.cdac_sw_2_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1344 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1345 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1346 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1347 a_19338_33146# single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1348 a_51468_25713# single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1349 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1350 a_23436_25722# SWN_IN[7] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1351 single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.cdac_sw_16_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1352 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1353 single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1354 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1355 VSREF single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1356 single_10b_cdac_0.cdac_sw_4_1.x1.x4.A CF[4] a_47463_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1357 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1358 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1359 single_10b_cdac_0.cdac_sw_1_1.x2.swn single_10b_cdac_0.cdac_sw_1_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1360 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1361 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1362 VSREF single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1363 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x8.A single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1364 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1365 a_21680_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1366 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1367 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1368 VCM single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1369 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1370 VDREF single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1371 VSREF single_10b_cdac_0.x8[6].x1.x9.A single_10b_cdac_0.x8[6].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1372 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1373 single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.cdac_sw_8_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1374 single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1375 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1376 VDREF single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1377 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1378 a_7336_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1379 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1380 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1381 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1382 single_10b_cdac_0.x8[7].x3.ck single_10b_cdac_0.x8[7].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1383 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1384 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1385 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1386 single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1387 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1388 single_10b_cdac_0.cdac_sw_1_0.x3.ck single_10b_cdac_0.cdac_sw_1_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1389 VCM single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1390 single_10b_cdac_1.cdac_sw_8_1.x1.x4.A CF[2] a_7429_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1391 single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.cdac_sw_4_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1392 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1393 single_10b_cdac_1.x6[4].x3.ck single_10b_cdac_1.x6[4].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1394 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1395 single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.cdac_sw_8_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1396 single_10b_cdac_1.cdac_sw_4_1.x1.x8.A single_10b_cdac_1.cdac_sw_4_1.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1397 VSREF single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1398 single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1399 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1400 single_10b_cdac_1.cdac_sw_4_1.x1.x7.A single_10b_cdac_1.cdac_sw_4_1.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1401 VDREF single_10b_cdac_0.x10[8].x1.x6.A single_10b_cdac_0.x10[8].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1402 single_10b_cdac_0.x4[2].x2.swn single_10b_cdac_0.x4[2].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1403 VSREF single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1404 single_10b_cdac_0.x4[3].x3.ck single_10b_cdac_0.x4[3].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1405 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1406 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1407 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1408 single_10b_cdac_0.x10b_cap_array_0.SW[7] single_10b_cdac_0.cdac_sw_2_0.x3.ckb a_57030_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1409 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1410 VSREF single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1411 single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1412 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1413 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1414 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1415 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1416 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1417 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1418 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1419 VDREF single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1420 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1421 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1422 single_10b_cdac_1.x3[0].x3.ck single_10b_cdac_1.x3[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1423 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1424 single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1425 single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1426 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x3.ck a_55274_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1427 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1428 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1429 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1430 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1431 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1432 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1433 VDREF single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1434 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1435 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1436 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1437 single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1438 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1439 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1440 single_10b_cdac_1.x8[6].x2.swn single_10b_cdac_1.x8[6].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1441 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1442 VDREF single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1443 single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1444 single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.cdac_sw_16_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1445 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1446 VSREF single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1447 single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1448 single_10b_cdac_1.x10b_cap_array_0.SW[4] single_10b_cdac_1.cdac_sw_4_1.x3.ckb a_13776_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1449 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1450 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1451 single_10b_cdac_1.cdac_sw_4_0.x1.x6.A single_10b_cdac_1.cdac_sw_4_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1452 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1453 single_10b_cdac_0.x10b_cap_array_0.SW[7] single_10b_cdac_0.cdac_sw_2_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1454 single_10b_cdac_0.cdac_sw_4_0.x1.x3.Y CF[5] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1455 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1456 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1457 single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1458 VSREF single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1459 single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.cdac_sw_4_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1460 single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1461 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1462 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1463 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1464 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1465 single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.cdac_sw_16_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1466 VDREF single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1467 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1468 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1469 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1470 VDREF single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1471 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1472 VSREF CF[1] single_10b_cdac_0.x3[1].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1473 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1474 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1475 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x9.A single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1476 single_10b_cdac_1.cdac_sw_1_1.x3.ck single_10b_cdac_1.cdac_sw_1_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1477 a_59372_31002# single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1478 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1479 single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1480 single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1481 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1482 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1483 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1484 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1485 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x3.Y a_36971_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1486 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1487 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1488 single_10b_cdac_0.x4[2].x3.ck single_10b_cdac_0.x4[2].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1489 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1490 VCM single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1491 VDREF single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1492 VSREF single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1493 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1494 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1495 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1496 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1497 single_10b_cdac_1.x8[7].x3.ck single_10b_cdac_1.x8[7].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1498 single_10b_cdac_1.x6[5].x3.ck single_10b_cdac_1.x6[5].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1499 a_19477_35702# CF[4] single_10b_cdac_1.x6[4].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1500 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1501 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1502 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1503 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1504 single_10b_cdac_0.x2[0].x1.x5.A single_10b_cdac_0.x2[0].x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1505 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1506 single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1507 a_11434_25713# single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1508 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1509 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1510 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1511 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x8.A single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1512 single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1513 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1514 VDREF single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1515 single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1516 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1517 VSREF single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1518 single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x2[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1519 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1520 VDREF SWP_IN[3] a_22558_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1521 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1522 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1523 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1524 VSREF single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1525 VSREF single_10b_cdac_1.x4[2].x1.x3.Y a_25917_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1526 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1527 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1528 VDREF single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1529 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1530 single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1531 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1532 single_10b_cdac_0.x2[0].x1.x7.A single_10b_cdac_0.x2[0].x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1533 VDREF single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1534 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1535 VDREF single_10b_cdac_0.x3[1].x1.x8.A single_10b_cdac_0.x3[1].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1536 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1537 VSREF single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1538 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1539 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1540 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1541 single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1542 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1543 VDREF single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1544 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1545 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1546 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1547 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1548 single_10b_cdac_1.x4[3].x3.ck single_10b_cdac_1.x4[3].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1549 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1550 single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1551 VSREF single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1552 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1553 single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.cdac_sw_8_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1554 single_10b_cdac_1.x4[3].x3.ck single_10b_cdac_1.x4[3].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1555 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1556 VSREF single_10b_cdac_1.x4[2].x1.x7.A single_10b_cdac_1.x4[2].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1557 single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.cdac_sw_16_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1558 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1559 VSREF SWN_IN[3] a_45028_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1560 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1561 VCN single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1562 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1563 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1564 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1565 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1566 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1567 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1568 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1569 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1570 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1571 single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1572 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1573 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1574 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x8.A single_10b_cdac_1.cdac_sw_1_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1575 VCM single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1576 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1577 VSREF single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1578 VDREF SWP_IN[3] a_22558_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1579 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1580 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1581 single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1582 VDREF single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1583 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1584 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1585 single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1586 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1587 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1588 VSREF single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1589 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1590 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1591 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1592 VCM single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1593 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1594 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1595 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1596 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1597 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1598 VDREF single_10b_cdac_1.x4[3].x1.x9.A single_10b_cdac_1.x4[3].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1599 single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x2[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1600 VSREF single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1601 single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1602 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1603 VDREF single_10b_cdac_1.x3[1].x1.x7.A single_10b_cdac_1.x3[1].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1604 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1605 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1606 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1607 single_10b_cdac_1.cdac_sw_2_0.x1.x3.Y CF[7] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1608 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1609 a_26749_24080# single_10b_cdac_1.cdac_sw_1_1.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1610 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1611 single_10b_cdac_0.x10b_cap_array_0.SW[6] single_10b_cdac_0.cdac_sw_2_1.x3.ckb a_53810_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1612 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1613 VDREF single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1614 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1615 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1616 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1617 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1618 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1619 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1620 single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1621 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1622 single_10b_cdac_0.cdac_sw_2_0.x1.x7.A single_10b_cdac_0.cdac_sw_2_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1623 single_10b_cdac_0.x8[7].x2.swn single_10b_cdac_0.x8[7].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1624 single_10b_cdac_1.x6[5].dac_out single_10b_cdac_1.x6[5].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1625 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1626 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1627 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1628 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x3.ckb a_40930_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1629 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1630 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1631 VDREF single_10b_cdac_1.x4[3].x1.x4.A single_10b_cdac_1.x4[3].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1632 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1633 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1634 VSREF single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1635 single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1636 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1637 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1638 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1639 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1640 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1641 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1642 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1643 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1644 single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1645 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1646 single_10b_cdac_1.x6[5].x3.ck single_10b_cdac_1.x6[5].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1647 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1648 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1649 single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.cdac_sw_8_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1650 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1651 VDREF single_10b_cdac_0.x6[4].x1.x9.A single_10b_cdac_0.x6[4].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1652 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1653 single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1654 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1655 single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.cdac_sw_16_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1656 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1657 single_10b_cdac_1.x6[5].x3.ck single_10b_cdac_1.x6[5].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1658 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x6.A single_10b_cdac_0.cdac_sw_1_2.x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1659 single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1660 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1661 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1662 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1663 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1664 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1665 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1666 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1667 single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1668 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1669 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1670 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1671 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1672 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1673 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1674 single_10b_cdac_1.x10[8].x1.x5.A single_10b_cdac_1.x10[8].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1675 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1676 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1677 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1678 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1679 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1680 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1681 VSREF single_10b_cdac_0.x3[0].x1.x9.A a_65951_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1682 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1683 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1684 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1685 VDREF single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1686 single_10b_cdac_1.x10b_cap_array_0.SW[4] single_10b_cdac_1.cdac_sw_4_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1687 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1688 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1689 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1690 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1691 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x3.ck a_21680_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1692 VCP single_10b_cdac_0.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1693 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1694 single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1695 single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1696 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1697 VCM single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1698 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1699 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x9.A single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1700 single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1701 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x3.ckb a_40930_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1702 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1703 single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1704 single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1705 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1706 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1707 single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1708 VSREF single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1709 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1710 single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.cdac_sw_4_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1711 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1712 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1713 a_57908_25713# single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[7] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1714 single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1715 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1716 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1717 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1718 VSREF single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1719 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1720 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1721 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1722 VDREF single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1723 a_10556_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1724 single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1725 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1726 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x8.A single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1727 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1728 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1729 single_10b_cdac_0.cdac_sw_1_2.x2.swn single_10b_cdac_0.cdac_sw_1_2.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1730 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1731 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1732 single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1733 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1734 single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1735 a_9678_34218# single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1736 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1737 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1738 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1739 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1740 single_10b_cdac_0.cdac_sw_4_0.x1.x9.A single_10b_cdac_0.cdac_sw_4_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1741 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1742 VCM single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1743 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1744 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1745 single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1746 VSREF single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1747 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1748 VSREF single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1749 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1750 VSREF single_10b_cdac_0.x6[4].x1.x9.A single_10b_cdac_0.x6[4].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1751 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1752 single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1753 VDREF single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1754 single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1755 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1756 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x9.A single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1757 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1758 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1759 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1760 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1761 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1762 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1763 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1764 VSREF single_10b_cdac_1.x3[1].x1.x9.A single_10b_cdac_1.x3[1].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1765 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1766 VDREF single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1767 single_10b_cdac_0.x10b_cap_array_0.SW[8] single_10b_cdac_0.cdac_sw_1_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1768 single_10b_cdac_0.x6[5].x1.x5.A single_10b_cdac_0.x6[5].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1769 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1770 VDREF single_10b_cdac_0.x3[1].x1.x3.Y single_10b_cdac_0.x3[1].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1771 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x6.A single_10b_cdac_1.cdac_sw_1_2.x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1772 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1773 single_10b_cdac_1.cdac_sw_1_0.x2.swn single_10b_cdac_1.cdac_sw_1_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1774 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1775 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1776 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1777 single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.cdac_sw_2_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1778 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1779 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1780 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1781 single_10b_cdac_0.x6[4].x2.swn single_10b_cdac_0.x6[4].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1782 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x3.ck a_24900_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1783 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1784 single_10b_cdac_0.cdac_sw_2_1.x1.x8.A single_10b_cdac_0.cdac_sw_2_1.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1785 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1786 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1787 VSREF single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1788 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1789 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1790 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1791 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1792 a_15240_34009# SWP_IN[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1793 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1794 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1795 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1796 VDREF single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1797 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1798 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x3.ckb a_44150_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1799 VSREF single_10b_cdac_0.x10[8].x1.x9.A single_10b_cdac_0.x10[8].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1800 single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1801 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1802 single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1803 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x9.A single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1804 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1805 VDREF single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1806 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x9.A single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1807 VDREF single_10b_cdac_0.x3[1].x1.x7.A single_10b_cdac_0.x3[1].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1808 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1809 a_41023_24944# single_10b_cdac_0.cdac_sw_8_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1810 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1811 VCM single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1812 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1813 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1814 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1815 VCM single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1816 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1817 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1818 a_65951_36566# single_10b_cdac_0.x3[0].x1.x8.A single_10b_cdac_0.x3[0].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1819 a_13776_25722# SWN_IN[4] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1820 VSREF single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1821 single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.cdac_sw_2_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1822 VCM single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1823 single_10b_cdac_0.x6[4].x2.swn single_10b_cdac_0.x6[4].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1824 VDREF SWP_IN[2] a_25778_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1825 VDREF single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1826 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1827 single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1828 VSREF single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1829 VDREF single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1830 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1831 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1832 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1833 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1834 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1835 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1836 VDREF single_10b_cdac_1.x8[6].x1.x7.A single_10b_cdac_1.x8[6].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1837 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1838 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1839 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1840 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1841 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1842 a_10649_24080# single_10b_cdac_1.cdac_sw_8_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1843 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1844 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1845 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1846 VSREF single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1847 VSREF single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1848 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1849 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1850 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1851 single_10b_cdac_0.cdac_sw_4_1.x1.x7.A single_10b_cdac_0.cdac_sw_4_1.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1852 VDREF single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1853 single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1854 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1855 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x9.A single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1856 VDREF single_10b_cdac_0.x8[6].x1.x5.A single_10b_cdac_0.x8[6].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1857 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1858 single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1859 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1860 single_10b_cdac_0.cdac_sw_8_1.x1.x7.A single_10b_cdac_0.cdac_sw_8_1.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1861 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1862 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1863 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1864 VDREF single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1865 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1866 single_10b_cdac_0.x6[5].dac_out single_10b_cdac_0.x6[5].x3.ck a_48834_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1867 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1868 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1869 a_46492_34218# single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1870 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1871 single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1872 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1873 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1874 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x8.A single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1875 single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.cdac_sw_2_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1876 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1877 VSREF single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1878 VSREF single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1879 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1880 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1881 VDREF single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1882 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1883 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1884 VSREF single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1885 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1886 single_10b_cdac_1.cdac_sw_8_1.x1.x8.A single_10b_cdac_1.cdac_sw_8_1.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1887 single_10b_cdac_0.x3[1].x3.ck single_10b_cdac_0.x3[1].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1888 single_10b_cdac_0.x10b_cap_array_0.SW[4] single_10b_cdac_0.cdac_sw_4_1.x3.ckb a_47370_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1889 VSREF single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1890 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1891 single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1892 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1893 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1894 single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1895 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1896 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1897 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x3.ck a_58494_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1898 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1899 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1900 single_10b_cdac_1.cdac_sw_16_0.x1.x7.A single_10b_cdac_1.cdac_sw_16_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1901 single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1902 VSREF single_10b_cdac_0.x3[1].x1.x5.A single_10b_cdac_0.x3[1].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1903 VDREF CF[1] single_10b_cdac_1.x3[1].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1904 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1905 single_10b_cdac_0.cdac_sw_1_2.x3.ck single_10b_cdac_0.cdac_sw_1_2.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1906 VSREF single_10b_cdac_0.x6[5].x1.x8.A single_10b_cdac_0.x6[5].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1907 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1908 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1909 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1910 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1911 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1912 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1913 VCM single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1914 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1915 single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1916 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1917 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1918 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1919 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1920 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1921 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1922 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1923 single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1924 a_7429_24944# single_10b_cdac_1.cdac_sw_8_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1925 single_10b_cdac_0.x8[6].x2.swn single_10b_cdac_0.x8[6].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1926 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1927 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1928 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x8.A single_10b_cdac_0.cdac_sw_8_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1929 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1930 single_10b_cdac_1.cdac_sw_1_1.x1.x6.A single_10b_cdac_1.cdac_sw_1_1.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1931 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1932 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1933 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1934 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1935 VSREF single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1936 single_10b_cdac_0.x6[5].x3.ck single_10b_cdac_0.x6[5].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1937 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1938 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1939 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1940 a_41808_25713# single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1941 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1942 a_45028_25713# single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1943 single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1944 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1945 VDREF single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1946 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1947 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1948 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1949 single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1950 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1951 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1952 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1953 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1954 VSREF single_10b_cdac_1.x6[4].x1.x3.Y a_19477_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1955 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1956 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1957 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1958 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1959 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1960 VSREF single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1961 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1962 VDREF single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1963 VDREF single_10b_cdac_0.x4[3].x1.x8.A single_10b_cdac_0.x4[3].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1964 VSREF single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1965 VSREF single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1966 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1967 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1968 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1969 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1970 VDREF single_10b_cdac_1.x10[8].x1.x8.A single_10b_cdac_1.x10[8].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1971 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1972 VSREF single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1973 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1974 single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1975 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1976 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1977 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1978 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1979 single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1980 single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.cdac_sw_16_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1981 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1982 VSREF single_10b_cdac_1.x8[6].x1.x9.A single_10b_cdac_1.x8[6].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1983 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1984 single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1985 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1986 single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.cdac_sw_2_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1987 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1988 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1989 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1990 VDREF single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1991 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1992 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1993 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1994 single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1995 VSREF single_10b_cdac_0.x4[2].x1.x7.A single_10b_cdac_0.x4[2].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1996 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1997 single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1998 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1999 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2000 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2001 VSREF single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2002 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2003 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2004 VDREF SWP_IN[5] a_16118_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2005 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2006 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2007 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x8.A single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2008 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2009 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2010 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2011 single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2012 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2013 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2014 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x8.A single_10b_cdac_0.cdac_sw_1_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2015 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2016 VSREF single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2017 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2018 single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2019 VSREF single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2020 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2021 single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.cdac_sw_2_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2022 a_22558_31002# single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2023 VDREF single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2024 VDREF single_10b_cdac_1.x6[5].x1.x9.A single_10b_cdac_1.x6[5].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2025 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2026 single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.cdac_sw_4_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2027 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2028 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2029 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2030 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2031 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2032 single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.cdac_sw_8_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2033 single_10b_cdac_1.cdac_sw_4_1.x1.x4.A CF[4] a_13869_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2034 VSREF SWN_IN[7] a_24314_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2035 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2036 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2037 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2038 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2039 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2040 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2041 single_10b_cdac_0.cdac_sw_2_0.x1.x3.Y CF[7] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2042 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2043 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2044 a_25917_36566# single_10b_cdac_1.x4[2].x1.x8.A single_10b_cdac_1.x4[2].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2045 a_8214_25713# single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2046 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2047 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2048 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2049 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2050 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2051 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2052 VSREF single_10b_cdac_1.x3[1].x1.x9.A a_29137_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2053 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2054 single_10b_cdac_0.x4[2].x3.ck single_10b_cdac_0.x4[2].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2055 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2056 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x8.A single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2057 VDREF single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2058 VDREF single_10b_cdac_0.x6[5].x1.x8.A single_10b_cdac_0.x6[5].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2059 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2060 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2061 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2062 VSREF single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2063 single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2064 single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2065 single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2066 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2067 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2068 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2069 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2070 single_10b_cdac_1.cdac_sw_1_0.x1.x9.A single_10b_cdac_1.cdac_sw_1_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2071 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2072 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2073 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2074 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2075 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2076 VSREF single_10b_cdac_1.x3[0].x1.x9.A single_10b_cdac_1.x3[0].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2077 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2078 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2079 VSREF single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2080 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2081 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2082 VDREF single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2083 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2084 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2085 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2086 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2087 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2088 VDREF single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2089 VCM single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2090 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2091 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2092 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2093 single_10b_cdac_1.x6[4].dac_out single_10b_cdac_1.x6[4].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2094 single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2095 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2096 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2097 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2098 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2099 VDREF SWP_IN[3] a_56152_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2100 single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2101 single_10b_cdac_1.x4[2].x2.swn single_10b_cdac_1.x4[2].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2102 a_55274_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2103 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2104 VDREF SWP_IN[4] a_19338_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2105 single_10b_cdac_1.x10b_cap_array_0.SW[7] single_10b_cdac_1.cdac_sw_2_0.x3.ckb a_23436_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2106 VSREF SWN_IN[5] a_51468_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2107 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2108 single_10b_cdac_0.cdac_sw_16_0.x1.x6.A single_10b_cdac_0.cdac_sw_16_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2109 VSREF single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2110 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x8.A single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2111 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2112 single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.cdac_sw_8_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2113 single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2114 single_10b_cdac_0.x6[4].dac_out single_10b_cdac_0.x6[4].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2115 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2116 VDREF CF[6] single_10b_cdac_1.x8[6].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2117 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2118 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2119 single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2120 single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2122 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2123 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2124 VDREF single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2125 single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2126 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2127 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2128 VSREF single_10b_cdac_1.x6[4].x1.x6.A single_10b_cdac_1.x6[4].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2129 single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.cdac_sw_8_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2130 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x3.ckb a_7336_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2131 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2132 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2133 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2134 VDREF single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2135 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2136 VCP single_10b_cdac_1.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2137 VCP single_10b_cdac_1.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2138 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2139 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2140 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2141 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2142 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2143 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2144 single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2145 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2146 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2147 VCM single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2148 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2149 single_10b_cdac_0.cdac_sw_4_0.x1.x6.A single_10b_cdac_0.cdac_sw_4_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2150 single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2151 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2152 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2153 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2154 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2155 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2156 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2157 single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2158 single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2159 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2160 single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.cdac_sw_4_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2161 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2162 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2163 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2164 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2165 single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2166 VSREF single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2167 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2168 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2169 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2170 single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2171 single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x2[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2172 VDREF single_10b_cdac_1.x4[2].x1.x5.A single_10b_cdac_1.x4[2].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2173 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2174 VSREF single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2175 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2176 VDREF single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2177 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2178 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2179 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2180 single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2181 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2182 a_25778_31002# single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2183 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2184 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2185 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2186 VDREF single_10b_cdac_0.x4[3].x1.x3.Y single_10b_cdac_0.x4[3].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2187 VCP single_10b_cdac_0.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2188 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2189 single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2190 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2191 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2192 single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2193 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2194 VSREF single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2195 VDREF single_10b_cdac_1.x6[5].x1.x8.A single_10b_cdac_1.x6[5].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2196 single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2197 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2198 single_10b_cdac_0.cdac_sw_4_1.x1.x8.A single_10b_cdac_0.cdac_sw_4_1.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2199 single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2200 single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2201 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2202 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2203 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2204 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2205 VSREF single_10b_cdac_0.x8[7].x1.x7.A single_10b_cdac_0.x8[7].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2206 single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2207 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2208 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x8.A single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2209 a_48834_34009# SWP_IN[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2210 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2211 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2212 single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.cdac_sw_8_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2213 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2214 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2215 single_10b_cdac_0.x6[4].dac_out single_10b_cdac_0.x6[4].x3.ck a_52054_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2216 VSREF SWN_IN[5] a_17874_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2217 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2218 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2219 VDREF single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2220 single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x2[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2221 a_34583_24944# single_10b_cdac_0.cdac_sw_16_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2222 VSREF single_10b_cdac_1.x3[1].x1.x8.A single_10b_cdac_1.x3[1].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2223 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2224 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2225 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2226 VSREF single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2227 VSREF single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2228 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2229 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2230 single_10b_cdac_0.x8[6].x2.swn single_10b_cdac_0.x8[6].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2231 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2232 single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2233 single_10b_cdac_1.x10[8].x2.swn single_10b_cdac_1.x10[8].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2234 a_18460_34009# SWP_IN[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2235 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2236 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2237 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2238 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2239 single_10b_cdac_0.cdac_sw_1_0.x1.x8.A single_10b_cdac_0.cdac_sw_1_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2240 VDREF SWP_IN[2] a_59372_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2241 single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2242 VSREF SWN_IN[3] a_11434_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2243 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2244 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2245 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2246 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2247 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2248 VSREF single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2249 a_52932_33146# single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2250 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2251 single_10b_cdac_0.cdac_sw_8_1.x1.x3.Y CF[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2252 single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2253 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x9.A single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2254 VDREF single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2255 VCM single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2256 single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2257 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2258 VDREF single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2259 VCM single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2260 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2261 VDREF CF[5] single_10b_cdac_0.cdac_sw_4_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2262 VSREF single_10b_cdac_1.x8[6].x1.x9.A a_13037_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2263 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2264 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2265 single_10b_cdac_0.x8[7].x3.ck single_10b_cdac_0.x8[7].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2266 VDREF single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2267 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2268 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2269 single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2270 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2271 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2272 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2273 VCM single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2274 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2275 single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2276 VDREF single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2277 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2278 VSREF single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2279 single_10b_cdac_0.x3[1].x2.swn single_10b_cdac_0.x3[1].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2280 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2281 VSREF single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2282 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2283 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2284 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2285 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2286 single_10b_cdac_0.cdac_sw_1_2.x2.swn single_10b_cdac_0.cdac_sw_1_2.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2287 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2288 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2289 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2290 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2291 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2292 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2293 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2294 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2295 VDREF single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2296 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2297 single_10b_cdac_0.x4[3].x1.x4.A CF[3] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2298 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2299 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2300 single_10b_cdac_1.cdac_sw_2_0.x1.x7.A single_10b_cdac_1.cdac_sw_2_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2301 single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2302 VSREF single_10b_cdac_0.x4[3].x1.x5.A single_10b_cdac_0.x4[3].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2303 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2304 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2305 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2306 single_10b_cdac_0.cdac_sw_1_1.x2.swn single_10b_cdac_0.cdac_sw_1_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2307 single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2308 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2309 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2310 single_10b_cdac_0.cdac_sw_2_0.x1.x9.A single_10b_cdac_0.cdac_sw_2_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2311 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2312 single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2313 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2314 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2315 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2316 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2317 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2318 VDREF single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2319 VSREF single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2320 VSREF single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2321 VDREF single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2322 a_29969_24944# single_10b_cdac_1.cdac_sw_1_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2323 single_10b_cdac_1.cdac_sw_1_0.x2.swn single_10b_cdac_1.cdac_sw_1_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2324 single_10b_cdac_0.x10[8].x2.swn single_10b_cdac_0.x10[8].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2325 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2326 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2327 VDREF single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2328 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2329 single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2330 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2331 VSREF single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2332 a_50590_25722# SWN_IN[5] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2333 VDREF single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2334 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2335 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2336 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2337 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2338 single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2339 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2340 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2341 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2342 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2343 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2344 a_57123_24080# single_10b_cdac_0.cdac_sw_2_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2345 single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2346 VDREF single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2347 VSREF single_10b_cdac_1.x3[0].x1.x9.A a_32357_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2348 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2349 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2350 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2351 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2352 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2353 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2354 VSREF single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2355 single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2356 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2357 single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2358 single_10b_cdac_0.x10b_cap_array_0.SW[5] single_10b_cdac_0.cdac_sw_4_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2359 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2360 VDREF single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2361 VSREF single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2362 single_10b_cdac_0.x4[3].x2.swn single_10b_cdac_0.x4[3].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2363 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2364 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2365 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2366 VSREF single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2367 single_10b_cdac_1.cdac_sw_2_1.x1.x5.A single_10b_cdac_1.cdac_sw_2_1.x1.x8.A a_20309_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2368 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2369 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2370 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2371 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2372 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2373 single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2374 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2375 single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2376 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2377 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2378 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2379 single_10b_cdac_1.cdac_sw_1_0.x3.ck single_10b_cdac_1.cdac_sw_1_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2380 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2381 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2382 single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.cdac_sw_4_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2383 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2384 single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.cdac_sw_4_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2385 single_10b_cdac_1.x3[0].x2.swn single_10b_cdac_1.x3[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2386 VDREF single_10b_cdac_0.x10[8].x1.x3.Y single_10b_cdac_0.x10[8].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2387 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2388 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2389 single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2390 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2391 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2392 single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2393 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2394 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2395 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2396 single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2397 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2398 VCP single_10b_cdac_0.x3[0].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2399 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2400 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2401 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x8.A single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2402 single_10b_cdac_0.cdac_sw_2_0.x1.x4.A CF[7] a_57123_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2403 VDREF single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2404 single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2405 VSREF single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2406 single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2407 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2408 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x9.A single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2409 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x3.ck a_21680_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2410 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2411 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2412 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2413 VSREF single_10b_cdac_1.x8[6].x1.x8.A single_10b_cdac_1.x8[6].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2414 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2415 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2416 single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.cdac_sw_4_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2417 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2418 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2419 single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2420 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2421 VDREF single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2422 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2423 single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2424 a_11434_25713# single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2425 VSREF single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2426 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2427 single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.cdac_sw_2_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2428 single_10b_cdac_1.x8[7].x3.ck single_10b_cdac_1.x8[7].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2429 single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2430 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2431 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2432 single_10b_cdac_0.x6[4].x3.ck single_10b_cdac_0.x6[4].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2433 VDREF single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2434 VDREF SWP_IN[7] a_43272_34218# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2435 single_10b_cdac_1.x6[5].x2.swn single_10b_cdac_1.x6[5].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2436 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2437 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2438 a_19477_36566# single_10b_cdac_1.x6[4].x1.x8.A single_10b_cdac_1.x6[4].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2439 single_10b_cdac_1.x3[0].x2.swn single_10b_cdac_1.x3[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2440 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x3.ckb a_10556_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2441 VCP single_10b_cdac_1.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2442 VCP single_10b_cdac_1.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2443 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2444 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2445 single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2446 single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2447 single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2448 VDREF SWP_IN[7] a_9678_34218# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2449 single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2450 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2451 single_10b_cdac_1.cdac_sw_2_0.x1.x8.A single_10b_cdac_1.cdac_sw_2_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2452 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2453 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2454 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2455 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2456 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2457 single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2458 VDREF single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2459 single_10b_cdac_0.x3[0].x3.ck single_10b_cdac_0.x3[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2460 VDREF single_10b_cdac_0.x4[2].x1.x9.A single_10b_cdac_0.x4[2].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2461 VSREF single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2462 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2463 single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.cdac_sw_2_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2464 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2465 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2466 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2467 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2468 single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2469 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2470 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2471 VDREF single_10b_cdac_1.x8[7].x1.x9.A single_10b_cdac_1.x8[7].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2472 a_56152_31002# single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2473 VDREF single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2474 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2475 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2476 single_10b_cdac_0.x10[8].x3.ck single_10b_cdac_0.x10[8].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2477 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2478 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2479 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2480 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2481 single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2482 single_10b_cdac_1.cdac_sw_16_0.x1.x4.A single_10b_cdac_1.cdac_sw_16_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2483 single_10b_cdac_1.x6[4].x2.swn single_10b_cdac_1.x6[4].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2484 VDREF single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2485 VSREF SWN_IN[3] a_45028_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2486 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2487 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2488 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x8.A single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2489 single_10b_cdac_1.x4[3].x2.swn single_10b_cdac_1.x4[3].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2490 single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2491 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2492 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2493 VSREF single_10b_cdac_1.x2[0].x1.x8.A single_10b_cdac_1.x2[0].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2494 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2495 single_10b_cdac_0.x8[6].dac_out single_10b_cdac_0.x8[6].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2496 single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2497 VSREF single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2498 single_10b_cdac_0.x10[8].x1.x4.A CF[8] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2499 single_10b_cdac_1.cdac_sw_1_1.x1.x8.A single_10b_cdac_1.cdac_sw_1_1.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2500 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2501 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2502 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2503 single_10b_cdac_0.cdac_sw_1_1.x1.x3.Y CF[8] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2504 VDREF single_10b_cdac_1.x8[7].x1.x4.A single_10b_cdac_1.x8[7].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2505 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2506 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2507 VDREF CF[6] single_10b_cdac_0.x8[6].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2508 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2509 VDREF single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2510 single_10b_cdac_0.cdac_sw_8_1.x1.x9.A single_10b_cdac_0.cdac_sw_8_1.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2511 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2512 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2513 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2514 VDREF single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2515 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2516 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2517 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2518 a_58494_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2519 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2520 a_13869_24944# single_10b_cdac_1.cdac_sw_4_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2521 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2522 VDREF single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2523 single_10b_cdac_1.x10b_cap_array_0.SW[5] single_10b_cdac_1.cdac_sw_4_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2524 VCM single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2525 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2526 VSREF single_10b_cdac_0.x2[0].x1.x9.A single_10b_cdac_0.x2[0].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2527 a_53071_35702# CF[4] single_10b_cdac_0.x6[4].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2528 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2529 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2530 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2531 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2532 VSREF single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2533 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2534 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2535 single_10b_cdac_1.x4[2].x2.swn single_10b_cdac_1.x4[2].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2536 single_10b_cdac_0.cdac_sw_8_0.x1.x6.A single_10b_cdac_0.cdac_sw_8_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2537 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2538 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2539 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2540 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2541 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2542 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x8.A single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2543 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2544 single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2545 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2546 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2547 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2548 single_10b_cdac_1.cdac_sw_1_2.x2.swn single_10b_cdac_1.cdac_sw_1_2.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2549 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2550 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2551 single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2552 single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.cdac_sw_8_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2553 single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2554 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2555 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2556 a_52054_34009# SWP_IN[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2557 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2558 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2559 single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2560 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2561 a_17874_25713# single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2562 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2563 single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2564 VDREF CF[8] single_10b_cdac_1.x10[8].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2565 VCN single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2566 VDREF single_10b_cdac_1.x6[4].x1.x5.A single_10b_cdac_1.x6[4].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2567 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2568 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2569 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2570 single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2571 a_19338_33146# single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2572 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2573 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2574 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2575 single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2576 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2577 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2578 single_10b_cdac_1.x2[0].x1.x6.A single_10b_cdac_1.x2[0].x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2579 VDREF single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2580 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2581 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2582 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2583 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2584 VDREF single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2585 VSREF single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2586 single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2587 single_10b_cdac_1.x6[5].x2.swn single_10b_cdac_1.x6[5].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2588 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2589 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2590 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2591 single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2592 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2593 single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2594 single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2595 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2596 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2597 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x7.A single_10b_cdac_0.cdac_sw_1_2.x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2598 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2599 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2600 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2601 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2602 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2603 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2604 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2605 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2606 single_10b_cdac_1.x3[0].x3.ck single_10b_cdac_1.x3[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2607 single_10b_cdac_0.cdac_sw_1_1.x1.x9.A single_10b_cdac_0.cdac_sw_1_1.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2608 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2609 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2610 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2611 single_10b_cdac_0.cdac_sw_8_1.x1.x4.A CF[2] a_41023_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2612 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2613 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x9.A single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2614 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2615 single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2616 VCN single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2617 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2618 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2619 single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2620 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2621 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2622 VSREF single_10b_cdac_0.x3[0].x1.x3.Y a_65951_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2623 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2624 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2625 single_10b_cdac_1.cdac_sw_8_1.x1.x6.A single_10b_cdac_1.cdac_sw_8_1.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2626 VCM single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2627 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2628 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2629 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2630 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2631 VDREF single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2632 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2633 VSREF single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2634 single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2635 single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2636 VDREF single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2637 VCM single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2638 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2639 single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2640 a_60343_24080# single_10b_cdac_0.cdac_sw_1_1.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2641 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2642 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2643 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2644 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2645 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2646 a_8214_25713# single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2647 single_10b_cdac_0.cdac_sw_16_0.x1.x3.Y CF[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2648 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2649 single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2650 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2651 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2652 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2653 VSREF single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2654 VSREF single_10b_cdac_1.x6[5].x1.x4.A single_10b_cdac_1.x6[5].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2655 single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2656 VDREF single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2657 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2658 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x8.A single_10b_cdac_1.cdac_sw_16_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2659 single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2660 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2661 VDREF single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2662 VDREF single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2663 VCM single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2664 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2665 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2666 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2667 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2668 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2669 VSREF single_10b_cdac_0.x8[6].x1.x9.A a_46631_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2670 single_10b_cdac_1.x10[8].x3.ck single_10b_cdac_1.x10[8].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2671 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2672 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2673 single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2674 VDREF single_10b_cdac_0.x8[7].x1.x9.A single_10b_cdac_0.x8[7].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2675 VSREF single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2676 single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2677 VCM single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2678 VDREF single_10b_cdac_1.x3[0].x1.x4.A single_10b_cdac_1.x3[0].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2679 single_10b_cdac_1.x10b_cap_array_0.SW[4] single_10b_cdac_1.cdac_sw_4_1.x3.ckb a_13776_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2680 VSREF single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2681 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2682 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2683 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2684 single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2685 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2686 VDREF single_10b_cdac_1.x6[4].x1.x9.A single_10b_cdac_1.x6[4].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2687 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2688 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2689 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2690 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2691 single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.cdac_sw_2_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2692 single_10b_cdac_1.x4[2].x3.ck single_10b_cdac_1.x4[2].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2693 VSREF single_10b_cdac_0.x8[6].x1.x6.A single_10b_cdac_0.x8[6].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2694 VDREF single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2695 VDREF CF[1] single_10b_cdac_1.x2[0].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2696 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2697 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2698 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2699 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2700 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2701 single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2702 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2703 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2704 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2705 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2706 single_10b_cdac_1.cdac_sw_8_0.x1.x8.A single_10b_cdac_1.cdac_sw_8_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2707 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2708 single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2709 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2710 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x8.A single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2711 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2712 single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2713 single_10b_cdac_0.cdac_sw_1_2.x3.ck single_10b_cdac_0.cdac_sw_1_2.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2714 VCM single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2715 VSREF single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2716 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2717 single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.cdac_sw_2_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2718 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2719 VDREF single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2720 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2721 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2722 VDREF single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2723 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2724 a_44150_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2725 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2726 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2727 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2728 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2729 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2730 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2731 VDREF SWP_IN[3] a_22558_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2732 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2733 single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.cdac_sw_2_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2734 single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2735 a_21680_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2736 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2737 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2738 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2739 VSREF single_10b_cdac_1.x10[8].x1.x4.A single_10b_cdac_1.x10[8].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2740 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2741 VSREF single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2742 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2743 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2744 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2745 single_10b_cdac_0.cdac_sw_1_1.x2.swn single_10b_cdac_0.cdac_sw_1_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2746 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2747 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2748 single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.cdac_sw_16_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2749 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2750 VSREF single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2751 VSREF SWN_IN[2] a_8214_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2752 single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2753 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2754 VDREF single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2755 VDREF single_10b_cdac_0.x6[4].x1.x6.A single_10b_cdac_0.x6[4].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2756 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2757 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2758 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2759 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x8.A single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2760 single_10b_cdac_0.x8[6].x2.swn single_10b_cdac_0.x8[6].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2761 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2762 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2763 single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.cdac_sw_8_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2764 VSREF single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2765 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2766 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2767 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2768 single_10b_cdac_0.x8[7].x3.ck single_10b_cdac_0.x8[7].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2769 single_10b_cdac_0.cdac_sw_2_1.x1.x5.A single_10b_cdac_0.cdac_sw_2_1.x1.x8.A a_53903_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2770 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2771 single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2772 VDREF single_10b_cdac_1.x8[7].x1.x9.A single_10b_cdac_1.x8[7].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2773 single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2774 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2775 single_10b_cdac_0.cdac_sw_1_0.x3.ck single_10b_cdac_0.cdac_sw_1_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2776 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x9.A single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2777 single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2778 VSREF single_10b_cdac_0.x3[0].x1.x6.A single_10b_cdac_0.x3[0].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2779 single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.cdac_sw_4_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2780 VDREF single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2781 single_10b_cdac_1.x6[4].x3.ck single_10b_cdac_1.x6[4].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2782 VCM single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2783 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2784 single_10b_cdac_1.cdac_sw_1_0.x1.x6.A single_10b_cdac_1.cdac_sw_1_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2785 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x4.A single_10b_cdac_0.cdac_sw_1_2.x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2786 single_10b_cdac_0.x4[2].x1.x5.A single_10b_cdac_0.x4[2].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2787 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x3.ck a_55274_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2788 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2789 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2790 a_53810_25722# SWN_IN[6] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2791 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2792 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2793 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2794 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2795 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x8.A single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2796 single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2797 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2798 VSREF single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2799 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2800 single_10b_cdac_0.x3[1].x2.swn single_10b_cdac_0.x3[1].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2801 single_10b_cdac_1.x10[8].x3.ck single_10b_cdac_1.x10[8].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2802 single_10b_cdac_1.x6[5].dac_out single_10b_cdac_1.x6[5].x3.ck a_15240_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2803 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2804 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2805 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2806 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2807 VSREF SWN_IN[2] a_41808_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2808 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2809 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2810 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2811 single_10b_cdac_1.x3[0].x3.ck single_10b_cdac_1.x3[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2812 VDREF single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2813 single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2814 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2815 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2816 VSREF single_10b_cdac_0.x6[5].x1.x9.A single_10b_cdac_0.x6[5].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2817 VDREF single_10b_cdac_1.x4[3].x1.x3.Y single_10b_cdac_1.x4[3].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2818 VDREF single_10b_cdac_0.x3[0].x1.x9.A single_10b_cdac_0.x3[0].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2819 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2820 single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2821 single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2822 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2823 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2824 single_10b_cdac_1.cdac_sw_2_1.x1.x9.A single_10b_cdac_1.cdac_sw_2_1.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2825 single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2826 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2827 single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2828 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2829 single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.cdac_sw_8_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2830 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2831 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2832 a_45028_25713# single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2833 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2834 VSREF single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2835 single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.cdac_sw_16_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2836 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2837 a_32357_35702# CF[0] single_10b_cdac_1.x3[0].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2838 VDREF SWP_IN[9] a_36832_34754# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2839 a_41808_25713# single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2840 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2841 single_10b_cdac_0.cdac_sw_4_0.x1.x5.A single_10b_cdac_0.cdac_sw_4_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2842 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2843 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2844 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2845 single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2846 single_10b_cdac_1.x10[8].dac_out single_10b_cdac_1.x10[8].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2847 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2848 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2849 VSREF single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2850 single_10b_cdac_0.x6[5].x2.swn single_10b_cdac_0.x6[5].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2851 VDREF single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2852 single_10b_cdac_0.x3[0].x2.swn single_10b_cdac_0.x3[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2853 VSREF single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2854 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2855 VDREF single_10b_cdac_1.x4[3].x1.x7.A single_10b_cdac_1.x4[3].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2856 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2857 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2858 a_20309_24080# single_10b_cdac_1.cdac_sw_2_1.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2859 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2860 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2861 single_10b_cdac_1.cdac_sw_1_1.x3.ck single_10b_cdac_1.cdac_sw_1_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2862 a_11434_25713# single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2863 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2864 single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2865 VSREF CF[9] single_10b_cdac_0.cdac_sw_1_2.x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2866 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2867 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2868 single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.cdac_sw_4_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2869 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2870 VDREF single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2871 single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2872 VDREF single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2873 VSREF single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2874 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2875 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2876 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2877 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2878 single_10b_cdac_0.cdac_sw_2_1.x1.x4.A single_10b_cdac_0.cdac_sw_2_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2879 VSREF single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2880 single_10b_cdac_1.x8[7].x3.ck single_10b_cdac_1.x8[7].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2881 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2882 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2883 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2884 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2885 VSREF single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2886 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2887 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2888 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2889 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x8.A single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2890 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2891 single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2892 VSREF single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2893 single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2894 single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x2[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2895 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2896 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2897 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2898 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2899 VSREF single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2900 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2901 VSREF single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2902 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2903 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2904 single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2905 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2906 VDREF single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2907 VSREF single_10b_cdac_0.x3[1].x1.x8.A single_10b_cdac_0.x3[1].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2908 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2909 single_10b_cdac_0.cdac_sw_16_0.x1.x9.A single_10b_cdac_0.cdac_sw_16_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2910 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2911 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2912 VDREF single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2913 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2914 single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.cdac_sw_4_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2915 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2916 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2917 single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.cdac_sw_8_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2918 VDREF single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2919 VDREF single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2920 single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2921 VSREF single_10b_cdac_1.x2[0].x1.x9.A single_10b_cdac_1.x2[0].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2922 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2923 VDREF single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2924 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2925 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2926 VSREF SWN_IN[3] a_45028_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2927 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2928 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2929 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2930 single_10b_cdac_1.x4[3].x3.ck single_10b_cdac_1.x4[3].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2931 single_10b_cdac_0.x6[5].dac_out single_10b_cdac_0.x6[5].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2932 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2933 single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2934 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2935 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2936 single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.cdac_sw_8_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2937 VSREF single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2938 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2939 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2940 VDREF single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2941 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2942 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2943 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2944 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2945 a_45614_34645# SWP_IN[6] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2946 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2947 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2948 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2949 a_51468_25713# single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2950 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2951 a_24900_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2952 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2953 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2954 single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2955 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2956 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2957 VDREF SWP_IN[2] a_25778_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2958 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2959 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2960 VDREF single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2961 single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2962 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2963 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2964 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2965 VSREF single_10b_cdac_1.x3[1].x1.x3.Y a_29137_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2966 VDREF single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2967 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2968 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2969 single_10b_cdac_1.x2[0].x1.x3.Y CF[1] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2970 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2971 VDREF single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2972 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2973 VDREF single_10b_cdac_1.x4[3].x1.x9.A single_10b_cdac_1.x4[3].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2974 VDREF single_10b_cdac_0.x3[0].x1.x8.A single_10b_cdac_0.x3[0].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2975 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2976 single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2977 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2978 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2979 single_10b_cdac_1.cdac_sw_1_1.x2.swn single_10b_cdac_1.cdac_sw_1_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2980 single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2981 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2982 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2983 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x9.A single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2984 a_5580_34963# SWP_IN[8] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2985 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2986 VCM single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2987 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2988 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2989 single_10b_cdac_1.x3[1].x1.x4.A CF[1] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2990 single_10b_cdac_0.x8[7].x1.x5.A single_10b_cdac_0.x8[7].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2991 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2992 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2993 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2994 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2995 single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2996 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2997 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2998 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x9.A single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2999 single_10b_cdac_0.x3[0].x3.ck single_10b_cdac_0.x3[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3000 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3001 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3002 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3003 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3004 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3005 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3006 a_13776_25722# SWN_IN[4] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3007 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3008 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3009 VCM single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3010 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3011 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3012 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3013 single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3014 single_10b_cdac_1.x6[5].x3.ck single_10b_cdac_1.x6[5].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3015 VDREF SWP_IN[2] a_25778_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3016 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3017 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3018 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3019 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3020 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x8.A single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3021 VSREF single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3022 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3023 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3024 single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3025 single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3026 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3027 VDREF single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3028 single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3029 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3030 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3031 VSREF single_10b_cdac_1.x6[4].x1.x7.A single_10b_cdac_1.x6[4].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3032 single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3033 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3034 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3035 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3036 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3037 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3038 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3039 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3040 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3041 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3042 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3043 single_10b_cdac_1.cdac_sw_2_0.x1.x4.A CF[7] a_23529_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3044 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3045 VSREF single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3046 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3047 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3048 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3049 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3050 VDREF single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3051 a_46492_34218# single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3052 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3053 single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3054 VDREF single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3055 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3056 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3057 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3058 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3059 VSREF single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3060 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3061 single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.cdac_sw_8_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3062 VCM single_10b_cdac_1.cdac_sw_1_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[9] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3063 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3064 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3065 single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3066 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x8.A single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3067 VDREF single_10b_cdac_0.x4[2].x1.x8.A single_10b_cdac_0.x4[2].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3068 VSREF single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3069 single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3070 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3071 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3072 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3073 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3074 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3075 single_10b_cdac_1.cdac_sw_4_0.x1.x3.Y CF[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3076 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3077 single_10b_cdac_0.x10b_cap_array_0.SW[4] single_10b_cdac_0.cdac_sw_4_1.x3.ckb a_47370_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3078 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3079 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3080 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3081 VDREF single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3082 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3083 single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3084 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3085 single_10b_cdac_0.cdac_sw_1_0.x3.ck single_10b_cdac_0.cdac_sw_1_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3086 single_10b_cdac_0.x3[1].x1.x5.A single_10b_cdac_0.x3[1].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3087 VDREF single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3088 VDREF CF[8] single_10b_cdac_1.cdac_sw_1_1.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3089 single_10b_cdac_1.x6[4].x3.ck single_10b_cdac_1.x6[4].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3090 VDREF single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3091 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3092 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x8.A single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3093 single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3094 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3095 single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3096 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3097 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3098 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3099 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3100 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3101 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3102 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3103 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3104 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3105 VCM single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3106 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3107 VSREF single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3108 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3109 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3110 VSREF single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3111 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3112 single_10b_cdac_1.cdac_sw_16_0.x1.x9.A single_10b_cdac_1.cdac_sw_16_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3113 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3114 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3115 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x8.A single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3116 single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3117 single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3118 VDREF single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3119 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3120 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x9.A single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3121 VSREF single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3122 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3123 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3124 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3125 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3126 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x3.ck a_24900_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3127 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3128 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3129 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3130 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3131 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3132 single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3133 VSREF single_10b_cdac_1.x3[1].x1.x9.A single_10b_cdac_1.x3[1].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3134 VDREF single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3135 VSREF SWN_IN[3] a_11434_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3136 VDREF single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3137 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3138 single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.cdac_sw_2_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3139 VSREF single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3140 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3141 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3142 single_10b_cdac_1.x4[2].x3.ck single_10b_cdac_1.x4[2].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3143 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3144 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3145 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3146 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3147 single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3148 VSREF single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3149 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3150 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3151 single_10b_cdac_1.x2[0].x1.x8.A single_10b_cdac_1.x2[0].x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3152 VSREF single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3153 VDREF single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3154 single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3155 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3156 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3157 single_10b_cdac_0.cdac_sw_1_1.x1.x7.A single_10b_cdac_0.cdac_sw_1_1.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3158 VDREF single_10b_cdac_1.x10[8].x1.x9.A single_10b_cdac_1.x10[8].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3159 single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3160 VDREF single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3161 VSREF single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3162 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3163 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3164 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3165 single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3166 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3167 single_10b_cdac_0.cdac_sw_4_1.x1.x5.A single_10b_cdac_0.cdac_sw_4_1.x1.x8.A a_47463_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3168 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3169 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3170 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3171 VSREF single_10b_cdac_1.x8[6].x1.x3.Y a_13037_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3172 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3173 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3174 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3175 single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.cdac_sw_2_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3176 single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3177 single_10b_cdac_1.cdac_sw_8_0.x1.x6.A single_10b_cdac_1.cdac_sw_8_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3178 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3179 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3180 VDREF single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3181 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3182 single_10b_cdac_1.x2[0].x1.x4.A single_10b_cdac_1.x2[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3183 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3184 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3185 single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.cdac_sw_8_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3186 VDREF single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3187 single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3188 single_10b_cdac_0.x10b_cap_array_0.SW[9] single_10b_cdac_0.cdac_sw_1_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3189 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3190 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3191 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3192 VDREF single_10b_cdac_1.x10[8].x1.x6.A single_10b_cdac_1.x10[8].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3193 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3194 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3195 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3196 single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3197 VSREF single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3198 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3199 single_10b_cdac_1.x3[1].x2.swn single_10b_cdac_1.x3[1].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3200 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3201 single_10b_cdac_0.cdac_sw_1_0.x1.x6.A single_10b_cdac_0.cdac_sw_1_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3202 single_10b_cdac_0.cdac_sw_8_0.x1.x9.A single_10b_cdac_0.cdac_sw_8_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3203 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3204 VSREF single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3205 a_56152_31002# single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3206 single_10b_cdac_1.x8[6].x1.x4.A CF[6] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3207 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3208 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3209 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3210 VDREF single_10b_cdac_0.x2[0].x1.x9.A single_10b_cdac_0.x2[0].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3211 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3212 single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3213 single_10b_cdac_1.cdac_sw_8_1.x1.x5.A single_10b_cdac_1.cdac_sw_8_1.x1.x8.A a_7429_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3214 VDREF single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3215 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3216 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3217 VDREF single_10b_cdac_1.x6[5].x1.x3.Y single_10b_cdac_1.x6[5].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3218 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3219 single_10b_cdac_1.cdac_sw_4_1.x1.x9.A single_10b_cdac_1.cdac_sw_4_1.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3220 a_58494_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3221 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3222 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3223 single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3224 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3225 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3226 VDREF single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3227 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3228 single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3229 VDREF single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3230 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3231 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3232 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x3.ck a_58494_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3233 single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.cdac_sw_4_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3234 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3235 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3236 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3237 single_10b_cdac_0.cdac_sw_8_0.x1.x5.A single_10b_cdac_0.cdac_sw_8_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3238 VDREF single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3239 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3240 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3241 single_10b_cdac_1.x6[4].dac_out single_10b_cdac_1.x6[4].x3.ck a_18460_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3242 single_10b_cdac_0.x3[1].x3.ck single_10b_cdac_0.x3[1].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3243 VSREF single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3244 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3245 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3246 VDREF single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3247 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3248 single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3249 single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.cdac_sw_2_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3250 single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3251 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3252 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3253 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3254 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3255 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3256 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3257 VSREF single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3258 single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3259 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3260 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3261 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3262 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3263 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3264 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3265 VDREF single_10b_cdac_0.x4[3].x1.x7.A single_10b_cdac_0.x4[3].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3266 VCM single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3267 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3268 VDREF single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3269 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3270 VSREF single_10b_cdac_1.x3[0].x1.x3.Y a_32357_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3271 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3272 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3273 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3274 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3275 a_45028_25713# single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3276 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3277 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3278 VCM single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3279 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3280 single_10b_cdac_0.cdac_sw_4_1.x1.x4.A single_10b_cdac_0.cdac_sw_4_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3281 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3282 VDREF CF[8] single_10b_cdac_0.cdac_sw_1_1.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3283 VDREF SWP_IN[4] a_19338_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3284 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3285 VCM single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3286 single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.cdac_sw_8_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3287 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3288 VDREF single_10b_cdac_0.x8[7].x1.x8.A single_10b_cdac_0.x8[7].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3289 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3290 single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.cdac_sw_16_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3291 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3292 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3293 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3294 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3295 single_10b_cdac_1.cdac_sw_1_1.x2.swn single_10b_cdac_1.cdac_sw_1_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3296 single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3297 single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3298 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3299 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3300 single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3301 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3302 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3303 VDREF CF[3] single_10b_cdac_1.cdac_sw_8_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3304 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3305 VDREF single_10b_cdac_0.x10[8].x1.x5.A single_10b_cdac_0.x10[8].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3306 single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3307 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3308 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3309 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x3.ckb a_40930_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3310 VSREF CF[4] single_10b_cdac_1.x6[4].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3311 a_25778_31002# single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3312 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3313 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3314 VSREF single_10b_cdac_0.x4[3].x1.x8.A single_10b_cdac_0.x4[3].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3315 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3316 a_40052_34754# single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3317 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3318 single_10b_cdac_1.x4[3].x1.x5.A single_10b_cdac_1.x4[3].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3319 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3320 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3321 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3322 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3323 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3324 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x9.A single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3325 a_63563_24944# single_10b_cdac_0.cdac_sw_1_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3326 VDREF single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3327 VDREF single_10b_cdac_1.x10[8].x1.x8.A single_10b_cdac_1.x10[8].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3328 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3329 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3330 VSREF single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3331 VDREF single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3332 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3333 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3334 VCM single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3335 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3336 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3337 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3338 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3339 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3340 VSREF single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3341 single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.cdac_sw_16_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3342 VSREF single_10b_cdac_1.x8[6].x1.x9.A single_10b_cdac_1.x8[6].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3343 single_10b_cdac_0.x4[3].x3.ck single_10b_cdac_0.x4[3].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3344 VDREF single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3345 single_10b_cdac_0.x6[5].x2.swn single_10b_cdac_0.x6[5].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3346 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3347 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3348 single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x2[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3349 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3350 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3351 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3352 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3353 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3354 VSREF SWN_IN[2] a_8214_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3355 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3356 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3357 VSREF single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3358 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3359 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3360 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3361 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3362 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3363 VDREF single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3364 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3365 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3366 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3367 VDREF single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3368 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3369 single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3370 a_25778_31002# single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3371 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3372 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3373 VDREF SWP_IN[2] a_59372_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3374 VSREF single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3375 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3376 VDREF single_10b_cdac_0.x2[0].x1.x8.A single_10b_cdac_0.x2[0].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3377 single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3378 single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3379 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3380 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3381 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3382 single_10b_cdac_1.x4[3].x3.ck single_10b_cdac_1.x4[3].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3383 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3384 single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.cdac_sw_4_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3385 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3386 single_10b_cdac_0.x3[0].x2.swn single_10b_cdac_0.x3[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3387 single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3388 VSREF single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3389 VCM single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3390 single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.cdac_sw_8_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3391 a_10556_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3392 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3393 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3394 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3395 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3396 VDREF single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3397 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3398 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3399 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3400 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3401 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3402 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3403 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3404 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3405 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x9.A a_3377_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3406 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3407 single_10b_cdac_1.cdac_sw_1_1.x3.ck single_10b_cdac_1.cdac_sw_1_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3408 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3409 single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3410 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3411 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3412 VDREF single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3413 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3414 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3415 single_10b_cdac_1.x8[6].x2.swn single_10b_cdac_1.x8[6].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3416 single_10b_cdac_0.x4[2].x3.ck single_10b_cdac_0.x4[2].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3417 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3418 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3419 VDREF single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3420 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3421 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3422 VSREF single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3423 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3424 single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3425 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3426 single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3427 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3428 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3429 single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3430 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3431 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3432 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3433 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3434 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3435 single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3436 VCP single_10b_cdac_0.x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3437 VSREF single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3438 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3439 VDREF single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3440 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3441 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3442 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3443 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3444 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x9.A single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3445 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3446 VDREF single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3447 single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.cdac_sw_16_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3448 VSREF single_10b_cdac_1.x3[0].x1.x6.A single_10b_cdac_1.x3[0].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3449 VCN single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3450 VDREF single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3451 VDREF SWP_IN[2] a_59372_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3452 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3453 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3454 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3455 a_52932_33146# single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3456 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3457 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3458 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3459 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3460 single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3461 single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3462 single_10b_cdac_1.x8[6].dac_out single_10b_cdac_1.x8[6].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3463 a_53071_36566# single_10b_cdac_0.x6[4].x1.x8.A single_10b_cdac_0.x6[4].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3464 VSREF single_10b_cdac_0.x3[0].x1.x4.A single_10b_cdac_0.x3[0].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3465 single_10b_cdac_1.cdac_sw_4_0.x1.x4.A CF[5] a_17089_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3466 VCM single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3467 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3468 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3469 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3470 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3471 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3472 single_10b_cdac_1.cdac_sw_1_0.x2.swn single_10b_cdac_1.cdac_sw_1_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3473 VSREF single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3474 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x3.ckb a_44150_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3475 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3476 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3477 single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.cdac_sw_8_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3478 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3479 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3480 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x8.A single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3481 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3482 single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3483 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3484 single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3485 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3486 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3487 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3488 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3489 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3490 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3491 VSREF single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3492 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3493 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3494 single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3495 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3496 VCM single_10b_cdac_0.cdac_sw_1_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[9] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3497 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3498 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3499 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3500 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3501 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3502 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3503 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3504 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3505 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3506 single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.cdac_sw_4_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3507 single_10b_cdac_1.cdac_sw_1_2.x2.swn single_10b_cdac_1.cdac_sw_1_2.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3508 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3509 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3510 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3511 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3512 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3513 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3514 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3515 single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3516 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3517 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3518 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x9.A single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3519 VSREF single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3520 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3521 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3522 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3523 single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.cdac_sw_4_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3524 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3525 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3526 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3527 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3528 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3529 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3530 single_10b_cdac_0.x2[0].x1.x6.A single_10b_cdac_0.x2[0].x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3531 VSREF single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3532 single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3533 single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3534 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3535 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3536 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3537 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3538 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3539 VSREF single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3540 single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x2[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3541 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3542 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3543 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x9.A single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3544 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3545 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3546 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3547 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x9.A single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3548 VDREF CF[3] single_10b_cdac_0.x4[3].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3549 VDREF single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3550 single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3551 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3552 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3553 VDREF single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3554 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3555 single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3556 VSREF single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3557 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3558 a_47370_25722# SWN_IN[4] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3559 a_23529_24944# single_10b_cdac_1.cdac_sw_2_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3560 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3561 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3562 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3563 single_10b_cdac_1.cdac_sw_2_1.x1.x3.Y CF[6] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3564 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3565 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3566 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3567 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3568 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3569 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3570 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3571 VSREF single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3572 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3573 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3574 single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3575 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3576 single_10b_cdac_0.cdac_sw_2_1.x1.x6.A single_10b_cdac_0.cdac_sw_2_1.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3577 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3578 VSREF single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3579 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3580 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3581 single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3582 VDREF single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3583 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3584 VSREF single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3585 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3586 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3587 VDREF single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3588 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3589 single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3590 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3591 VSREF single_10b_cdac_1.x6[5].x1.x5.A single_10b_cdac_1.x6[5].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3592 single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3593 single_10b_cdac_1.cdac_sw_1_2.dac_out single_10b_cdac_1.cdac_sw_1_2.x3.ck a_2360_34963# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3594 VSREF SWN_IN[3] a_11434_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3595 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3596 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3597 single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3598 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3599 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3600 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3601 VSREF single_10b_cdac_0.x8[6].x1.x3.Y a_46631_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3602 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3603 single_10b_cdac_1.x10[8].x2.swn single_10b_cdac_1.x10[8].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3604 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3605 single_10b_cdac_1.cdac_sw_1_1.x1.x4.A single_10b_cdac_1.cdac_sw_1_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3606 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3607 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3608 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3609 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3610 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3611 VSREF single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3612 VDREF single_10b_cdac_1.x4[3].x1.x8.A single_10b_cdac_1.x4[3].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3613 a_12020_34645# SWP_IN[6] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3614 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3615 VDREF single_10b_cdac_1.x3[1].x1.x6.A single_10b_cdac_1.x3[1].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3616 single_10b_cdac_0.x2[0].x1.x8.A single_10b_cdac_0.x2[0].x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3617 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3618 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3619 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3620 a_41023_24080# single_10b_cdac_0.cdac_sw_8_1.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3621 single_10b_cdac_0.cdac_sw_2_0.x1.x6.A single_10b_cdac_0.cdac_sw_2_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3622 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3623 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3624 single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.cdac_sw_8_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3625 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3626 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3627 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3628 single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3629 single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3630 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3631 VDREF single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3632 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3633 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x9.A single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3634 single_10b_cdac_0.x8[7].x3.ck single_10b_cdac_0.x8[7].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3635 VDREF single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3636 VSREF single_10b_cdac_0.x8[6].x1.x7.A single_10b_cdac_0.x8[6].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3637 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3638 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3639 single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3640 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3641 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3642 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3643 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3644 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3645 VDREF single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3646 VDREF single_10b_cdac_0.x6[5].x1.x3.Y single_10b_cdac_0.x6[5].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3647 single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3648 VSREF single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3649 single_10b_cdac_0.cdac_sw_1_2.x2.swn single_10b_cdac_0.cdac_sw_1_2.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3650 VDREF single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3651 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3652 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3653 VDREF SWP_IN[7] a_43272_34218# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3654 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3655 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3656 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3657 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3658 single_10b_cdac_0.x4[3].x3.ck single_10b_cdac_0.x4[3].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3659 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3660 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3661 VSREF single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3662 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3663 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3664 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3665 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3666 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3667 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3668 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3669 single_10b_cdac_1.x3[1].x2.swn single_10b_cdac_1.x3[1].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3670 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3671 single_10b_cdac_1.x10[8].x1.x4.A CF[8] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3672 single_10b_cdac_0.x8[6].dac_out single_10b_cdac_0.x8[6].x3.ck a_45614_34645# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3673 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3674 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3675 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3676 VSREF single_10b_cdac_1.x10[8].x1.x5.A single_10b_cdac_1.x10[8].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3677 VDREF single_10b_cdac_0.x6[5].x1.x7.A single_10b_cdac_0.x6[5].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3678 a_56152_31002# single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3679 a_55274_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3680 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3681 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3682 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3683 VSREF SWN_IN[5] a_51468_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3684 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3685 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3686 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3687 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3688 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3689 VDREF single_10b_cdac_1.x8[7].x1.x3.Y single_10b_cdac_1.x8[7].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3690 VSREF single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3691 single_10b_cdac_1.cdac_sw_8_1.x1.x9.A single_10b_cdac_1.cdac_sw_8_1.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3692 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3693 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3694 VDREF single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3695 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3696 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x8.A single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3697 single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3698 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3699 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3700 single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3701 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3702 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3703 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3704 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3705 VDREF single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3706 single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3707 a_40930_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3708 VDREF single_10b_cdac_0.x6[4].x1.x9.A single_10b_cdac_0.x6[4].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3709 VSREF single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3710 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3711 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3712 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3713 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3714 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3715 single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3716 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3717 VDREF single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3718 VDREF single_10b_cdac_1.x8[7].x1.x7.A single_10b_cdac_1.x8[7].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3719 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3720 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3721 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3722 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3723 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3724 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3725 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3726 VSREF single_10b_cdac_0.x3[0].x1.x7.A single_10b_cdac_0.x3[0].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3727 single_10b_cdac_0.cdac_sw_1_2.x3.ck single_10b_cdac_0.cdac_sw_1_2.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3728 a_7429_24080# single_10b_cdac_1.cdac_sw_8_1.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3729 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3730 single_10b_cdac_1.cdac_sw_1_1.x1.x7.A single_10b_cdac_1.cdac_sw_1_1.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3731 single_10b_cdac_1.x6[5].x1.x5.A single_10b_cdac_1.x6[5].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3732 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3733 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3734 single_10b_cdac_0.cdac_sw_1_0.x2.swn single_10b_cdac_0.cdac_sw_1_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3735 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3736 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3737 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3738 single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3739 VDREF single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3740 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3741 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3742 single_10b_cdac_0.x6[4].x2.swn single_10b_cdac_0.x6[4].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3743 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3744 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3745 single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3746 single_10b_cdac_0.x10b_cap_array_0.SW[5] single_10b_cdac_0.cdac_sw_4_0.x3.ckb a_50590_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3747 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3748 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3749 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3750 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3751 single_10b_cdac_1.x10[8].x2.swn single_10b_cdac_1.x10[8].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3752 single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3753 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3754 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3755 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3756 single_10b_cdac_1.cdac_sw_1_0.x3.ck single_10b_cdac_1.cdac_sw_1_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3757 VSREF single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3758 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3759 single_10b_cdac_0.x6[5].x3.ck single_10b_cdac_0.x6[5].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3760 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3761 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3762 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3763 VDREF CF[8] single_10b_cdac_0.x10[8].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3764 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3765 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3766 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3767 single_10b_cdac_1.x3[0].x2.swn single_10b_cdac_1.x3[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3768 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3769 VSREF single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3770 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3771 single_10b_cdac_0.x6[5].x1.x4.A CF[5] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3772 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3773 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3774 single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3775 single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3776 VDREF single_10b_cdac_0.x3[1].x1.x9.A single_10b_cdac_0.x3[1].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3777 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x3.ck a_21680_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3778 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3779 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3780 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3781 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3782 a_32357_36566# single_10b_cdac_1.x3[0].x1.x8.A single_10b_cdac_1.x3[0].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3783 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3784 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3785 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3786 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x8.A single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3787 VDREF single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3788 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3789 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3790 single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3791 a_19338_33146# single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3792 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3793 VDREF single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3794 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3795 single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3796 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3797 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3798 VDREF single_10b_cdac_0.x3[1].x1.x6.A single_10b_cdac_0.x3[1].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3799 VDREF single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3800 single_10b_cdac_1.x8[7].x3.ck single_10b_cdac_1.x8[7].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3801 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3802 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3803 VCP single_10b_cdac_0.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3804 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3805 VDREF single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3806 single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3807 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3808 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3809 single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.cdac_sw_2_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3810 VDREF single_10b_cdac_0.x8[6].x1.x9.A single_10b_cdac_0.x8[6].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3811 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3812 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3813 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3814 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3815 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3816 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3817 single_10b_cdac_1.cdac_sw_8_0.x1.x4.A single_10b_cdac_1.cdac_sw_8_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3818 a_27534_25713# single_10b_cdac_1.cdac_sw_1_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[8] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3819 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3820 single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3821 single_10b_cdac_0.x6[4].x3.ck single_10b_cdac_0.x6[4].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3822 VDREF single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3823 a_7336_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3824 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3825 VDREF single_10b_cdac_1.x8[6].x1.x6.A single_10b_cdac_1.x8[6].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3826 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3827 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3828 single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3829 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3830 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3831 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3832 single_10b_cdac_0.cdac_sw_8_1.x1.x6.A single_10b_cdac_0.cdac_sw_8_1.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3833 VSREF single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3834 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3835 single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.cdac_sw_2_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3836 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3837 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3838 single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.cdac_sw_4_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3839 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3840 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3841 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3842 single_10b_cdac_1.cdac_sw_4_1.x1.x5.A single_10b_cdac_1.cdac_sw_4_1.x1.x8.A a_13869_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3843 VDREF single_10b_cdac_0.x8[6].x1.x4.A single_10b_cdac_0.x8[6].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3844 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3845 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3846 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3847 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3848 single_10b_cdac_0.x3[0].x3.ck single_10b_cdac_0.x3[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3849 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3850 VSREF single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3851 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3852 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3853 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3854 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3855 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3856 single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.cdac_sw_2_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3857 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x9.A single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3858 VSREF single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3859 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x3.ck a_24900_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3860 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3861 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3862 VDREF single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3863 single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3864 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3865 VDREF single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3866 VSREF single_10b_cdac_0.x3[1].x1.x9.A single_10b_cdac_0.x3[1].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3867 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3868 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3869 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3870 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3871 VCN single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3872 single_10b_cdac_1.x10b_cap_array_0.SW[9] single_10b_cdac_1.cdac_sw_1_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3873 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3874 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x9.A single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3875 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3876 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3877 VSREF single_10b_cdac_0.x4[2].x1.x4.A single_10b_cdac_0.x4[2].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3878 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3879 single_10b_cdac_1.cdac_sw_16_0.x1.x6.A single_10b_cdac_1.cdac_sw_16_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3880 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3881 single_10b_cdac_1.x4[3].x2.swn single_10b_cdac_1.x4[3].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3882 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3883 a_26656_25722# SWN_IN[8] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3884 a_54688_25713# single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[6] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3885 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3886 single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3887 single_10b_cdac_1.x8[6].x2.swn single_10b_cdac_1.x8[6].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3888 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3889 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3890 VSREF single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3891 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3892 single_10b_cdac_0.cdac_sw_1_0.x2.swn single_10b_cdac_0.cdac_sw_1_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3893 VCM single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3894 a_51468_25713# single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3895 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3896 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3897 VSREF single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3898 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3899 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3900 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3901 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3902 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3903 VSREF single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3904 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3905 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3906 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3907 single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.cdac_sw_4_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3908 VCP single_10b_cdac_1.x3[1].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3909 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3910 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3911 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3912 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3913 single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3914 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3915 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3916 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3917 single_10b_cdac_0.x8[6].x3.ck single_10b_cdac_0.x8[6].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3918 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3919 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3920 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3921 a_3377_35702# CF[9] single_10b_cdac_1.cdac_sw_1_2.x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3922 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3923 single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3924 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3925 single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3926 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3927 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3928 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3929 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3930 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3931 VCM single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3932 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x8.A single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3933 single_10b_cdac_1.cdac_sw_1_2.x2.swn single_10b_cdac_1.cdac_sw_1_2.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3934 single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3935 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3936 single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.cdac_sw_8_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3937 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3938 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3939 single_10b_cdac_1.cdac_sw_4_0.x1.x8.A single_10b_cdac_1.cdac_sw_4_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3940 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3941 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3942 single_10b_cdac_1.cdac_sw_4_0.x1.x7.A single_10b_cdac_1.cdac_sw_4_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3943 single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3944 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3945 single_10b_cdac_0.x4[2].x3.ck single_10b_cdac_0.x4[2].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3946 VDREF single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3947 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3948 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3949 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3950 single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3951 single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.cdac_sw_4_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3952 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3953 VDREF single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3954 single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3955 VCN single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3956 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3957 single_10b_cdac_0.cdac_sw_4_0.x1.x7.A single_10b_cdac_0.cdac_sw_4_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3958 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3959 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3960 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3961 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3962 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3963 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3964 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3965 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3966 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x3.ck a_58494_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3967 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3968 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3969 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3970 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3971 VDREF single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3972 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3973 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3974 a_17089_24944# single_10b_cdac_1.cdac_sw_4_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3975 single_10b_cdac_1.x6[5].x2.swn single_10b_cdac_1.x6[5].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3976 single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3977 single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3978 single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3979 VDREF single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3980 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3981 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3982 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3983 VSREF single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3984 single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x2[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3985 VSREF single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3986 VSREF single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3987 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3988 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3989 single_10b_cdac_1.x10b_cap_array_0.SW[5] single_10b_cdac_1.cdac_sw_4_0.x3.ckb a_16996_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3990 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3991 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3992 single_10b_cdac_0.cdac_sw_2_1.x1.x3.Y CF[6] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3993 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3994 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3995 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3996 single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3997 single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3998 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3999 single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4000 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4001 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4002 single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x2[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4003 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4004 a_55274_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4005 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4006 VDREF single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4007 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4008 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4009 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4010 VSREF CF[0] single_10b_cdac_0.x3[0].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4011 single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4012 a_46631_35702# CF[6] single_10b_cdac_0.x8[6].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4013 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4014 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4015 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4016 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4017 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4018 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4019 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4020 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4021 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4022 VDREF single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4023 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4024 VSREF single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4025 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4026 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4027 VDREF single_10b_cdac_1.x6[5].x1.x8.A single_10b_cdac_1.x6[5].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4028 VDREF single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4029 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4030 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4031 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4032 a_11434_25713# single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4033 single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x2[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4034 a_34583_24080# single_10b_cdac_0.cdac_sw_16_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4035 single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4036 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4037 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4038 single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4039 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4040 single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4041 VDREF single_10b_cdac_1.x3[0].x1.x9.A single_10b_cdac_1.x3[0].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4042 VSREF single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4043 single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4044 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4045 VDREF single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4046 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4047 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4048 VSREF single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4049 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4050 single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.cdac_sw_8_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4051 VDREF single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4052 single_10b_cdac_0.cdac_sw_1_0.x1.x9.A single_10b_cdac_0.cdac_sw_1_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4053 VDREF single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4054 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4055 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4056 VSREF single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4057 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4058 VSREF single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4059 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4060 single_10b_cdac_0.x10b_cap_array_0.SW[4] single_10b_cdac_0.cdac_sw_4_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4061 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4062 VSREF single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4063 VDREF single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4064 single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4065 VSREF single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4066 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4067 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4068 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4069 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4070 VSREF single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4071 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4072 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4073 VSREF single_10b_cdac_0.x8[7].x1.x4.A single_10b_cdac_0.x8[7].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4074 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4075 single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.cdac_sw_8_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4076 single_10b_cdac_1.x4[2].x3.ck single_10b_cdac_1.x4[2].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4077 single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4078 VSREF single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4079 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4080 a_10556_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4081 single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x2[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4082 single_10b_cdac_0.cdac_sw_16_0.x1.x4.A CF[0] a_34583_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4083 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4084 VSREF SWN_IN[3] a_45028_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4085 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4086 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4087 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4088 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4089 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4090 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4091 VSREF single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4092 single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4093 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4094 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4095 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4096 single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4097 VDREF single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4098 VSREF single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4099 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4100 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4101 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4102 a_8214_25713# single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4103 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4104 VSREF single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4105 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4106 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4107 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4108 single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4109 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4110 single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4111 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4112 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4113 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4114 single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4115 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4116 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4117 VDREF single_10b_cdac_1.x4[2].x1.x9.A single_10b_cdac_1.x4[2].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4118 VSREF single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4119 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x3.ckb a_10556_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4120 single_10b_cdac_0.cdac_sw_1_1.x3.ck single_10b_cdac_0.cdac_sw_1_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4121 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4122 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4123 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4124 single_10b_cdac_1.cdac_sw_1_1.x1.x3.Y CF[8] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4125 single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.cdac_sw_4_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4126 a_29969_24080# single_10b_cdac_1.cdac_sw_1_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4127 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4128 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4129 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4130 single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.cdac_sw_16_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4131 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4132 VSREF single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4133 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4134 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x8.A single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4135 VDREF single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4136 VCM single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4137 single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4138 single_10b_cdac_0.x8[6].x2.swn single_10b_cdac_0.x8[6].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4139 single_10b_cdac_1.x6[4].dac_out single_10b_cdac_1.x6[4].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4140 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4141 single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4142 single_10b_cdac_0.x8[7].x3.ck single_10b_cdac_0.x8[7].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4143 a_10556_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4144 VSREF single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4145 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4146 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x3.ckb a_44150_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4147 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4148 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4149 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4150 single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4151 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4152 VSREF single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4153 VDREF single_10b_cdac_1.x4[2].x1.x4.A single_10b_cdac_1.x4[2].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4154 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4155 single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4156 VDREF single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4157 single_10b_cdac_1.x6[4].x3.ck single_10b_cdac_1.x6[4].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4158 single_10b_cdac_0.x6[4].dac_out single_10b_cdac_0.x6[4].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4159 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4160 single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4161 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4162 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4163 single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4164 VDREF single_10b_cdac_0.x4[3].x1.x9.A single_10b_cdac_0.x4[3].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4165 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4166 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4167 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4168 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4169 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4170 VSREF single_10b_cdac_0.x10[8].x1.x6.A single_10b_cdac_0.x10[8].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4171 single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4172 VDREF SWP_IN[2] a_25778_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4173 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4174 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4175 VSREF SWN_IN[6] a_21094_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4176 single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4177 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4178 single_10b_cdac_1.x8[7].x1.x5.A single_10b_cdac_1.x8[7].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4179 single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4180 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4181 single_10b_cdac_0.x3[1].x2.swn single_10b_cdac_0.x3[1].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4182 VSREF single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4183 single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.cdac_sw_4_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4184 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4185 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4186 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4187 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4188 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4189 VDREF single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4190 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4191 VDREF CF[3] single_10b_cdac_1.x4[3].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4192 single_10b_cdac_1.x10b_cap_array_0.SW[5] single_10b_cdac_1.cdac_sw_4_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4193 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4194 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4195 single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4196 single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4197 VSREF CF[5] single_10b_cdac_0.x6[5].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4198 single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.cdac_sw_4_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4199 VDREF single_10b_cdac_0.x10[8].x1.x9.A single_10b_cdac_0.x10[8].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4200 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4201 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4202 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x3.ckb a_44150_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4203 single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4204 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4205 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4206 single_10b_cdac_0.x8[6].x3.ck single_10b_cdac_0.x8[6].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4207 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4208 single_10b_cdac_0.cdac_sw_2_0.x1.x5.A single_10b_cdac_0.cdac_sw_2_0.x1.x8.A a_57123_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4209 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4210 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4211 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4212 VCP VCM sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4213 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4214 single_10b_cdac_1.cdac_sw_2_1.x1.x6.A single_10b_cdac_1.cdac_sw_2_1.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4215 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4216 VDREF single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4217 single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4218 VDREF single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4219 VSREF single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4220 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4221 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x8.A single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4222 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4223 single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4224 single_10b_cdac_0.x10[8].x2.swn single_10b_cdac_0.x10[8].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4225 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4226 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4227 single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4228 single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4229 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4230 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4231 single_10b_cdac_0.x4[2].x3.ck single_10b_cdac_0.x4[2].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4232 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4233 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4234 single_10b_cdac_0.cdac_sw_2_1.x1.x9.A single_10b_cdac_0.cdac_sw_2_1.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4235 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4236 VDREF single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4237 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4238 VDREF single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4239 single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4240 single_10b_cdac_1.x8[7].x3.ck single_10b_cdac_1.x8[7].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4241 VSREF single_10b_cdac_0.x4[3].x1.x9.A single_10b_cdac_0.x4[3].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4242 VDREF single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4243 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4244 single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4245 VDREF single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4246 single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4247 VDREF SWP_IN[4] a_52932_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4248 single_10b_cdac_1.cdac_sw_2_0.x1.x9.A single_10b_cdac_1.cdac_sw_2_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4249 single_10b_cdac_0.x6[4].dac_out single_10b_cdac_0.x6[4].x3.ck a_52054_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4250 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4251 single_10b_cdac_1.cdac_sw_2_0.x1.x6.A single_10b_cdac_1.cdac_sw_2_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4252 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4253 VCP single_10b_cdac_0.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4254 a_48248_25713# single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4255 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4256 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4257 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4258 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4259 single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.cdac_sw_2_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4260 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4261 single_10b_cdac_0.x4[3].x2.swn single_10b_cdac_0.x4[3].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4262 VDREF single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4263 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4264 single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4265 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4266 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4267 single_10b_cdac_0.cdac_sw_2_0.x1.x8.A single_10b_cdac_0.cdac_sw_2_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4268 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4269 VSREF single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4270 a_18460_34009# SWP_IN[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4271 VSREF single_10b_cdac_0.x3[1].x1.x8.A single_10b_cdac_0.x3[1].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4272 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4273 VDREF single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4274 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4275 single_10b_cdac_1.cdac_sw_1_0.x3.ck single_10b_cdac_1.cdac_sw_1_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4276 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4277 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4278 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4279 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4280 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4281 single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4282 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4283 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4284 single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4285 a_40930_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4286 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4287 a_41808_25713# single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4288 VDREF single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4289 VDREF single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4290 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4291 VSREF single_10b_cdac_1.x2[0].x1.x9.A single_10b_cdac_1.x2[0].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4292 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4293 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4294 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4295 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4296 single_10b_cdac_0.x10[8].x3.ck single_10b_cdac_0.x10[8].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4297 VDREF single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4298 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4299 single_10b_cdac_1.x4[3].x3.ck single_10b_cdac_1.x4[3].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4300 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4301 VSREF single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4302 a_24900_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4303 VCM single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4304 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4305 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4306 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4307 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4308 a_16996_25722# SWN_IN[5] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4309 single_10b_cdac_0.cdac_sw_2_0.x1.x4.A single_10b_cdac_0.cdac_sw_2_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4310 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4311 VCM single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4312 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4313 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4314 single_10b_cdac_1.x4[3].x2.swn single_10b_cdac_1.x4[3].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4315 single_10b_cdac_0.x4[3].x2.swn single_10b_cdac_0.x4[3].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4316 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4317 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4318 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4319 VDREF single_10b_cdac_1.x6[5].x1.x7.A single_10b_cdac_1.x6[5].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4320 a_21680_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4321 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4322 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4323 single_10b_cdac_1.cdac_sw_8_0.x1.x3.Y CF[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4324 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4325 a_13869_24080# single_10b_cdac_1.cdac_sw_4_1.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4326 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4327 VCN single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4328 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4329 VSREF single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4330 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4331 VDREF single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4332 VDREF CF[6] single_10b_cdac_1.cdac_sw_2_1.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4333 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x3.Y a_3377_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4334 single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4335 single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4336 VDREF single_10b_cdac_0.x6[5].x1.x5.A single_10b_cdac_0.x6[5].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4337 single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4338 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4339 single_10b_cdac_0.cdac_sw_8_0.x1.x7.A single_10b_cdac_0.cdac_sw_8_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4340 single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4341 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4342 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x9.A single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4343 VDREF single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4344 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4345 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4346 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4347 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4348 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4349 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4350 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4351 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4352 single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4353 single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4354 VSREF single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4355 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4356 VDREF single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4357 single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4358 VDREF single_10b_cdac_0.x10[8].x1.x9.A single_10b_cdac_0.x10[8].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4359 VSREF single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4360 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4361 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4362 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4363 VSREF single_10b_cdac_1.x3[0].x1.x7.A single_10b_cdac_1.x3[0].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4364 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4365 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4366 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4367 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4368 single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4369 VSREF single_10b_cdac_1.x4[3].x1.x4.A single_10b_cdac_1.x4[3].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4370 single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4371 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4372 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4373 single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4374 single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4375 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4376 single_10b_cdac_1.x2[0].x1.x7.A single_10b_cdac_1.x2[0].x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4377 VSREF single_10b_cdac_0.x3[0].x1.x5.A single_10b_cdac_0.x3[0].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4378 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4379 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x3.ck a_55274_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4380 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4381 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4382 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4383 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4384 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4385 VDREF single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4386 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4387 single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4388 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4389 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4390 VSREF single_10b_cdac_0.x6[4].x1.x9.A a_53071_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4391 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4392 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4393 single_10b_cdac_1.x6[5].x3.ck single_10b_cdac_1.x6[5].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4394 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4395 VDREF single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4396 a_7336_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4397 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4398 single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4399 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4400 single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4401 single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4402 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4403 single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4404 VSREF single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4405 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4406 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4407 single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4408 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4409 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4410 single_10b_cdac_1.cdac_sw_8_1.x1.x3.Y CF[2] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4411 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4412 single_10b_cdac_0.cdac_sw_8_1.x1.x5.A single_10b_cdac_0.cdac_sw_8_1.x1.x8.A a_41023_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4413 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4414 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4415 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4416 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4417 VDREF single_10b_cdac_1.x4[2].x1.x9.A single_10b_cdac_1.x4[2].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4418 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4419 a_45028_25713# single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4420 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4421 single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4422 single_10b_cdac_1.x3[0].x3.ck single_10b_cdac_1.x3[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4423 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4424 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4425 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4426 single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.cdac_sw_16_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4427 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4428 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4429 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4430 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4431 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4432 single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4433 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4434 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4435 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4436 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4437 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4438 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4439 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4440 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4441 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4442 VDREF single_10b_cdac_0.x4[2].x1.x8.A single_10b_cdac_0.x4[2].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4443 VSREF single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4444 VSREF single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4445 single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4446 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4447 single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4448 single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4449 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4450 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4451 VDREF single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4452 VDREF single_10b_cdac_1.x8[7].x1.x8.A single_10b_cdac_1.x8[7].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4453 single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4454 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x9.A single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4455 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4456 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4457 single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4458 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4459 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x3.ck a_21680_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4460 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4461 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4462 single_10b_cdac_1.x6[4].x3.ck single_10b_cdac_1.x6[4].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4463 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4464 VSREF single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4465 VDREF single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4466 single_10b_cdac_0.cdac_sw_1_2.x1.x5.A single_10b_cdac_0.cdac_sw_1_2.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4467 single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.cdac_sw_2_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4468 VDREF single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4469 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4470 VCM single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4471 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4472 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4473 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4474 single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4475 single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.cdac_sw_8_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4476 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4477 VCN single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4478 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4479 single_10b_cdac_0.cdac_sw_8_1.x1.x8.A single_10b_cdac_0.cdac_sw_8_1.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4480 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4481 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4482 VSREF single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4483 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4484 VSREF single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4485 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4486 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4487 VDREF SWP_IN[4] a_19338_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4488 single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4489 VDREF single_10b_cdac_0.x2[0].x1.x8.A single_10b_cdac_0.x2[0].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4490 single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4491 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4492 single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4493 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4494 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4495 VSREF single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4496 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x6.A single_10b_cdac_1.cdac_sw_1_2.x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4497 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4498 single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4499 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4500 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4501 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4502 VDREF single_10b_cdac_1.x6[4].x1.x9.A single_10b_cdac_1.x6[4].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4503 a_25778_31002# single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4504 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4505 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4506 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4507 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4508 single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.cdac_sw_2_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4509 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4510 a_21094_25713# single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[6] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4511 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4512 VSREF SWN_IN[8] a_27534_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4513 single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.cdac_sw_8_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4514 single_10b_cdac_1.x4[2].x3.ck single_10b_cdac_1.x4[2].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4515 VDREF SWP_IN[6] a_12898_34218# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4516 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4517 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4518 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x3.ckb a_7336_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4519 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4520 single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4521 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4522 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4523 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4524 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4525 single_10b_cdac_1.cdac_sw_1_2.x3.ck single_10b_cdac_1.cdac_sw_1_2.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4526 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4527 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4528 VSREF single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4529 VDREF single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4530 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4531 single_10b_cdac_0.x10[8].x2.swn single_10b_cdac_0.x10[8].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4532 single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4533 single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4534 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4535 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4536 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4537 single_10b_cdac_0.cdac_sw_16_0.x1.x7.A single_10b_cdac_0.cdac_sw_16_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4538 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x8.A single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4539 VDREF single_10b_cdac_1.x6[4].x1.x4.A single_10b_cdac_1.x6[4].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4540 VSREF single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4541 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x9.A single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4542 single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4543 single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4544 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4545 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4546 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4547 VSREF single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4548 single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4549 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4550 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4551 VDREF single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4552 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4553 VDREF single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4554 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4555 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x9.A single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4556 single_10b_cdac_0.cdac_sw_1_1.x3.ck single_10b_cdac_0.cdac_sw_1_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4557 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4558 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4559 single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.cdac_sw_8_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4560 VDREF single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4561 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4562 single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4563 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4564 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4565 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4566 single_10b_cdac_0.cdac_sw_1_1.x1.x8.A single_10b_cdac_0.cdac_sw_1_1.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4567 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4568 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4569 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4570 single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4571 VDREF SWP_IN[2] a_59372_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4572 single_10b_cdac_1.x3[1].x2.swn single_10b_cdac_1.x3[1].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4573 a_58494_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4574 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4575 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4576 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4577 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4578 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4579 VSREF single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4580 single_10b_cdac_1.x10b_cap_array_0.SW[8] single_10b_cdac_1.cdac_sw_1_1.x3.ckb a_26656_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4581 VSREF SWN_IN[6] a_54688_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4582 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4583 single_10b_cdac_0.x4[3].x2.swn single_10b_cdac_0.x4[3].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4584 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4585 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x8.A single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4586 VSREF single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4587 VSREF SWN_IN[5] a_51468_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4588 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4589 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4590 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4591 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4592 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4593 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4594 VDREF CF[5] single_10b_cdac_1.x6[5].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4595 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4596 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4597 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x8.A single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4598 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4599 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4600 VCM single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4601 single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4602 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4603 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4604 VDREF single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4605 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4606 VSREF single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4607 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4608 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4609 a_52054_34009# SWP_IN[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4610 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4611 single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.cdac_sw_4_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4612 single_10b_cdac_0.cdac_sw_1_1.x1.x4.A single_10b_cdac_0.cdac_sw_1_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4613 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4614 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4615 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4616 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4617 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4618 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4619 VDREF single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4620 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4621 VDREF single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4622 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4623 single_10b_cdac_1.cdac_sw_4_1.x1.x6.A single_10b_cdac_1.cdac_sw_4_1.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4624 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4625 single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4626 VDREF single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4627 single_10b_cdac_0.cdac_sw_1_2.x3.ck single_10b_cdac_0.cdac_sw_1_2.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4628 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4629 single_10b_cdac_1.x10[8].x2.swn single_10b_cdac_1.x10[8].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4630 single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4631 VSREF single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4632 a_21680_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4633 VDREF single_10b_cdac_0.x6[4].x1.x5.A single_10b_cdac_0.x6[4].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4634 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4635 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4636 single_10b_cdac_0.cdac_sw_4_1.x1.x9.A single_10b_cdac_0.cdac_sw_4_1.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4637 VSREF CF[0] single_10b_cdac_1.x3[0].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4638 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4639 a_52932_33146# single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4640 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4641 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4642 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4643 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4644 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4645 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4646 single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4647 VDREF single_10b_cdac_1.x3[1].x1.x5.A single_10b_cdac_1.x3[1].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4648 VSREF single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4649 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4650 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4651 single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.cdac_sw_8_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4652 VDREF single_10b_cdac_0.x8[7].x1.x8.A single_10b_cdac_0.x8[7].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4653 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4654 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4655 VSREF single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4656 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4657 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4658 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4659 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4660 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4661 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4662 VCM single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4663 VDREF single_10b_cdac_0.x4[2].x1.x3.Y single_10b_cdac_0.x4[2].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4664 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4665 single_10b_cdac_1.cdac_sw_1_1.x2.swn single_10b_cdac_1.cdac_sw_1_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4666 single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4667 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4668 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4669 VDREF single_10b_cdac_1.x6[4].x1.x8.A single_10b_cdac_1.x6[4].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4670 single_10b_cdac_0.x3[1].x2.swn single_10b_cdac_0.x3[1].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4671 VSREF single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4672 single_10b_cdac_0.x6[5].x2.swn single_10b_cdac_0.x6[5].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4673 VDREF single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4674 single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4675 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4676 VSREF single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4677 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4678 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4679 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4680 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4681 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4682 VSREF single_10b_cdac_0.x4[3].x1.x8.A single_10b_cdac_0.x4[3].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4683 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4684 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4685 single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.cdac_sw_2_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4686 single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4687 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4688 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4689 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4690 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4691 VSREF single_10b_cdac_1.x10[8].x1.x8.A single_10b_cdac_1.x10[8].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4692 VSREF single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4693 single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4694 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x3.ck a_55274_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4695 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4696 single_10b_cdac_1.x10b_cap_array_0.SW[4] single_10b_cdac_1.cdac_sw_4_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4697 VCN single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4698 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4699 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x9.A single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4700 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4701 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4702 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4703 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4704 VDREF single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4705 a_37803_24944# single_10b_cdac_0.x2[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4706 VDREF single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4707 VSREF single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4708 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4709 VDREF single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4710 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x8.A single_10b_cdac_0.cdac_sw_4_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4711 VCN single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4712 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4713 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4714 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4715 VSREF single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4716 VSREF single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4717 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4718 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4719 single_10b_cdac_0.x6[5].x2.swn single_10b_cdac_0.x6[5].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4720 VCM single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4721 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4722 single_10b_cdac_1.x8[7].x2.swn single_10b_cdac_1.x8[7].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4723 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4724 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4725 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4726 single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4727 VCN single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4728 single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x2[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4729 VSREF SWN_IN[3] a_11434_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4730 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4731 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4732 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4733 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4734 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4735 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4736 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4737 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4738 single_10b_cdac_0.cdac_sw_8_0.x1.x3.Y CF[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4739 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4740 single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4741 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4742 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4743 VDREF single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4744 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4745 single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4746 single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4747 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4748 VDREF single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4749 VDREF single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4750 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4751 VCM single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4752 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4753 VDREF CF[6] single_10b_cdac_0.cdac_sw_2_1.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4754 single_10b_cdac_0.x8[6].x3.ck single_10b_cdac_0.x8[6].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4755 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4756 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4757 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4758 single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4759 a_20216_25722# SWN_IN[6] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4760 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4761 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4762 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4763 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4764 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4765 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4766 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4767 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4768 VDREF single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4769 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4770 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4771 single_10b_cdac_0.x3[0].x2.swn single_10b_cdac_0.x3[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4772 single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4773 VSREF single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4774 VDREF single_10b_cdac_1.x8[7].x1.x8.A single_10b_cdac_1.x8[7].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4775 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4776 single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.cdac_sw_16_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4777 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4778 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4779 VDREF single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4780 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4781 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4782 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4783 single_10b_cdac_0.x4[2].x3.ck single_10b_cdac_0.x4[2].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4784 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4785 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4786 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4787 VSREF single_10b_cdac_0.x6[5].x1.x8.A single_10b_cdac_0.x6[5].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4788 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4789 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4790 single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4791 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4792 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4793 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4794 VDREF single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4795 single_10b_cdac_1.cdac_sw_1_0.x1.x4.A CF[9] a_29969_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4796 single_10b_cdac_1.x8[6].x2.swn single_10b_cdac_1.x8[6].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4797 single_10b_cdac_0.x4[2].x1.x4.A CF[2] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4798 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4799 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4800 VSREF single_10b_cdac_0.x4[2].x1.x5.A single_10b_cdac_0.x4[2].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4801 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4802 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x3.ckb a_10556_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4803 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4804 single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4805 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4806 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4807 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4808 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4809 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4810 single_10b_cdac_1.cdac_sw_2_1.x1.x8.A single_10b_cdac_1.cdac_sw_2_1.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4811 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4812 VSREF single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4813 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4814 single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4815 VSREF single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4816 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4817 VSREF single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4818 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4819 single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.cdac_sw_16_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4820 VDREF single_10b_cdac_1.x4[3].x1.x9.A single_10b_cdac_1.x4[3].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4821 VDREF single_10b_cdac_0.x3[0].x1.x8.A single_10b_cdac_0.x3[0].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4822 single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4823 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4824 VDREF single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4825 single_10b_cdac_1.cdac_sw_1_0.x1.x3.Y CF[9] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4826 VDREF single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4827 VSREF SWN_IN[2] a_8214_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4828 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4829 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4830 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4831 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4832 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4833 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4834 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4835 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4836 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4837 single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4838 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4839 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4840 single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4841 VCP single_10b_cdac_0.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4842 VCP single_10b_cdac_0.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4843 single_10b_cdac_1.cdac_sw_1_0.x2.swn single_10b_cdac_1.cdac_sw_1_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4844 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4845 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4846 single_10b_cdac_1.cdac_sw_2_1.x1.x4.A single_10b_cdac_1.cdac_sw_2_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4847 a_3377_36566# single_10b_cdac_1.cdac_sw_1_2.x1.x8.A single_10b_cdac_1.cdac_sw_1_2.x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4848 VCM single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4849 VDREF single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4850 single_10b_cdac_0.x3[0].x3.ck single_10b_cdac_0.x3[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4851 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4852 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4853 single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4854 single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4855 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4856 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4857 VDREF single_10b_cdac_1.x4[3].x1.x6.A single_10b_cdac_1.x4[3].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4858 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4859 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4860 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4861 VSREF single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4862 single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4863 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x3.ckb a_10556_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4864 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4865 VDREF single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4866 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4867 single_10b_cdac_0.x10b_cap_array_0.SW[6] single_10b_cdac_0.cdac_sw_2_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4868 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4869 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4870 single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4871 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4872 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4873 single_10b_cdac_0.x4[2].x2.swn single_10b_cdac_0.x4[2].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4874 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4875 VSREF single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4876 single_10b_cdac_1.cdac_sw_2_0.x1.x5.A single_10b_cdac_1.cdac_sw_2_0.x1.x8.A a_23529_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4877 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x9.A single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4878 VDREF single_10b_cdac_1.x8[6].x1.x5.A single_10b_cdac_1.x8[6].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4879 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4880 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4881 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4882 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4883 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4884 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4885 single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4886 single_10b_cdac_1.x6[5].dac_out single_10b_cdac_1.x6[5].x3.ck a_15240_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4887 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4888 a_12898_34218# single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4889 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4890 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4891 single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.cdac_sw_4_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4892 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4893 VDREF single_10b_cdac_0.x8[7].x1.x3.Y single_10b_cdac_0.x8[7].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4894 single_10b_cdac_1.cdac_sw_1_2.x2.swn single_10b_cdac_1.cdac_sw_1_2.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4895 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4896 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4897 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4898 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4899 single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.cdac_sw_8_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4900 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4901 a_56152_31002# single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4902 single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4903 a_60250_25722# SWN_IN[8] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4904 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4905 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4906 single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4907 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4908 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x9.A single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4909 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4910 single_10b_cdac_0.cdac_sw_16_0.x1.x8.A single_10b_cdac_0.cdac_sw_16_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4911 single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4912 single_10b_cdac_1.x6[5].dac_out single_10b_cdac_1.x6[5].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4913 VSREF single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4914 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4915 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4916 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4917 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4918 single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4919 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4920 single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.cdac_sw_8_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4921 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4922 single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4923 a_41808_25713# single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4924 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4925 VDREF single_10b_cdac_1.x2[0].x1.x8.A single_10b_cdac_1.x2[0].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4926 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4927 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4928 single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4929 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4930 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4931 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4932 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4933 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x9.A single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4934 VSREF single_10b_cdac_1.x6[5].x1.x8.A single_10b_cdac_1.x6[5].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4935 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4936 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4937 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4938 VDREF single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4939 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4940 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4941 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4942 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4943 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4944 single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4945 VDREF single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4946 a_46631_36566# single_10b_cdac_0.x8[6].x1.x8.A single_10b_cdac_0.x8[6].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4947 a_14654_25713# single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4948 VSREF single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4949 VCM single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4950 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4951 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4952 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4953 a_11434_25713# single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4954 single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.cdac_sw_2_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4955 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4956 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4957 VDREF single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4958 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4959 VDREF SWP_IN[6] a_46492_34218# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4960 single_10b_cdac_0.cdac_sw_4_0.x1.x8.A single_10b_cdac_0.cdac_sw_4_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4961 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4962 single_10b_cdac_1.cdac_sw_16_0.x1.x5.A single_10b_cdac_1.cdac_sw_16_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4963 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4964 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4965 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4966 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4967 single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4968 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4969 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x8.A single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4970 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4971 single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4972 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x9.A single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4973 VSREF single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4974 single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4975 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4976 single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.cdac_sw_2_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4977 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4978 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x5.A single_10b_cdac_1.cdac_sw_1_2.x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4979 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4980 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4981 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4982 single_10b_cdac_1.cdac_sw_1_1.x1.x9.A single_10b_cdac_1.cdac_sw_1_1.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4983 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4984 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4985 a_3238_34754# single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4986 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4987 single_10b_cdac_1.cdac_sw_1_1.x3.ck single_10b_cdac_1.cdac_sw_1_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4988 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4989 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4990 VDREF single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4991 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4992 single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.cdac_sw_2_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4993 a_59372_31002# single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4994 VDREF single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4995 VDREF single_10b_cdac_1.x4[3].x1.x8.A single_10b_cdac_1.x4[3].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4996 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4997 VSREF single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4998 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4999 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5000 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5001 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5002 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5003 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5004 VSREF SWN_IN[4] a_48248_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5005 single_10b_cdac_0.x8[7].x3.ck single_10b_cdac_0.x8[7].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5006 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x8.A single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5007 single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5008 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5009 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5010 VSREF SWN_IN[3] a_45028_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5011 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5012 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x8.A single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5013 single_10b_cdac_1.cdac_sw_8_0.x1.x7.A single_10b_cdac_1.cdac_sw_8_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5014 single_10b_cdac_0.x8[7].x1.x4.A CF[7] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5015 single_10b_cdac_0.x6[5].dac_out single_10b_cdac_0.x6[5].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5016 VSREF single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5017 VSREF single_10b_cdac_0.x8[7].x1.x5.A single_10b_cdac_0.x8[7].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5018 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5019 single_10b_cdac_0.cdac_sw_1_0.x1.x3.Y CF[9] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5020 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5021 single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5022 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5023 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5024 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5025 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5026 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5027 a_45614_34645# SWP_IN[6] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5028 single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5029 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5030 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5031 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5032 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5033 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5034 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5035 a_24900_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5036 single_10b_cdac_1.cdac_sw_4_1.x1.x3.Y CF[4] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5037 a_56291_35702# CF[3] single_10b_cdac_0.x4[3].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5038 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5039 VDREF single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5040 VDREF SWP_IN[5] a_49712_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5041 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5042 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5043 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5044 single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5045 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5046 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5047 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5048 single_10b_cdac_1.x3[1].x2.swn single_10b_cdac_1.x3[1].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5049 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5050 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5051 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5052 single_10b_cdac_0.cdac_sw_4_1.x1.x6.A single_10b_cdac_0.cdac_sw_4_1.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5053 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5054 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x8.A single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5055 single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5056 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5057 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5058 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5059 a_15240_34009# SWP_IN[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5060 single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5061 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5062 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5063 VSREF CF[2] single_10b_cdac_1.x4[2].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5064 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5065 single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.cdac_sw_4_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5066 single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5067 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5068 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5069 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5070 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5071 single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5072 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5073 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5074 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5075 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5076 single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5077 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5078 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5079 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5080 VSREF single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5081 single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5082 VDREF single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5083 VCM single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5084 single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5085 single_10b_cdac_0.x8[7].x2.swn single_10b_cdac_0.x8[7].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5086 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5087 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5088 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5089 VSREF single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5090 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5091 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5092 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5093 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5094 VSREF single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5095 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5096 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5097 VDREF single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5098 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5099 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5100 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5101 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5102 single_10b_cdac_1.cdac_sw_8_1.x1.x7.A single_10b_cdac_1.cdac_sw_8_1.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5103 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x9.A single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5104 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5105 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5106 single_10b_cdac_1.x6[4].x2.swn single_10b_cdac_1.x6[4].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5107 single_10b_cdac_0.x3[1].x1.x4.A CF[1] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5108 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5109 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5110 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5111 single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5112 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5113 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5114 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5115 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5116 VSREF single_10b_cdac_0.x10[8].x1.x7.A single_10b_cdac_0.x10[8].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5117 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5118 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5119 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5120 single_10b_cdac_0.x6[5].dac_out single_10b_cdac_0.x6[5].x3.ck a_48834_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5121 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5122 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5123 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5124 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5125 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5126 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5127 single_10b_cdac_0.cdac_sw_8_0.x1.x4.A CF[3] a_44243_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5128 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5129 single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5130 VSREF single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5131 single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5132 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5133 VCN single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5134 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5135 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5136 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5137 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5138 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x3.ckb a_7336_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5139 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5140 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5141 VCM single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5142 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5143 VSREF single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5144 single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5145 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5146 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5147 single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5148 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5149 single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5150 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5151 single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5152 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5153 a_63563_24080# single_10b_cdac_0.cdac_sw_1_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5154 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5155 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5156 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5157 a_44150_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5158 a_49712_33146# single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5159 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5160 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5161 single_10b_cdac_0.x2[0].x1.x3.Y CF[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5162 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5163 VSREF single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5164 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5165 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5166 single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5167 VDREF single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5168 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5169 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5170 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5171 VDREF CF[4] single_10b_cdac_0.cdac_sw_4_1.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5172 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5173 VCP single_10b_cdac_1.x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5174 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5175 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5176 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5177 VDREF single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5178 VDREF single_10b_cdac_1.x2[0].x1.x8.A single_10b_cdac_1.x2[0].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5179 VSREF single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5180 single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5181 VDREF single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5182 single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x2[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5183 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5184 single_10b_cdac_1.x8[7].x3.ck single_10b_cdac_1.x8[7].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5185 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5186 single_10b_cdac_1.cdac_sw_8_0.x1.x9.A single_10b_cdac_1.cdac_sw_8_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5187 single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5188 single_10b_cdac_0.x4[2].x2.swn single_10b_cdac_0.x4[2].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5189 single_10b_cdac_0.x6[4].x3.ck single_10b_cdac_0.x6[4].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5190 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5191 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5192 single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.cdac_sw_2_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5193 VSREF single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5194 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x9.A single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5195 VDREF single_10b_cdac_0.x8[6].x1.x9.A single_10b_cdac_0.x8[6].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5196 VSREF single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5197 single_10b_cdac_0.x10b_cap_array_0.SW[6] single_10b_cdac_0.cdac_sw_2_1.x3.ckb a_53810_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5198 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5199 single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5200 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5201 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5202 single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.cdac_sw_8_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5203 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5204 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5205 single_10b_cdac_1.x8[7].x2.swn single_10b_cdac_1.x8[7].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5206 single_10b_cdac_1.x10b_cap_array_0.SW[5] single_10b_cdac_1.cdac_sw_4_0.x3.ckb a_16996_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5207 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5208 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5209 single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5210 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5211 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5212 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5213 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5214 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5215 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5216 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5217 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x3.ck a_24900_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5218 single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.cdac_sw_2_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5219 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5220 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5221 single_10b_cdac_1.x3[1].x3.ck single_10b_cdac_1.x3[1].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5222 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5223 VDREF CF[2] single_10b_cdac_1.cdac_sw_8_1.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5224 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5225 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5226 single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.cdac_sw_4_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5227 single_10b_cdac_0.cdac_sw_1_0.x1.x4.A CF[9] a_63563_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5228 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5229 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5230 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5231 single_10b_cdac_1.cdac_sw_4_1.x1.x8.A single_10b_cdac_1.cdac_sw_4_1.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5232 single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5233 single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5234 single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5235 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5236 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5237 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5238 single_10b_cdac_0.x10[8].x3.ck single_10b_cdac_0.x10[8].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5239 VSREF single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5240 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5241 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5242 VDREF single_10b_cdac_1.x6[5].x1.x9.A single_10b_cdac_1.x6[5].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5243 single_10b_cdac_1.cdac_sw_1_1.x2.swn single_10b_cdac_1.cdac_sw_1_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5244 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5245 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5246 VSREF single_10b_cdac_0.x3[1].x1.x9.A single_10b_cdac_0.x3[1].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5247 VDREF single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5248 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5249 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5250 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5251 VDREF single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5252 a_47370_25722# SWN_IN[4] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5253 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5254 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5255 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5256 single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5257 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5258 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5259 a_40191_35702# CF[8] single_10b_cdac_0.x10[8].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5260 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5261 single_10b_cdac_1.x4[3].x2.swn single_10b_cdac_1.x4[3].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5262 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5263 VSREF single_10b_cdac_1.x8[7].x1.x4.A single_10b_cdac_1.x8[7].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5264 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5265 single_10b_cdac_1.x8[6].x2.swn single_10b_cdac_1.x8[6].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5266 VDREF single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5267 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5268 single_10b_cdac_0.cdac_sw_1_0.x2.swn single_10b_cdac_0.cdac_sw_1_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5269 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5270 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5271 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5272 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5273 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5274 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5275 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5276 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5277 single_10b_cdac_1.cdac_sw_1_0.x1.x8.A single_10b_cdac_1.cdac_sw_1_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5278 single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5279 VSREF single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5280 VSREF CF[7] single_10b_cdac_1.x8[7].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5281 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5282 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5283 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5284 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5285 single_10b_cdac_1.cdac_sw_1_0.x1.x7.A single_10b_cdac_1.cdac_sw_1_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5286 single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5287 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5288 VDREF single_10b_cdac_0.x4[3].x1.x6.A single_10b_cdac_0.x4[3].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5289 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5290 VSREF single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5291 single_10b_cdac_0.x10b_cap_array_0.SW[4] single_10b_cdac_0.cdac_sw_4_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5292 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5293 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5294 single_10b_cdac_1.cdac_sw_4_0.x1.x5.A single_10b_cdac_1.cdac_sw_4_0.x1.x8.A a_17089_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5295 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x9.A single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5296 VSREF single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5297 single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.cdac_sw_16_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5298 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5299 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5300 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5301 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5302 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5303 VDREF CF[1] single_10b_cdac_0.x3[1].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5304 single_10b_cdac_1.cdac_sw_1_1.x3.ck single_10b_cdac_1.cdac_sw_1_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5305 single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5306 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5307 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x3.Y single_10b_cdac_0.cdac_sw_1_2.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5308 single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5309 VDREF single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5310 single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5311 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5312 single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5313 VDREF single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5314 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5315 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5316 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5317 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5318 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5319 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5320 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5321 VCM single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5322 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5323 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5324 VSREF single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5325 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5326 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5327 single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5328 VDREF single_10b_cdac_0.x10[8].x1.x4.A single_10b_cdac_0.x10[8].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5329 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5330 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x3.ck a_58494_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5331 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5332 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5333 a_57030_25722# SWN_IN[7] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5334 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5335 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5336 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5337 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5338 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5339 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5340 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x8.A single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5341 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5342 single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5343 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5344 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5345 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5346 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5347 single_10b_cdac_1.x6[4].dac_out single_10b_cdac_1.x6[4].x3.ck a_18460_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5348 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5349 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5350 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5351 single_10b_cdac_1.x4[3].x1.x4.A CF[3] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5352 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5353 VDREF single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5354 VSREF single_10b_cdac_1.x4[3].x1.x5.A single_10b_cdac_1.x4[3].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5355 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5356 VSREF SWN_IN[2] a_41808_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5357 VDREF single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5358 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5359 VDREF single_10b_cdac_1.x4[2].x1.x3.Y single_10b_cdac_1.x4[2].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5360 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5361 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5362 single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5363 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5364 VSREF single_10b_cdac_0.x6[4].x1.x3.Y a_53071_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5365 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5366 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5367 a_50590_25722# SWN_IN[5] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5368 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5369 single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.cdac_sw_4_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5370 VCM single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5371 single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5372 VDREF single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5373 single_10b_cdac_1.x6[5].x2.swn single_10b_cdac_1.x6[5].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5374 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5375 single_10b_cdac_0.x6[5].x3.ck single_10b_cdac_0.x6[5].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5376 VDREF single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5377 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5378 single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x2[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5379 VSREF single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5380 single_10b_cdac_1.x3[0].x3.ck single_10b_cdac_1.x3[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5381 single_10b_cdac_0.cdac_sw_2_1.x1.x5.A single_10b_cdac_0.cdac_sw_2_1.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5382 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5383 a_45028_25713# single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5384 single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5385 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5386 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5387 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5388 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5389 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5390 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5391 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5392 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5393 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5394 single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5395 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5396 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5397 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5398 VSREF single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5399 single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5400 VDREF single_10b_cdac_1.x4[2].x1.x7.A single_10b_cdac_1.x4[2].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5401 VDREF single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5402 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5403 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5404 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5405 a_23529_24080# single_10b_cdac_1.cdac_sw_2_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5406 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5407 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5408 single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5409 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5410 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5411 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5412 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5413 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5414 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5415 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5416 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5417 single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5418 single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5419 single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5420 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5421 single_10b_cdac_0.cdac_sw_2_1.x1.x7.A single_10b_cdac_0.cdac_sw_2_1.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5422 VDREF single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5423 VDREF single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5424 VSREF single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5425 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5426 single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5427 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5428 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5429 single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5430 VDREF single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5431 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5432 VSREF single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5433 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5434 single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5435 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5436 VSREF single_10b_cdac_0.x3[1].x1.x10.A single_10b_cdac_0.x3[1].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5437 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5438 VDREF single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5439 single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5440 VSREF single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5441 single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.cdac_sw_8_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5442 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5443 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5444 single_10b_cdac_1.x8[6].x3.ck single_10b_cdac_1.x8[6].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5445 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5446 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5447 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5448 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5449 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5450 VDREF single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5451 single_10b_cdac_0.x10b_cap_array_0.SW[5] single_10b_cdac_0.cdac_sw_4_0.x3.ckb a_50590_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5452 VSREF single_10b_cdac_1.x3[0].x1.x4.A single_10b_cdac_1.x3[0].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5453 single_10b_cdac_0.x2[0].x1.x9.A single_10b_cdac_0.x2[0].x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5454 single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5455 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5456 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5457 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5458 VSREF single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5459 single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.cdac_sw_8_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5460 VDREF single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5461 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5462 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5463 single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5464 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5465 single_10b_cdac_1.x4[2].x3.ck single_10b_cdac_1.x4[2].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5466 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5467 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5468 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5469 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5470 VSREF single_10b_cdac_1.cdac_sw_1_2.x1.x7.A single_10b_cdac_1.cdac_sw_1_2.x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5471 single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5472 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x8.A single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5473 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5474 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5475 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5476 single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.cdac_sw_8_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5477 VSREF single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5478 single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5479 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5480 VSREF single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5481 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5482 single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5483 a_48834_34009# SWP_IN[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5484 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5485 a_54688_25713# single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[6] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5486 VSREF CF[2] single_10b_cdac_0.x4[2].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5487 single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5488 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5489 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5490 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5491 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5492 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5493 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5494 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5495 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5496 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5497 VSREF single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5498 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5499 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5500 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5501 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5502 VDREF SWP_IN[4] a_52932_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5503 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5504 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5505 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5506 single_10b_cdac_1.x10b_cap_array_0.SW[6] single_10b_cdac_1.cdac_sw_2_1.x3.ckb a_20216_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5507 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5508 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5509 VCP single_10b_cdac_1.x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5510 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5511 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5512 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5513 VSREF single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5514 single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5515 single_10b_cdac_0.cdac_sw_1_1.x3.ck single_10b_cdac_0.cdac_sw_1_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5516 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5517 VDREF single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5518 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5519 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5520 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5521 single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.cdac_sw_4_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5522 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x9.A single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5523 a_22558_31002# single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5524 single_10b_cdac_1.cdac_sw_1_2.x3.ck single_10b_cdac_1.cdac_sw_1_2.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5525 VSREF single_10b_cdac_0.x6[4].x1.x6.A single_10b_cdac_0.x6[4].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5526 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5527 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5528 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5529 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5530 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5531 a_40930_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5532 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5533 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5534 single_10b_cdac_1.x10b_cap_array_0.SW[6] single_10b_cdac_1.cdac_sw_2_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5535 single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5536 single_10b_cdac_0.x8[7].x3.ck single_10b_cdac_0.x8[7].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5537 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x8.A single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5538 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5539 VSREF single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5540 single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5541 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5542 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5543 single_10b_cdac_1.x8[6].dac_out single_10b_cdac_1.x8[6].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5544 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5545 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5546 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5547 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5548 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5549 a_16996_25722# SWN_IN[5] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5550 single_10b_cdac_1.x6[4].x3.ck single_10b_cdac_1.x6[4].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5551 VCM single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5552 VDREF single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5553 single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5554 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5555 single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5556 VCP single_10b_cdac_0.x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5557 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5558 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5559 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x9.A single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5560 VDREF single_10b_cdac_0.x6[4].x1.x9.A single_10b_cdac_0.x6[4].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5561 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x4.A single_10b_cdac_0.cdac_sw_1_2.x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5562 single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5563 single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5564 VSREF single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5565 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5566 VDREF single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5567 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5568 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5569 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5570 VDREF single_10b_cdac_1.x3[1].x1.x9.A single_10b_cdac_1.x3[1].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5571 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5572 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5573 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5574 single_10b_cdac_0.cdac_sw_1_0.x2.swn single_10b_cdac_0.cdac_sw_1_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5575 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5576 VDREF SWP_IN[3] a_56152_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5577 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x8.A single_10b_cdac_1.cdac_sw_1_1.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5578 single_10b_cdac_0.cdac_sw_1_2.x2.swn single_10b_cdac_0.cdac_sw_1_2.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5579 single_10b_cdac_0.x6[4].x2.swn single_10b_cdac_0.x6[4].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5580 VSREF single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5581 single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5582 VDREF single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5583 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5584 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5585 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5586 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5587 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5588 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5589 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5590 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5591 single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.cdac_sw_4_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5592 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5593 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5594 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5595 VDREF single_10b_cdac_0.x10[8].x1.x9.A single_10b_cdac_0.x10[8].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5596 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5597 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5598 single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5599 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5600 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5601 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x9.A single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5602 single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5603 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5604 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5605 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5606 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5607 single_10b_cdac_0.cdac_sw_8_1.x1.x4.A single_10b_cdac_0.cdac_sw_8_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5608 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5609 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5610 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5611 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5612 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5613 single_10b_cdac_0.x3[0].x1.x5.A single_10b_cdac_0.x3[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5614 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5615 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5616 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5617 VDREF single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5618 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x8.A single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5619 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5620 single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.cdac_sw_2_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5621 single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5622 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5623 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5624 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5625 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5626 a_7336_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5627 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5628 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5629 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5630 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5631 VDREF single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5632 VSREF single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5633 single_10b_cdac_1.x8[7].x3.ck single_10b_cdac_1.x8[7].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5634 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5635 VSREF single_10b_cdac_0.x4[3].x1.x9.A single_10b_cdac_0.x4[3].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5636 single_10b_cdac_1.x2[0].x1.x9.A single_10b_cdac_1.x2[0].x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5637 single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.cdac_sw_2_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5638 VDREF single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5639 single_10b_cdac_1.x8[6].dac_out single_10b_cdac_1.x8[6].x3.ck a_12020_34645# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5640 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5641 single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5642 VDREF single_10b_cdac_0.x6[5].x1.x9.A single_10b_cdac_0.x6[5].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5643 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5644 VSREF single_10b_cdac_1.x10[8].x1.x9.A single_10b_cdac_1.x10[8].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5645 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5646 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5647 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5648 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5649 VDREF single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5650 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5651 single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5652 VSREF SWN_IN[4] a_14654_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5653 single_10b_cdac_0.cdac_sw_1_2.dac_out single_10b_cdac_0.cdac_sw_1_2.x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5654 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5655 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5656 VSREF SWN_IN[3] a_11434_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5657 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5658 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5659 single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.cdac_sw_2_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5660 VSREF single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5661 VDREF single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5662 single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5663 single_10b_cdac_1.x3[1].x3.ck single_10b_cdac_1.x3[1].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5664 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5665 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5666 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5667 single_10b_cdac_1.x2[0].x1.x5.A single_10b_cdac_1.x2[0].x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5668 single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5669 VSREF single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5670 VCM single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5671 VDREF single_10b_cdac_0.x6[5].x1.x6.A single_10b_cdac_0.x6[5].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5672 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5673 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5674 single_10b_cdac_1.cdac_sw_8_1.x1.x8.A single_10b_cdac_1.cdac_sw_8_1.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5675 VSREF single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5676 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5677 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5678 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5679 VDREF single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5680 VSREF single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5681 single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5682 VSREF CF[7] single_10b_cdac_0.x8[7].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5683 a_12020_34645# SWP_IN[6] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5684 VSREF single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5685 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5686 single_10b_cdac_0.cdac_sw_1_0.x1.x7.A single_10b_cdac_0.cdac_sw_1_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5687 single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5688 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5689 VDREF single_10b_cdac_1.x8[7].x1.x9.A single_10b_cdac_1.x8[7].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5690 VDREF single_10b_cdac_0.x3[1].x1.x5.A single_10b_cdac_0.x3[1].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5691 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5692 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5693 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5694 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5695 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5696 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5697 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5698 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5699 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5700 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5701 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5702 VDREF single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5703 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5704 VDREF SWP_IN[9] a_3238_34754# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5705 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5706 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5707 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5708 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5709 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5710 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5711 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5712 VDREF single_10b_cdac_0.x6[4].x1.x8.A single_10b_cdac_0.x6[4].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5713 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5714 VDREF single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5715 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5716 single_10b_cdac_1.cdac_sw_8_1.x1.x4.A single_10b_cdac_1.cdac_sw_8_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5717 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5718 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5719 VSREF single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5720 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5721 single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.cdac_sw_4_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5722 single_10b_cdac_1.cdac_sw_1_1.x1.x6.A single_10b_cdac_1.cdac_sw_1_1.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5723 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5724 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5725 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5726 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5727 VDREF single_10b_cdac_1.x8[7].x1.x6.A single_10b_cdac_1.x8[7].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5728 VSREF single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5729 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5730 single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5731 VSREF CF[9] single_10b_cdac_1.cdac_sw_1_2.x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5732 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5733 VSREF single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5734 a_59372_31002# single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5735 single_10b_cdac_0.x4[2].x2.swn single_10b_cdac_0.x4[2].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5736 single_10b_cdac_1.x6[5].x1.x4.A CF[5] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5737 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5738 VSREF single_10b_cdac_0.x6[5].x1.x9.A single_10b_cdac_0.x6[5].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5739 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5740 single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.cdac_sw_2_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5741 single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5742 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5743 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5744 VDREF single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5745 VSREF single_10b_cdac_0.x3[0].x1.x8.A single_10b_cdac_0.x3[0].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5746 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x9.A single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5747 single_10b_cdac_0.x6[4].x3.ck single_10b_cdac_0.x6[4].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5748 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x3.ckb a_40930_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5749 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5750 VDREF single_10b_cdac_1.x6[4].x1.x3.Y single_10b_cdac_1.x6[4].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5751 single_10b_cdac_1.cdac_sw_4_0.x1.x9.A single_10b_cdac_1.cdac_sw_4_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5752 single_10b_cdac_0.x8[6].dac_out single_10b_cdac_0.x8[6].x3.ck a_45614_34645# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5753 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5754 a_44150_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5755 single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5756 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5757 VSREF single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5758 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5759 VDREF SWP_IN[6] a_12898_34218# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5760 VDREF single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5761 VSREF single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5762 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5763 a_29137_35702# CF[1] single_10b_cdac_1.x3[1].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5764 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5765 single_10b_cdac_0.cdac_sw_4_1.x1.x5.A single_10b_cdac_0.cdac_sw_4_1.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5766 single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5767 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x8.A single_10b_cdac_0.cdac_sw_1_1.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5768 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5769 a_10556_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5770 VCN single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5771 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5772 single_10b_cdac_0.x3[0].x3.ck single_10b_cdac_0.x3[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5773 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5774 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5775 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5776 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5777 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5778 VDREF single_10b_cdac_1.x8[6].x1.x9.A single_10b_cdac_1.x8[6].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5779 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5780 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5781 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5782 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5783 VSREF SWN_IN[6] a_21094_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5784 a_17089_24080# single_10b_cdac_1.cdac_sw_4_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5785 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5786 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x8.A single_10b_cdac_1.cdac_sw_8_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5787 single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5788 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5789 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5790 VDREF single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5791 VDREF single_10b_cdac_0.x4[2].x1.x7.A single_10b_cdac_0.x4[2].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5792 VCM single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5793 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5794 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5795 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5796 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5797 VDREF single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5798 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5799 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5800 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5801 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5802 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5803 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5804 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5805 VSREF single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5806 single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5807 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5808 VDREF single_10b_cdac_0.x8[6].x1.x8.A single_10b_cdac_0.x8[6].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5809 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5810 VDREF single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5811 VCN single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5812 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5813 single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x2[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5814 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5815 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5816 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5817 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5818 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5819 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5820 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5821 VSREF single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5822 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5823 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5824 single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5825 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5826 single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.cdac_sw_4_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5827 single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5828 VSREF single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5829 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5830 single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.cdac_sw_16_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5831 VDREF CF[4] single_10b_cdac_1.cdac_sw_4_1.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5832 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5833 VDREF single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5834 VCN VCM sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5835 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x3.ckb a_44150_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5836 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5837 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5838 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5839 VSREF single_10b_cdac_0.x4[2].x1.x8.A single_10b_cdac_0.x4[2].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5840 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5841 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5842 single_10b_cdac_1.x4[2].x1.x5.A single_10b_cdac_1.x4[2].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5843 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x3.ck a_21680_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5844 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5845 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5846 VSREF single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5847 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x8.A single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5848 single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5849 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5850 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5851 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5852 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5853 VSREF single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5854 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5855 single_10b_cdac_1.x6[4].x3.ck single_10b_cdac_1.x6[4].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5856 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5857 VSREF single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5858 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5859 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5860 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5861 single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5862 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5863 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5864 single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5865 VSREF single_10b_cdac_1.x6[5].x1.x9.A single_10b_cdac_1.x6[5].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5866 VDREF single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5867 VDREF single_10b_cdac_1.x3[0].x1.x9.A single_10b_cdac_1.x3[0].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5868 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5869 VSREF single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5870 single_10b_cdac_1.cdac_sw_16_0.x1.x4.A CF[0] a_989_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5871 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5872 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5873 single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.cdac_sw_8_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5874 single_10b_cdac_1.x8[6].x3.ck single_10b_cdac_1.x8[6].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5875 a_52932_33146# single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5876 a_48248_25713# single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5877 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5878 VSREF single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5879 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5880 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5881 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5882 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5883 VCM single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5884 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5885 VDREF single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5886 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5887 single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5888 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5889 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5890 VSREF single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5891 VSREF single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5892 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5893 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5894 single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5895 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5896 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5897 single_10b_cdac_0.cdac_sw_16_0.x1.x5.A single_10b_cdac_0.cdac_sw_16_0.x1.x8.A a_34583_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5898 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5899 single_10b_cdac_1.x4[2].x3.ck single_10b_cdac_1.x4[2].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5900 single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.cdac_sw_2_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5901 single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5902 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5903 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5904 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5905 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5906 single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5907 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5908 single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.cdac_sw_8_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5909 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5910 single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5911 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5912 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5913 single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.cdac_sw_16_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5914 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5915 VDREF single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5916 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x3.ck a_24900_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5917 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5918 single_10b_cdac_1.cdac_sw_1_2.x3.ck single_10b_cdac_1.cdac_sw_1_2.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5919 single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5920 VSREF single_10b_cdac_1.x10[8].x1.x9.A a_6597_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5921 single_10b_cdac_0.x10b_cap_array_0.SW[5] single_10b_cdac_0.cdac_sw_4_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5922 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5923 single_10b_cdac_1.x10b_cap_array_0.SW[4] single_10b_cdac_1.cdac_sw_4_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5924 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5925 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5926 single_10b_cdac_0.cdac_sw_4_0.x1.x6.A single_10b_cdac_0.cdac_sw_4_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5927 single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5928 single_10b_cdac_0.x8[7].x2.swn single_10b_cdac_0.x8[7].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5929 VSREF single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5930 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5931 single_10b_cdac_0.cdac_sw_1_1.x2.swn single_10b_cdac_0.cdac_sw_1_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5932 single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5933 single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5934 single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5935 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5936 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x9.A single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5937 single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5938 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5939 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5940 single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5941 single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5942 a_51468_25713# single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5943 VSREF single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5944 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5945 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5946 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5947 single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x2[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5948 VDREF single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5949 VDREF single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5950 VSREF single_10b_cdac_1.x10[8].x1.x6.A single_10b_cdac_1.x10[8].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5951 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x9.A single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5952 single_10b_cdac_0.cdac_sw_1_1.x3.ck single_10b_cdac_0.cdac_sw_1_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5953 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5954 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5955 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5956 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5957 single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.cdac_sw_16_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5958 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5959 a_13037_35702# CF[6] single_10b_cdac_1.x8[6].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5960 VDREF single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5961 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5962 a_56291_36566# single_10b_cdac_0.x4[3].x1.x8.A single_10b_cdac_0.x4[3].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5963 VSREF single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5964 single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5965 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5966 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5967 VDREF single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5968 single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5969 single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5970 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5971 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5972 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5973 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5974 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5975 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5976 single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5977 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5978 VDREF single_10b_cdac_0.x8[7].x1.x7.A single_10b_cdac_0.x8[7].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5979 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5980 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5981 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5982 VSREF single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5983 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5984 single_10b_cdac_0.x2[0].x1.x7.A single_10b_cdac_0.x2[0].x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5985 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x8.A single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5986 single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5987 single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.cdac_sw_4_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5988 VSREF single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5989 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5990 VCN single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5991 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5992 single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x2[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5993 single_10b_cdac_0.cdac_sw_16_0.x1.x4.A single_10b_cdac_0.cdac_sw_16_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5994 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5995 VDREF single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5996 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5997 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5998 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5999 VCM single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6000 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6001 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6002 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6003 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6004 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6005 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6006 single_10b_cdac_1.x10[8].x2.swn single_10b_cdac_1.x10[8].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6007 single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6008 single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.cdac_sw_4_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6009 VDREF single_10b_cdac_1.x3[0].x1.x8.A single_10b_cdac_1.x3[0].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6010 VSREF single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6011 VSREF single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6012 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6013 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6014 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6015 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6016 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6017 single_10b_cdac_0.cdac_sw_1_0.x1.x8.A single_10b_cdac_0.cdac_sw_1_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6018 single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6019 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6020 VDREF single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6021 VSREF SWN_IN[7] a_57908_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6022 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6023 VSREF single_10b_cdac_0.x8[7].x1.x8.A single_10b_cdac_0.x8[7].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6024 single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6025 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6026 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6027 single_10b_cdac_1.cdac_sw_2_1.x1.x7.A single_10b_cdac_1.cdac_sw_2_1.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6028 single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.cdac_sw_8_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6029 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6030 VDREF single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6031 single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6032 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6033 a_50683_24944# single_10b_cdac_0.cdac_sw_4_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6034 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x9.A single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6035 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6036 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6037 VDREF single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6038 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6039 single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6040 a_55274_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6041 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6042 single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6043 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6044 VCM single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6045 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6046 single_10b_cdac_0.x3[1].x2.swn single_10b_cdac_0.x3[1].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6047 single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6048 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6049 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6050 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6051 single_10b_cdac_0.cdac_sw_1_2.x2.swn single_10b_cdac_0.cdac_sw_1_2.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6052 single_10b_cdac_1.cdac_sw_1_1.x1.x5.A single_10b_cdac_1.cdac_sw_1_1.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6053 single_10b_cdac_1.cdac_sw_2_0.x1.x3.Y CF[7] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6054 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6055 single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6056 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6057 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6058 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6059 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6060 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6061 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6062 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6063 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6064 single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6065 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6066 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6067 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6068 VSREF single_10b_cdac_1.x10[8].x1.x8.A single_10b_cdac_1.x10[8].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6069 single_10b_cdac_0.cdac_sw_2_0.x1.x7.A single_10b_cdac_0.cdac_sw_2_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6070 VSREF single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6071 single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6072 VDREF single_10b_cdac_0.x4[3].x1.x5.A single_10b_cdac_0.x4[3].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6073 VSREF single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6074 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6075 single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6076 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6077 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6078 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6079 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6080 VDREF single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6081 single_10b_cdac_1.x10[8].dac_out single_10b_cdac_1.x10[8].x3.ck a_5580_34963# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6082 VDREF single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6083 a_12898_34218# single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6084 a_56152_31002# single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6085 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6086 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6087 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6088 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6089 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6090 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6091 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6092 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6093 single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6094 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6095 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6096 VDREF single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6097 single_10b_cdac_1.x8[7].x2.swn single_10b_cdac_1.x8[7].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6098 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6099 single_10b_cdac_1.cdac_sw_1_0.x1.x4.A single_10b_cdac_1.cdac_sw_1_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6100 single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x2[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6101 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6102 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6103 single_10b_cdac_0.x6[4].x2.swn single_10b_cdac_0.x6[4].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6104 VCM single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6105 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6106 single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6107 VDREF single_10b_cdac_1.x4[2].x1.x8.A single_10b_cdac_1.x4[2].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6108 VSREF single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6109 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6110 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6111 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6112 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6113 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6114 a_21094_25713# single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[6] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6115 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6116 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6117 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6118 single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.cdac_sw_4_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6119 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6120 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6121 single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6122 single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6123 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6124 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6125 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6126 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6127 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6128 VDREF single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6129 single_10b_cdac_0.x8[6].x3.ck single_10b_cdac_0.x8[6].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6130 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6131 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6132 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6133 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6134 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6135 single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6136 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6137 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6138 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6139 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6140 VDREF single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6141 VCM single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6142 single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6143 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6144 VDREF single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6145 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6146 single_10b_cdac_0.x10[8].x2.swn single_10b_cdac_0.x10[8].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6147 single_10b_cdac_0.x4[3].x2.swn single_10b_cdac_0.x4[3].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6148 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6149 single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6150 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6151 VDREF SWP_IN[6] a_46492_34218# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6152 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6153 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6154 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6155 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6156 single_10b_cdac_0.x4[2].x3.ck single_10b_cdac_0.x4[2].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6157 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6158 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6159 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6160 single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.cdac_sw_4_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6161 single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6162 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6163 VDREF single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6164 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6165 single_10b_cdac_1.x3[0].x2.swn single_10b_cdac_1.x3[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6166 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6167 single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6168 a_40191_36566# single_10b_cdac_0.x10[8].x1.x8.A single_10b_cdac_0.x10[8].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6169 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6170 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6171 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6172 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6173 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6174 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6175 single_10b_cdac_1.x8[7].x1.x4.A CF[7] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6176 single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6177 VSREF single_10b_cdac_1.x8[7].x1.x5.A single_10b_cdac_1.x8[7].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6178 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6179 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6180 a_58494_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6181 a_59372_31002# single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6182 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6183 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6184 VSREF SWN_IN[6] a_54688_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6185 single_10b_cdac_0.cdac_sw_4_1.x1.x3.Y CF[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6186 VSREF single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6187 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6188 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6189 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6190 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6191 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6192 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6193 VSREF single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6194 VDREF CF[7] single_10b_cdac_0.cdac_sw_2_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6195 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6196 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6197 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6198 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6199 single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6200 VDREF single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6201 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x8.A single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6202 VDREF single_10b_cdac_0.x10[8].x1.x8.A single_10b_cdac_0.x10[8].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6203 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6204 single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6205 VSREF single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6206 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6207 VCM single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6208 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6209 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6210 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6211 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6212 single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6213 single_10b_cdac_1.cdac_sw_16_0.x1.x3.Y CF[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6214 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6215 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6216 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6217 single_10b_cdac_1.cdac_sw_1_0.x2.swn single_10b_cdac_1.cdac_sw_1_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6218 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6219 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6220 single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6221 VDREF SWP_IN[3] a_22558_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6222 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6223 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6224 single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6225 VDREF single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6226 single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6227 single_10b_cdac_0.x6[4].dac_out single_10b_cdac_0.x6[4].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6228 single_10b_cdac_0.x10[8].x3.ck single_10b_cdac_0.x10[8].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6229 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6230 single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6231 single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6232 single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6233 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6234 single_10b_cdac_1.x6[5].x2.swn single_10b_cdac_1.x6[5].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6235 single_10b_cdac_1.x6[4].x1.x5.A single_10b_cdac_1.x6[4].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6236 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6237 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6238 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6239 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6240 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6241 single_10b_cdac_1.x10b_cap_array_0.SW[4] single_10b_cdac_1.cdac_sw_4_1.x3.ckb a_13776_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6242 VSREF SWN_IN[2] a_41808_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6243 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6244 single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6245 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6246 a_22558_31002# single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6247 single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6248 single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6249 VDREF SWP_IN[5] a_49712_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6250 single_10b_cdac_1.cdac_sw_2_0.x1.x8.A single_10b_cdac_1.cdac_sw_2_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6251 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x9.A single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6252 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6253 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6254 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6255 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6256 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6257 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6258 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6259 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6260 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6261 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6262 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6263 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6264 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6265 VDREF single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6266 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6267 single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6268 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6269 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6270 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6271 single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6272 VDREF single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6273 single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6274 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6275 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6276 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6277 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6278 VCM single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6279 single_10b_cdac_1.cdac_sw_8_0.x1.x5.A single_10b_cdac_1.cdac_sw_8_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6280 VDREF single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6281 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6282 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6283 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6284 single_10b_cdac_1.x3[0].x2.swn single_10b_cdac_1.x3[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6285 single_10b_cdac_1.x4[3].x2.swn single_10b_cdac_1.x4[3].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6286 VDREF single_10b_cdac_1.x2[0].x1.x8.A single_10b_cdac_1.x2[0].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6287 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6288 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6289 single_10b_cdac_0.cdac_sw_8_1.x1.x7.A single_10b_cdac_0.cdac_sw_8_1.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6290 single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6291 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6292 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6293 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6294 VDREF single_10b_cdac_0.x8[6].x1.x11.A single_10b_cdac_0.x8[6].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6295 VSREF single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6296 VSREF single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6297 single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6298 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6299 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6300 single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6301 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6302 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6303 single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6304 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6305 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6306 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6307 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6308 VSREF single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6309 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6310 VDREF SWP_IN[3] a_56152_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6311 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6312 single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.cdac_sw_2_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6313 VDREF single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6314 single_10b_cdac_1.cdac_sw_4_1.x1.x4.A single_10b_cdac_1.cdac_sw_4_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6315 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6316 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6317 single_10b_cdac_0.x4[3].x3.ck single_10b_cdac_0.x4[3].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6318 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6319 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6320 single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6321 VDREF single_10b_cdac_1.x6[5].x1.x6.A single_10b_cdac_1.x6[5].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6322 single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6323 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6324 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6325 single_10b_cdac_1.cdac_sw_16_0.x1.x8.A single_10b_cdac_1.cdac_sw_16_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6326 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x3.ckb a_40930_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6327 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6328 single_10b_cdac_0.cdac_sw_8_0.x1.x6.A single_10b_cdac_0.cdac_sw_8_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6329 VSREF single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6330 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x8.A single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6331 single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6332 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6333 single_10b_cdac_1.cdac_sw_16_0.x1.x7.A single_10b_cdac_1.cdac_sw_16_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6334 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6335 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6336 single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.cdac_sw_2_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6337 single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6338 single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6339 single_10b_cdac_0.x6[4].dac_out single_10b_cdac_0.x6[4].x3.ck a_52054_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6340 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6341 VSREF single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6342 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6343 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6344 single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6345 VDREF single_10b_cdac_0.x6[5].x1.x4.A single_10b_cdac_0.x6[5].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6346 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6347 single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6348 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x3.ckb a_7336_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6349 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6350 single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6351 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6352 VSREF single_10b_cdac_1.x4[3].x1.x8.A single_10b_cdac_1.x4[3].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6353 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6354 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6355 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6356 VSREF single_10b_cdac_1.x3[1].x1.x6.A single_10b_cdac_1.x3[1].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6357 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6358 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6359 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6360 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6361 VSREF single_10b_cdac_1.x3[0].x1.x5.A single_10b_cdac_1.x3[0].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6362 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6363 a_49712_33146# single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6364 a_53810_25722# SWN_IN[6] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6365 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6366 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6367 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6368 VDREF single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6369 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6370 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6371 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6372 VSREF single_10b_cdac_0.cdac_sw_2_1.x1.x9.A single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6373 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6374 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6375 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6376 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6377 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6378 single_10b_cdac_0.x8[7].x3.ck single_10b_cdac_0.x8[7].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6379 a_41808_25713# single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6380 single_10b_cdac_1.x2[0].x1.x6.A single_10b_cdac_1.x2[0].x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6381 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6382 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6383 single_10b_cdac_1.x4[2].x2.swn single_10b_cdac_1.x4[2].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6384 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6385 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6386 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6387 single_10b_cdac_0.cdac_sw_1_1.x1.x6.A single_10b_cdac_0.cdac_sw_1_1.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6388 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6389 a_29876_25722# SWN_IN[9] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6390 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6391 single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6392 single_10b_cdac_1.x6[5].x2.swn single_10b_cdac_1.x6[5].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6393 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6394 a_24900_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6395 VCM single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6396 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6397 single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6398 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6399 single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6400 single_10b_cdac_0.cdac_sw_1_1.x2.swn single_10b_cdac_0.cdac_sw_1_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6401 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6402 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6403 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x7.A single_10b_cdac_0.cdac_sw_1_2.x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6404 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6405 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6406 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6407 single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6408 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6409 a_11434_25713# single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6410 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6411 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6412 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6413 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6414 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6415 VSREF single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6416 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6417 VDREF single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6418 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6419 VDREF CF[2] single_10b_cdac_0.cdac_sw_8_1.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6420 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6421 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6422 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6423 VDREF single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6424 single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6425 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6426 VDREF single_10b_cdac_0.x3[0].x1.x3.Y single_10b_cdac_0.x3[0].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6427 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6428 single_10b_cdac_0.cdac_sw_8_0.x1.x8.A single_10b_cdac_0.cdac_sw_8_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6429 a_6597_35702# CF[8] single_10b_cdac_1.x10[8].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6430 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6431 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6432 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6433 VDREF single_10b_cdac_1.x4[2].x1.x8.A single_10b_cdac_1.x4[2].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6434 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6435 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6436 single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6437 VSREF single_10b_cdac_0.x2[0].x1.x8.A single_10b_cdac_0.x2[0].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6438 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6439 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6440 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6441 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6442 single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6443 single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.cdac_sw_4_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6444 single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6445 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6446 VSREF single_10b_cdac_0.x6[4].x1.x7.A single_10b_cdac_0.x6[4].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6447 single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6448 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x8.A single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6449 single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6450 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6451 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6452 VDREF single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6453 single_10b_cdac_1.cdac_sw_4_1.x1.x7.A single_10b_cdac_1.cdac_sw_4_1.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6454 VDREF single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6455 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6456 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6457 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6458 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6459 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6460 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6461 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6462 a_44243_24944# single_10b_cdac_0.cdac_sw_8_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6463 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6464 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6465 single_10b_cdac_0.x8[7].x2.swn single_10b_cdac_0.x8[7].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6466 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6467 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6468 VDREF single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6469 single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6470 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6471 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6472 VSREF single_10b_cdac_1.x4[3].x1.x10.A single_10b_cdac_1.x4[3].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6473 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6474 VSREF SWN_IN[3] a_45028_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6475 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6476 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6477 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6478 single_10b_cdac_0.cdac_sw_1_2.x3.ck single_10b_cdac_0.cdac_sw_1_2.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6479 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6480 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6481 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6482 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6483 single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6484 single_10b_cdac_1.x6[4].x2.swn single_10b_cdac_1.x6[4].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6485 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6486 VDREF single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6487 single_10b_cdac_0.cdac_sw_1_2.x1.x4.A CF[9] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6488 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6489 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x3.ckb a_10556_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6490 VSREF single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6491 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x5.A single_10b_cdac_0.cdac_sw_1_2.x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6492 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6493 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6494 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6495 single_10b_cdac_0.cdac_sw_2_0.x1.x3.Y CF[7] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6496 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6497 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6498 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6499 single_10b_cdac_0.cdac_sw_4_0.x1.x3.Y CF[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6500 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6501 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6502 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6503 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6504 single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6505 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6506 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6507 single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.cdac_sw_8_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6508 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6509 a_58494_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6510 VDREF single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6511 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6512 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6513 single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6514 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6515 VSREF single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6516 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6517 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6518 single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6519 a_49851_35702# CF[5] single_10b_cdac_0.x6[5].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6520 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6521 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6522 VSREF single_10b_cdac_0.x3[1].x1.x9.A a_62731_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6523 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6524 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6525 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6526 VDREF single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6527 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6528 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6529 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6530 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6531 single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6532 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6533 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6534 VDREF single_10b_cdac_1.x6[4].x1.x8.A single_10b_cdac_1.x6[4].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6535 VSREF single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6536 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6537 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6538 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6539 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6540 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6541 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6542 a_14654_25713# single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6543 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6544 a_37803_24080# single_10b_cdac_0.x2[0].x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6545 single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6546 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6547 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6548 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6549 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6550 single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6551 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6552 VDREF single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6553 VDREF single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6554 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6555 VSREF single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6556 single_10b_cdac_0.x10[8].x3.ck single_10b_cdac_0.x10[8].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6557 VSREF single_10b_cdac_0.x3[1].x1.x6.A single_10b_cdac_0.x3[1].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6558 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6559 single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.cdac_sw_8_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6560 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6561 single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x2[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6562 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6563 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6564 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6565 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6566 a_50590_25722# SWN_IN[5] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6567 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6568 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6569 single_10b_cdac_0.x6[4].x3.ck single_10b_cdac_0.x6[4].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6570 VSREF single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6571 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6572 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x8.A single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6573 single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6574 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6575 VDREF single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6576 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6577 single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.cdac_sw_8_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6578 VSREF single_10b_cdac_1.x8[6].x1.x6.A single_10b_cdac_1.x8[6].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6579 single_10b_cdac_1.x8[7].x2.swn single_10b_cdac_1.x8[7].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6580 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6581 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6582 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6583 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6584 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6585 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6586 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6587 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6588 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6589 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6590 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6591 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6592 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6593 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6594 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6595 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6596 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6597 single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6598 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6599 VSREF single_10b_cdac_0.x8[6].x1.x4.A single_10b_cdac_0.x8[6].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6600 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6601 single_10b_cdac_1.x3[1].x3.ck single_10b_cdac_1.x3[1].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6602 VSREF single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6603 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6604 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6605 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6606 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6607 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6608 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6609 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6610 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6611 a_13776_25722# SWN_IN[4] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6612 VSREF SWN_IN[4] a_48248_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6613 single_10b_cdac_0.x2[0].x1.x4.A CF[1] a_37803_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6614 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6615 single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.cdac_sw_16_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6616 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6617 single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.cdac_sw_4_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6618 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6619 VCN VCM sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6620 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6621 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6622 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6623 VSREF single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6624 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6625 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6626 single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6627 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6628 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6629 VDREF single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6630 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6631 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6632 VSREF single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6633 single_10b_cdac_0.x3[1].x2.swn single_10b_cdac_0.x3[1].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6634 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6635 VSREF single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6636 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6637 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6638 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6639 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6640 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6641 single_10b_cdac_1.cdac_sw_1_0.x1.x5.A single_10b_cdac_1.cdac_sw_1_0.x1.x8.A a_29969_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6642 VSREF single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6643 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6644 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6645 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6646 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6647 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6648 single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6649 a_8214_25713# single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6650 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6651 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6652 VDREF single_10b_cdac_0.x6[5].x1.x9.A single_10b_cdac_0.x6[5].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6653 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6654 VCP VCM sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6655 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6656 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6657 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6658 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6659 VSREF single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6660 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6661 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6662 single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6663 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6664 VDREF single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6665 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6666 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6667 single_10b_cdac_1.x10[8].x3.ck single_10b_cdac_1.x10[8].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6668 VDREF single_10b_cdac_0.x6[4].x1.x4.A single_10b_cdac_0.x6[4].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6669 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6670 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6671 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6672 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6673 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6674 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6675 single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6676 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x8.A single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6677 VDREF single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6678 single_10b_cdac_0.x6[5].x2.swn single_10b_cdac_0.x6[5].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6679 single_10b_cdac_0.x8[6].x3.ck single_10b_cdac_0.x8[6].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6680 single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6681 VDREF single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6682 VSREF single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6683 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6684 VCM single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6685 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6686 single_10b_cdac_0.x10b_cap_array_0.SW[4] single_10b_cdac_0.cdac_sw_4_1.x3.ckb a_47370_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6687 VSREF single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6688 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6689 VDREF single_10b_cdac_1.x3[1].x1.x4.A single_10b_cdac_1.x3[1].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6690 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6691 single_10b_cdac_1.cdac_sw_1_1.x3.ck single_10b_cdac_1.cdac_sw_1_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6692 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6693 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6694 single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6695 VSREF SWN_IN[5] a_51468_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6696 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6697 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6698 VDREF CF[9] single_10b_cdac_0.cdac_sw_1_2.x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6699 VDREF single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6700 VSREF single_10b_cdac_0.x3[0].x1.x9.A single_10b_cdac_0.x3[0].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6701 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6702 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6703 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6704 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6705 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6706 single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6707 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6708 single_10b_cdac_1.cdac_sw_1_0.x3.ck single_10b_cdac_1.cdac_sw_1_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6709 single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6710 VDREF single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6711 VDREF single_10b_cdac_0.x4[2].x1.x9.A single_10b_cdac_0.x4[2].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6712 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6713 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6714 single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6715 single_10b_cdac_0.x3[1].x3.ck single_10b_cdac_0.x3[1].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6716 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6717 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6718 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6719 VDREF single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6720 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6721 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6722 VDREF SWP_IN[4] a_52932_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6723 VSREF SWN_IN[2] a_41808_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6724 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6725 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6726 a_29137_36566# single_10b_cdac_1.x3[1].x1.x8.A single_10b_cdac_1.x3[1].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6727 a_52054_34009# SWP_IN[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6728 single_10b_cdac_0.cdac_sw_8_1.x1.x3.Y CF[2] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6729 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6730 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x8.A single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6731 single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6732 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6733 single_10b_cdac_0.x3[0].x2.swn single_10b_cdac_0.x3[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6734 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6735 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6736 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6737 VDREF single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6738 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6739 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6740 single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6741 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6742 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6743 VCM single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[6] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6744 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6745 a_42394_34645# SWP_IN[7] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6746 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6747 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6748 VDREF single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6749 a_22558_31002# single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6750 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6751 VSREF CF[4] single_10b_cdac_0.x6[4].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6752 single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6753 a_21680_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6754 single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.cdac_sw_4_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6755 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6756 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6757 VDREF single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6758 single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6759 VDREF single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6760 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6761 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6762 a_40930_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6763 single_10b_cdac_0.x6[5].x3.ck single_10b_cdac_0.x6[5].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6764 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6765 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6766 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x8.A single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6767 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6768 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6769 single_10b_cdac_1.cdac_sw_2_0.x1.x7.A single_10b_cdac_1.cdac_sw_2_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6770 VDREF single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6771 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6772 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6773 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x8.A single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6774 VSREF single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6775 single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6776 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6777 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6778 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6779 single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6780 VSREF single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6781 VDREF single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6782 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6783 VSREF single_10b_cdac_1.x6[5].x1.x8.A single_10b_cdac_1.x6[5].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6784 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6785 VCM single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6786 single_10b_cdac_0.cdac_sw_2_0.x1.x9.A single_10b_cdac_0.cdac_sw_2_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6787 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6788 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6789 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6790 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6791 single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6792 single_10b_cdac_0.cdac_sw_4_0.x1.x9.A single_10b_cdac_0.cdac_sw_4_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6793 VSREF single_10b_cdac_0.x4[2].x1.x9.A single_10b_cdac_0.x4[2].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6794 VDREF single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6795 single_10b_cdac_1.cdac_sw_1_0.x2.swn single_10b_cdac_1.cdac_sw_1_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6796 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6797 VDREF single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6798 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6799 single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6800 single_10b_cdac_1.x10b_cap_array_0.SW[8] single_10b_cdac_1.cdac_sw_1_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6801 single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6802 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6803 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6804 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6805 VSREF single_10b_cdac_0.cdac_sw_4_1.x1.x9.A single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6806 VDREF SWP_IN[3] a_56152_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6807 VSREF single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6808 VDREF single_10b_cdac_1.x3[1].x1.x3.Y single_10b_cdac_1.x3[1].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6809 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6810 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x3.ck a_55274_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6811 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6812 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6813 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6814 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6815 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6816 single_10b_cdac_1.x6[4].x2.swn single_10b_cdac_1.x6[4].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6817 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6818 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6819 VSREF single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6820 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6821 single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6822 VSREF single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6823 VSREF single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6824 a_48248_25713# single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6825 single_10b_cdac_0.cdac_sw_2_0.x1.x5.A single_10b_cdac_0.cdac_sw_2_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6826 single_10b_cdac_1.x8[6].x3.ck single_10b_cdac_1.x8[6].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6827 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6828 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6829 single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.cdac_sw_2_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6830 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6831 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6832 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6833 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6834 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6835 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6836 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6837 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6838 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6839 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6840 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6841 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6842 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6843 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6844 VSREF single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6845 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6846 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x8.A single_10b_cdac_1.cdac_sw_2_1.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6847 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6848 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6849 a_45028_25713# single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6850 VDREF single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6851 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x9.A single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6852 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6853 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6854 VDREF single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6855 single_10b_cdac_1.x4[2].x3.ck single_10b_cdac_1.x4[2].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6856 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6857 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6858 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6859 VSREF single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6860 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6861 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6862 a_7336_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6863 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6864 single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6865 single_10b_cdac_1.x4[2].x2.swn single_10b_cdac_1.x4[2].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6866 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6867 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x8.A single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6868 single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6869 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6870 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6871 single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6872 VSREF single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6873 single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6874 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6875 VDREF single_10b_cdac_1.x6[4].x1.x7.A single_10b_cdac_1.x6[4].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6876 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6877 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6878 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6879 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6880 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6881 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6882 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6883 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6884 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6885 single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6886 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6887 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6888 VSREF single_10b_cdac_1.x10[8].x1.x3.Y a_6597_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6889 VDREF single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6890 VDREF CF[7] single_10b_cdac_1.cdac_sw_2_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6891 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6892 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6893 single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6894 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6895 single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6896 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6897 single_10b_cdac_0.cdac_sw_4_1.x1.x7.A single_10b_cdac_0.cdac_sw_4_1.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6898 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x9.A single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6899 single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6900 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6901 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6902 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6903 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6904 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6905 VDREF single_10b_cdac_1.x8[6].x1.x4.A single_10b_cdac_1.x8[6].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6906 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6907 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6908 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6909 single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.cdac_sw_8_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6910 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6911 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6912 single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6913 single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6914 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6915 VDREF single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6916 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x8.A single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6917 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6918 VDREF single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6919 single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6920 VSREF single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6921 single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6922 VDREF single_10b_cdac_0.x8[7].x1.x9.A single_10b_cdac_0.x8[7].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6923 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6924 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6925 single_10b_cdac_1.cdac_sw_1_2.x3.ck single_10b_cdac_1.cdac_sw_1_2.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6926 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6927 VSREF single_10b_cdac_1.x10[8].x1.x7.A single_10b_cdac_1.x10[8].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6928 single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6929 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6930 single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6931 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6932 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6933 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6934 a_13037_36566# single_10b_cdac_1.x8[6].x1.x8.A single_10b_cdac_1.x8[6].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6935 VSREF single_10b_cdac_1.x4[2].x1.x4.A single_10b_cdac_1.x4[2].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6936 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6937 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x8.A single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6938 single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6939 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6940 VSREF single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6941 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x3.ck a_58494_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6942 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6943 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6944 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6945 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6946 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6947 VSREF single_10b_cdac_0.x4[3].x1.x9.A a_56291_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6948 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6949 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6950 VDREF single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6951 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6952 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6953 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6954 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6955 single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6956 single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6957 VSREF single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6958 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6959 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x9.A single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6960 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6961 single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6962 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6963 single_10b_cdac_0.cdac_sw_8_0.x1.x5.A single_10b_cdac_0.cdac_sw_8_0.x1.x8.A a_44243_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6964 VDREF single_10b_cdac_1.x3[1].x1.x9.A single_10b_cdac_1.x3[1].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6965 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6966 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6967 single_10b_cdac_0.cdac_sw_1_0.x3.ck single_10b_cdac_0.cdac_sw_1_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6968 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6969 VCP single_10b_cdac_0.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6970 single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.cdac_sw_2_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6971 VCP single_10b_cdac_0.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6972 VDREF single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6973 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6974 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6975 VSREF single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6976 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6977 VSREF single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6978 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6979 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x4.A single_10b_cdac_1.cdac_sw_1_2.x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6980 a_44150_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6981 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6982 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6983 single_10b_cdac_0.x8[6].x3.ck single_10b_cdac_0.x8[6].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6984 single_10b_cdac_1.x10b_cap_array_0.SW[7] single_10b_cdac_1.cdac_sw_2_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6985 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6986 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6987 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6988 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6989 single_10b_cdac_0.cdac_sw_8_1.x1.x9.A single_10b_cdac_0.cdac_sw_8_1.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6990 VDREF SWP_IN[3] a_22558_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6991 single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6992 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6993 single_10b_cdac_1.x6[5].dac_out single_10b_cdac_1.x6[5].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6994 VSREF single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6995 VSREF single_10b_cdac_0.x8[7].x1.x9.A single_10b_cdac_0.x8[7].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6996 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6997 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6998 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6999 VDREF single_10b_cdac_0.x2[0].x1.x9.A single_10b_cdac_0.x2[0].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7000 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7001 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7002 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7003 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7004 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7005 VDREF single_10b_cdac_1.x8[6].x1.x3.Y single_10b_cdac_1.x8[6].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7006 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7007 single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7008 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7009 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7010 single_10b_cdac_1.cdac_sw_8_0.x1.x6.A single_10b_cdac_1.cdac_sw_8_0.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7011 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7012 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7013 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7014 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7015 single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7016 VSREF single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7017 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7018 single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7019 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7020 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7021 single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.cdac_sw_2_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7022 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7023 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7024 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7025 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7026 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7027 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7028 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7029 single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.cdac_sw_8_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7030 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7031 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7032 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7033 VSREF single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7034 a_11434_25713# single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7035 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7036 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7037 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7038 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7039 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7040 single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7041 VSREF single_10b_cdac_1.x10[8].x1.x9.A single_10b_cdac_1.x10[8].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7042 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7043 single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7044 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7045 VSREF single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7046 single_10b_cdac_0.cdac_sw_1_0.x1.x5.A single_10b_cdac_0.cdac_sw_1_0.x1.x8.A a_63563_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7047 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7048 single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7049 single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7050 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7051 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7052 single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.cdac_sw_2_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7053 VCM single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7054 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7055 single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.cdac_sw_4_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7056 VCM single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7057 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7058 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x11.A single_10b_cdac_1.cdac_sw_1_2.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7059 single_10b_cdac_1.x3[1].x3.ck single_10b_cdac_1.x3[1].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7060 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7061 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7062 VCP single_10b_cdac_1.x3[0].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7063 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7064 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7065 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7066 single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7067 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7068 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7069 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7070 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7071 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7072 VSREF single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7073 VDREF single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7074 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7075 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7076 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x8.A single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7077 single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7078 single_10b_cdac_0.cdac_sw_1_1.x1.x9.A single_10b_cdac_0.cdac_sw_1_1.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7079 single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7080 single_10b_cdac_0.x10[8].x3.ck single_10b_cdac_0.x10[8].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7081 VCM single_10b_cdac_1.cdac_sw_1_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[8] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7082 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7083 VSREF single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7084 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7085 VSREF single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7086 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7087 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7088 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7089 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7090 VDREF single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7091 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x9.A single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7092 single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7093 single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7094 VDREF single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7095 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7096 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7097 VSREF SWN_IN[3] a_45028_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7098 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7099 VDREF single_10b_cdac_1.x3[0].x1.x3.Y single_10b_cdac_1.x3[0].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7100 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7101 single_10b_cdac_0.x6[5].dac_out single_10b_cdac_0.x6[5].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7102 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7103 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7104 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7105 single_10b_cdac_1.cdac_sw_1_0.x1.x9.A single_10b_cdac_1.cdac_sw_1_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7106 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7107 VDREF single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7108 VDREF single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7109 single_10b_cdac_0.cdac_sw_1_0.x3.ck single_10b_cdac_0.cdac_sw_1_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7110 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7111 single_10b_cdac_0.cdac_sw_1_1.x1.x5.A single_10b_cdac_0.cdac_sw_1_1.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7112 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x8.A single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7113 VCN single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7114 VSREF SWN_IN[5] a_17874_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7115 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7116 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7117 single_10b_cdac_0.x10[8].dac_out single_10b_cdac_0.x10[8].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7118 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7119 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7120 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7121 single_10b_cdac_0.cdac_sw_16_0.x1.x3.Y CF[0] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7122 single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7123 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7124 VCM single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7125 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7126 a_24900_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7127 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7128 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7129 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7130 VSREF single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7131 single_10b_cdac_0.x4[2].x2.swn single_10b_cdac_0.x4[2].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7132 single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7133 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7134 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7135 single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7136 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7137 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7138 single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7139 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7140 single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7141 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7142 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7143 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7144 a_16118_33146# single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7145 VDREF CF[4] single_10b_cdac_1.x6[4].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7146 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7147 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7148 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7149 a_15240_34009# SWP_IN[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7150 VCM single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[6] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7151 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7152 VSREF single_10b_cdac_0.x10[8].x1.x9.A a_40191_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7153 VSREF SWN_IN[3] a_11434_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7154 single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7155 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7156 VCM single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7157 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7158 VSREF single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7159 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7160 single_10b_cdac_0.cdac_sw_1_0.x1.x4.A single_10b_cdac_0.cdac_sw_1_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7161 VCN single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7162 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7163 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7164 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7165 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7166 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7167 single_10b_cdac_1.cdac_sw_4_0.x1.x6.A single_10b_cdac_1.cdac_sw_4_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7168 VDREF single_10b_cdac_1.x8[6].x1.x9.A single_10b_cdac_1.x8[6].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7169 VSREF single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7170 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7171 single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7172 single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.cdac_sw_4_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7173 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7174 single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7175 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7176 single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x2[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7177 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7178 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7179 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7180 single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7181 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7182 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7183 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7184 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7185 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7186 VDREF single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7187 VCN single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7188 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7189 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7190 single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7191 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7192 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7193 single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.cdac_sw_2_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7194 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7195 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7196 VDREF single_10b_cdac_0.x8[6].x1.x8.A single_10b_cdac_0.x8[6].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7197 VSREF single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7198 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7199 single_10b_cdac_1.x3[0].x3.ck single_10b_cdac_1.x3[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7200 single_10b_cdac_0.x6[5].dac_out single_10b_cdac_0.x6[5].x3.ck a_48834_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7201 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7202 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7203 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7204 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7205 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7206 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7207 single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7208 single_10b_cdac_0.cdac_sw_4_0.x3.ck single_10b_cdac_0.cdac_sw_4_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7209 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7210 single_10b_cdac_0.x3[0].x2.swn single_10b_cdac_0.x3[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7211 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7212 single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7213 VDREF single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7214 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7215 VSREF single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7216 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7217 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7218 VSREF single_10b_cdac_0.x4[2].x1.x8.A single_10b_cdac_0.x4[2].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7219 single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7220 a_61128_25713# single_10b_cdac_0.cdac_sw_1_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[8] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7221 single_10b_cdac_1.cdac_sw_1_1.x3.ck single_10b_cdac_1.cdac_sw_1_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7222 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7223 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7224 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7225 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7226 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7227 VSREF single_10b_cdac_1.x8[7].x1.x8.A single_10b_cdac_1.x8[7].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7228 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7229 VSREF single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7230 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7231 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7232 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7233 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7234 single_10b_cdac_1.x10b_cap_array_0.SW[5] single_10b_cdac_1.cdac_sw_4_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7235 VCM single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7236 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x3.ck a_58494_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7237 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7238 single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7239 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7240 VDREF single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7241 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7242 VSREF single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7243 single_10b_cdac_1.x6[4].x3.ck single_10b_cdac_1.x6[4].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7244 single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7245 VSREF single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7246 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x8.A single_10b_cdac_0.cdac_sw_2_1.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7247 VSREF single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7248 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7249 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7250 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7251 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7252 single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7253 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7254 single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.cdac_sw_8_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7255 VCM single_10b_cdac_0.cdac_sw_1_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[8] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7256 VSREF SWN_IN[4] a_14654_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7257 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7258 single_10b_cdac_1.x8[6].x3.ck single_10b_cdac_1.x8[6].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7259 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7260 a_56152_31002# single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7261 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7262 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7263 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7264 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7265 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7266 single_10b_cdac_0.x6[4].x1.x5.A single_10b_cdac_0.x6[4].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7267 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7268 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7269 VDREF CF[5] single_10b_cdac_1.cdac_sw_4_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7270 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7271 VDREF single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7272 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7273 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7274 single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7275 single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7276 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x9.A single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7277 VCM single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7278 VSREF single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7279 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7280 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7281 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7282 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7283 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7284 single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7285 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7286 VSREF single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7287 single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7288 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x3.ck a_24900_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7289 single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7290 a_23436_25722# SWN_IN[7] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7291 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7292 single_10b_cdac_1.x4[2].x3.ck single_10b_cdac_1.x4[2].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7293 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7294 single_10b_cdac_1.cdac_sw_2_1.x1.x9.A single_10b_cdac_1.cdac_sw_2_1.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7295 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7296 single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7297 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7298 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7299 single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7300 VSREF single_10b_cdac_1.x4[3].x1.x9.A single_10b_cdac_1.x4[3].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7301 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x9.A single_10b_cdac_0.cdac_sw_1_2.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7302 single_10b_cdac_1.cdac_sw_1_2.x3.ck single_10b_cdac_1.cdac_sw_1_2.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7303 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7304 single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x2[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7305 VDREF single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7306 single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.cdac_sw_16_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7307 VSREF single_10b_cdac_1.x3[1].x1.x7.A single_10b_cdac_1.x3[1].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7308 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7309 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7310 VDREF single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7311 single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7312 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7313 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7314 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7315 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7316 VSREF single_10b_cdac_1.x6[4].x1.x4.A single_10b_cdac_1.x6[4].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7317 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7318 single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7319 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7320 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7321 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7322 single_10b_cdac_0.x8[7].x2.swn single_10b_cdac_0.x8[7].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7323 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7324 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7325 a_56152_31002# single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7326 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7327 single_10b_cdac_0.cdac_sw_1_1.x2.swn single_10b_cdac_0.cdac_sw_1_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7328 single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7329 single_10b_cdac_1.cdac_sw_2_1.x1.x5.A single_10b_cdac_1.cdac_sw_2_1.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7330 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7331 VDREF single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7332 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7333 single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7334 VSREF single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7335 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7336 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7337 single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7338 VSREF single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7339 VDREF single_10b_cdac_1.x4[2].x1.x9.A single_10b_cdac_1.x4[2].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7340 VDREF single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7341 single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x2[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7342 single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7343 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7344 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7345 VDREF single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7346 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7347 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7348 single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.cdac_sw_16_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7349 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7350 VSREF SWN_IN[2] a_8214_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7351 single_10b_cdac_0.x10b_cap_array_0.SW[7] single_10b_cdac_0.cdac_sw_2_0.x3.ckb a_57030_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7352 VDREF single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7353 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7354 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7355 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7356 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7357 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7358 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7359 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7360 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7361 single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7362 a_6597_36566# single_10b_cdac_1.x10[8].x1.x8.A single_10b_cdac_1.x10[8].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7363 single_10b_cdac_1.cdac_sw_2_0.x1.x4.A single_10b_cdac_1.cdac_sw_2_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7364 VCM single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7365 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7366 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7367 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7368 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7369 single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7370 VDREF single_10b_cdac_1.x4[2].x1.x6.A single_10b_cdac_1.x4[2].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7371 single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7372 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7373 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7374 VSREF single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7375 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7376 VCP single_10b_cdac_1.x3[1].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7377 single_10b_cdac_0.cdac_sw_2_1.x1.x6.A single_10b_cdac_0.cdac_sw_2_1.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7378 single_10b_cdac_0.cdac_sw_16_0.x1.x9.A single_10b_cdac_0.cdac_sw_16_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7379 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7380 VSREF single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7381 VDREF single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7382 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7383 single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7384 VSREF single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7385 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7386 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x9.A single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7387 single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7388 single_10b_cdac_0.x10b_cap_array_0.SW[7] single_10b_cdac_0.cdac_sw_2_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7389 single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.cdac_sw_8_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7390 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7391 single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7392 single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7393 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7394 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7395 VDREF single_10b_cdac_1.x6[5].x1.x5.A single_10b_cdac_1.x6[5].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7396 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7397 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7398 VDREF single_10b_cdac_1.x2[0].x1.x9.A single_10b_cdac_1.x2[0].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7399 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7400 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7401 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7402 VDREF single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7403 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7404 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7405 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7406 single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7407 single_10b_cdac_1.x6[4].dac_out single_10b_cdac_1.x6[4].x3.ck a_18460_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7408 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7409 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7410 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7411 single_10b_cdac_0.x8[7].dac_out single_10b_cdac_0.x8[7].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7412 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7413 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7414 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7415 VDREF single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7416 VDREF single_10b_cdac_0.x8[6].x1.x3.Y single_10b_cdac_0.x8[6].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7417 single_10b_cdac_1.x10[8].x2.swn single_10b_cdac_1.x10[8].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7418 single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.cdac_sw_4_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7419 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7420 VSREF single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7421 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7422 a_59372_31002# single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7423 a_63470_25722# SWN_IN[9] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7424 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7425 single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7426 single_10b_cdac_0.cdac_sw_1_2.x2.swn single_10b_cdac_0.cdac_sw_1_2.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7427 VDREF single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7428 single_10b_cdac_1.x6[4].dac_out single_10b_cdac_1.x6[4].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7429 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7430 single_10b_cdac_0.x2[0].x1.x8.A single_10b_cdac_0.x2[0].x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7431 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7432 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7433 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7434 VSREF single_10b_cdac_0.x8[7].x1.x8.A single_10b_cdac_0.x8[7].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7435 a_55274_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7436 single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.cdac_sw_8_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7437 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7438 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7439 a_45028_25713# single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7440 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7441 single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7442 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7443 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7444 single_10b_cdac_0.x8[7].dac_out single_10b_cdac_0.x8[7].x3.ck a_42394_34645# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7445 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x9.A single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7446 single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7447 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7448 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7449 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x3.ck a_21680_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7450 VDREF SWP_IN[3] a_22558_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7451 VDREF single_10b_cdac_0.x8[6].x1.x7.A single_10b_cdac_0.x8[6].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7452 VSREF single_10b_cdac_1.x6[4].x1.x8.A single_10b_cdac_1.x6[4].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7453 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7454 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7455 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7456 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7457 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7458 VSREF single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7459 a_17874_25713# single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7460 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7461 a_49851_36566# single_10b_cdac_0.x6[5].x1.x8.A single_10b_cdac_0.x6[5].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7462 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7463 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7464 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7465 VSREF single_10b_cdac_0.x3[1].x1.x3.Y a_62731_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7466 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7467 VSREF single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7468 VCM single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7469 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7470 single_10b_cdac_0.cdac_sw_1_2.x2.swn single_10b_cdac_0.cdac_sw_1_2.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7471 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7472 single_10b_cdac_1.cdac_sw_1_1.x2.swn single_10b_cdac_1.cdac_sw_1_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7473 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7474 a_14654_25713# single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7475 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7476 single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.cdac_sw_2_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7477 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7478 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7479 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7480 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7481 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7482 single_10b_cdac_0.cdac_sw_2_1.x1.x8.A single_10b_cdac_0.cdac_sw_2_1.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7483 VDREF SWP_IN[5] a_49712_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7484 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7485 VSREF single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7486 VSREF single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7487 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7488 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7489 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7490 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7491 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7492 VSREF single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7493 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7494 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7495 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7496 single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7497 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x9.A single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7498 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7499 single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7500 VDREF single_10b_cdac_1.x10[8].x1.x5.A single_10b_cdac_1.x10[8].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7501 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7502 VSREF single_10b_cdac_0.x3[1].x1.x7.A single_10b_cdac_0.x3[1].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7503 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7504 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7505 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7506 single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7507 a_6458_34754# single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7508 VCN single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7509 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7510 VDREF single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7511 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7512 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7513 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7514 single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.cdac_sw_2_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7515 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7516 single_10b_cdac_0.x6[4].x2.swn single_10b_cdac_0.x6[4].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7517 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7518 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7519 single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7520 VSREF single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7521 VSREF single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7522 VDREF single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7523 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7524 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7525 VSREF single_10b_cdac_1.x8[6].x1.x7.A single_10b_cdac_1.x8[6].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7526 single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7527 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7528 VSREF single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7529 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7530 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7531 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7532 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7533 single_10b_cdac_0.x8[6].x3.ck single_10b_cdac_0.x8[6].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7534 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7535 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7536 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7537 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7538 VSREF SWN_IN[4] a_48248_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7539 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7540 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7541 VSREF single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7542 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7543 VSREF single_10b_cdac_0.x8[6].x1.x5.A single_10b_cdac_0.x8[6].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7544 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7545 VDREF single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7546 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7547 VDREF single_10b_cdac_0.x3[0].x1.x7.A single_10b_cdac_0.x3[0].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7548 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7549 single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7550 single_10b_cdac_0.cdac_sw_1_1.x1.x3.Y CF[8] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7551 VSREF single_10b_cdac_1.x8[7].x1.x8.A single_10b_cdac_1.x8[7].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7552 VCM single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7553 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7554 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7555 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7556 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7557 VSREF single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7558 a_8214_25713# single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7559 a_48834_34009# SWP_IN[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7560 single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7561 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7562 single_10b_cdac_1.x8[7].dac_out single_10b_cdac_1.x8[7].x3.ck a_8800_34645# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7563 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7564 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7565 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7566 VDREF single_10b_cdac_0.x6[4].x1.x8.A single_10b_cdac_0.x6[4].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7567 single_10b_cdac_1.cdac_sw_4_0.x1.x3.Y CF[5] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7568 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7569 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7570 single_10b_cdac_1.x10[8].x2.swn single_10b_cdac_1.x10[8].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7571 a_59511_35702# CF[2] single_10b_cdac_0.x4[2].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7572 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7573 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7574 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7575 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7576 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7577 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x3.ckb a_40930_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7578 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7579 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7580 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7581 single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7582 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x3.ckb a_7336_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7583 single_10b_cdac_1.x3[0].x2.swn single_10b_cdac_1.x3[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7584 single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7585 VDREF single_10b_cdac_1.x3[1].x1.x8.A single_10b_cdac_1.x3[1].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7586 VDREF single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7587 a_18460_34009# SWP_IN[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7588 single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7589 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7590 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7591 VSREF CF[1] single_10b_cdac_1.x3[1].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7592 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7593 VSREF single_10b_cdac_1.x4[3].x1.x9.A a_22697_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7594 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7595 single_10b_cdac_0.x6[4].x3.ck single_10b_cdac_0.x6[4].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7596 VSREF single_10b_cdac_0.x3[0].x1.x8.A single_10b_cdac_0.x3[0].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7597 VCM single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7598 a_49712_33146# single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7599 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7600 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7601 single_10b_cdac_1.x3[0].x1.x5.A single_10b_cdac_1.x3[0].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7602 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7603 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7604 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7605 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7606 single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7607 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7608 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7609 VDREF single_10b_cdac_0.x10[8].x1.x8.A single_10b_cdac_0.x10[8].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7610 single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7611 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7612 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7613 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7614 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7615 single_10b_cdac_0.x8[6].x2.swn single_10b_cdac_0.x8[6].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7616 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7617 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7618 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7619 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7620 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7621 VSREF single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7622 single_10b_cdac_0.x3[0].x3.ck single_10b_cdac_0.x3[0].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7623 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7624 single_10b_cdac_0.x10b_cap_array_0.SW[5] single_10b_cdac_0.cdac_sw_4_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7625 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7626 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7627 single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.cdac_sw_2_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7628 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7629 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7630 VSREF single_10b_cdac_1.x4[3].x1.x6.A single_10b_cdac_1.x4[3].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7631 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7632 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7633 single_10b_cdac_0.x3[0].x1.x4.A CF[0] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7634 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7635 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7636 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7637 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7638 single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7639 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7640 VDREF single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7641 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7642 VSREF single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7643 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7644 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7645 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7646 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7647 VSREF SWN_IN[7] a_57908_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7648 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x8.A single_10b_cdac_0.cdac_sw_4_1.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7649 VSREF single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7650 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7651 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7652 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7653 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7654 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7655 VDREF single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7656 single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7657 single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7658 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7659 single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.cdac_sw_16_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7660 VDREF single_10b_cdac_0.x3[1].x1.x9.A single_10b_cdac_0.x3[1].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7661 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7662 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7663 single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7664 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7665 single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.cdac_sw_8_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7666 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7667 VDREF single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7668 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7669 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7670 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7671 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7672 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7673 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7674 VDREF SWP_IN[2] a_25778_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7675 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7676 single_10b_cdac_1.x4[3].x2.swn single_10b_cdac_1.x4[3].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7677 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7678 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7679 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7680 VDREF single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7681 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7682 single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7683 VSREF single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7684 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x8.A single_10b_cdac_1.cdac_sw_8_1.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7685 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x8.A single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7686 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7687 single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7688 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7689 single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7690 VDREF single_10b_cdac_0.x3[1].x1.x4.A single_10b_cdac_0.x3[1].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7691 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7692 VSREF single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7693 single_10b_cdac_1.cdac_sw_16_0.x1.x5.A single_10b_cdac_1.cdac_sw_16_0.x1.x8.A a_989_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7694 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7695 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7696 single_10b_cdac_1.cdac_sw_4_1.x1.x9.A single_10b_cdac_1.cdac_sw_4_1.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7697 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7698 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7699 single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7700 single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.cdac_sw_2_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7701 VSREF single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7702 VDREF single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7703 VSREF single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7704 VSREF single_10b_cdac_1.x6[5].x1.x9.A single_10b_cdac_1.x6[5].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7705 single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.cdac_sw_4_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7706 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7707 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7708 single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.cdac_sw_8_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7709 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7710 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7711 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7712 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7713 single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7714 single_10b_cdac_1.x8[6].dac_out single_10b_cdac_1.x8[6].x3.ck a_12020_34645# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7715 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7716 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7717 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7718 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7719 single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7720 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7721 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7722 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7723 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7724 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x8.A single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7725 single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.cdac_sw_2_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7726 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7727 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7728 VSREF single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7729 single_10b_cdac_1.cdac_sw_4_0.x1.x8.A single_10b_cdac_1.cdac_sw_4_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7730 single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7731 VSREF single_10b_cdac_1.x6[4].x3.ckb single_10b_cdac_1.x6[4].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7732 VSREF SWN_IN[3] a_11434_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7733 single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7734 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7735 VSREF single_10b_cdac_1.x4[3].x1.x8.A single_10b_cdac_1.x4[3].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7736 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7737 VDREF single_10b_cdac_1.x6[4].x1.x9.A single_10b_cdac_1.x6[4].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7738 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7739 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7740 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7741 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7742 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7743 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7744 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7745 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x3.ck a_21680_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7746 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7747 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7748 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7749 single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.cdac_sw_16_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7750 VDREF single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7751 a_43411_35702# CF[7] single_10b_cdac_0.x8[7].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7752 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7753 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7754 single_10b_cdac_1.cdac_sw_1_1.x2.swn single_10b_cdac_1.cdac_sw_1_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7755 single_10b_cdac_1.x4[2].x2.swn single_10b_cdac_1.x4[2].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7756 single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7757 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7758 single_10b_cdac_1.cdac_sw_4_0.x1.x4.A single_10b_cdac_1.cdac_sw_4_0.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7759 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7760 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7761 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7762 single_10b_cdac_1.x6[5].x2.swn single_10b_cdac_1.x6[5].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7763 single_10b_cdac_0.cdac_sw_16_0.x1.x6.A single_10b_cdac_0.cdac_sw_16_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7764 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x8.A single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7765 VDREF single_10b_cdac_1.x8[6].x1.x8.A single_10b_cdac_1.x8[6].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7766 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7767 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7768 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7769 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7770 VDREF single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7771 single_10b_cdac_0.cdac_sw_1_1.x2.swn single_10b_cdac_0.cdac_sw_1_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7772 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7773 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7774 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7775 single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.cdac_sw_16_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7776 VSREF CF[6] single_10b_cdac_1.x8[6].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7777 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7778 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7779 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7780 single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7781 single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7782 VDREF single_10b_cdac_0.x4[2].x1.x6.A single_10b_cdac_0.x4[2].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7783 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7784 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7785 VSREF single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7786 VSREF single_10b_cdac_1.x8[7].x1.x10.A single_10b_cdac_1.x8[7].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7787 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7788 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7789 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x9.A single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7790 single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x2[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7791 VDREF single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7792 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7793 VDREF single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7794 VDREF CF[0] single_10b_cdac_0.x3[0].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7795 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7796 VDREF single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7797 single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7798 VDREF single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7799 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7800 VDREF single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7801 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7802 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x9.A single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7803 single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7804 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7805 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7806 single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.cdac_sw_4_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7807 VSREF single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7808 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7809 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7810 single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7811 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7812 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7813 single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7814 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7815 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7816 single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7817 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7818 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7819 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7820 single_10b_cdac_1.x4[2].x1.x4.A CF[2] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7821 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7822 VDREF single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7823 single_10b_cdac_0.cdac_sw_1_2.dac_out single_10b_cdac_0.cdac_sw_1_2.x3.ck a_35954_34963# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7824 VSREF single_10b_cdac_1.x4[2].x1.x5.A single_10b_cdac_1.x4[2].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7825 VDREF SWP_IN[5] a_16118_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7826 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7827 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7828 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7829 VSREF SWN_IN[2] a_41808_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7830 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7831 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7832 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7833 single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7834 a_62731_35702# CF[1] single_10b_cdac_0.x3[1].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7835 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7836 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7837 VSREF single_10b_cdac_0.x4[3].x1.x3.Y a_56291_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7838 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7839 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7840 VSREF single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7841 VCM single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7842 single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7843 VDREF single_10b_cdac_1.x3[0].x1.x8.A single_10b_cdac_1.x3[0].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7844 VDREF single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7845 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7846 VCM single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7847 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7848 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7849 single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.cdac_sw_8_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7850 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7851 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7852 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7853 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7854 single_10b_cdac_0.cdac_sw_4_1.x1.x8.A single_10b_cdac_0.cdac_sw_4_1.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7855 single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7856 VDREF single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7857 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7858 a_50683_24080# single_10b_cdac_0.cdac_sw_4_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7859 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7860 VCN single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7861 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7862 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7863 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7864 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7865 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7866 single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7867 single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7868 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7869 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7870 VDREF single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7871 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7872 single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.cdac_sw_8_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7873 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7874 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7875 VDREF single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7876 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7877 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7878 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7879 VDREF single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7880 VDREF CF[0] single_10b_cdac_0.cdac_sw_16_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7881 single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7882 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7883 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7884 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7885 VCP single_10b_cdac_0.x4[2].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7886 VDREF single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7887 single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7888 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7889 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7890 single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7891 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7892 single_10b_cdac_0.x8[6].x2.swn single_10b_cdac_0.x8[6].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7893 VDREF single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7894 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7895 VSREF single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7896 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7897 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7898 VDREF SWP_IN[4] a_52932_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7899 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7900 VCN single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7901 VDREF single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7902 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7903 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7904 VSREF single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7905 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7906 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7907 single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7908 single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7909 VSREF single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7910 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7911 VDREF single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7912 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7913 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7914 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7915 single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7916 single_10b_cdac_0.cdac_sw_1_1.x3.ck single_10b_cdac_0.cdac_sw_1_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7917 single_10b_cdac_1.x10b_cap_array_0.SW[4] single_10b_cdac_1.cdac_sw_4_1.x3.ckb a_13776_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7918 VSREF single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7919 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7920 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7921 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7922 single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.cdac_sw_8_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7923 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7924 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7925 a_22558_31002# single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7926 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7927 single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x2[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7928 single_10b_cdac_0.cdac_sw_4_0.x1.x4.A CF[5] a_50683_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7929 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7930 VSREF SWN_IN[8] a_61128_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7931 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7932 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7933 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7934 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7935 single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7936 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7937 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7938 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7939 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x8.A single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7940 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7941 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7942 VSREF single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7943 single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7944 VDREF single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7945 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7946 single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.cdac_sw_4_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7947 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7948 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7949 VDREF single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7950 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7951 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7952 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7953 single_10b_cdac_1.x3[1].x3.ck single_10b_cdac_1.x3[1].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7954 a_34490_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7955 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7956 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7957 single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7958 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7959 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7960 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7961 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7962 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7963 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7964 VSREF single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7965 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7966 single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7967 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7968 single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7969 VDREF single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7970 VSREF single_10b_cdac_1.x6[5].x1.x9.A a_16257_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7971 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7972 single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.cdac_sw_4_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7973 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7974 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7975 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7976 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7977 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7978 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7979 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7980 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7981 a_8214_25713# single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7982 VCM single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7983 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7984 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7985 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7986 VSREF single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7987 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7988 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7989 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7990 single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7991 VDREF single_10b_cdac_0.x8[7].x1.x6.A single_10b_cdac_0.x8[7].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7992 single_10b_cdac_0.x3[1].x2.swn single_10b_cdac_0.x3[1].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7993 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7994 VSREF single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7995 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7996 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7997 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7998 VSREF single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7999 VDREF SWP_IN[3] a_56152_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8000 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8001 single_10b_cdac_0.x10b_cap_array_0.SW[8] single_10b_cdac_0.cdac_sw_1_1.x3.ckb a_60250_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8002 single_10b_cdac_0.x10[8].x2.swn single_10b_cdac_0.x10[8].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8003 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8004 VSREF single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8005 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x9.A single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8006 single_10b_cdac_1.x10b_cap_array_0.SW[7] single_10b_cdac_1.cdac_sw_2_0.x3.ckb a_23436_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8007 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8008 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8009 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8010 VSREF single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8011 VDREF CF[5] single_10b_cdac_0.x6[5].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8012 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8013 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8014 single_10b_cdac_1.x2[0].x1.x3.Y CF[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8015 single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.cdac_sw_4_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8016 VSREF single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8017 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8018 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8019 VDREF single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8020 single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8021 single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8022 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8023 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8024 VCM single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8025 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8026 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8027 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8028 VSREF single_10b_cdac_0.x4[3].x1.x6.A single_10b_cdac_0.x4[3].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8029 a_25778_31002# single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8030 single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8031 single_10b_cdac_1.x10[8].x3.ck single_10b_cdac_1.x10[8].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8032 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8033 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8034 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x9.A single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8035 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8036 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8037 single_10b_cdac_1.cdac_sw_2_1.x1.x6.A single_10b_cdac_1.cdac_sw_2_1.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8038 single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8039 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8040 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8041 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8042 single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8043 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8044 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x8.A single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8045 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8046 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8047 single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8048 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8049 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8050 VSREF single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8051 single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8052 single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8053 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8054 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8055 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8056 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8057 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8058 single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8059 single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8060 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8061 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8062 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8063 single_10b_cdac_1.cdac_sw_1_0.x3.ck single_10b_cdac_1.cdac_sw_1_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8064 VDREF single_10b_cdac_0.x4[3].x1.x9.A single_10b_cdac_0.x4[3].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8065 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8066 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8067 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8068 VSREF single_10b_cdac_0.x10[8].x1.x3.Y a_40191_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8069 VSREF single_10b_cdac_0.x10[8].x1.x4.A single_10b_cdac_0.x10[8].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8070 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8071 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8072 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8073 single_10b_cdac_0.x3[1].x3.ck single_10b_cdac_0.x3[1].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8074 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8075 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8076 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8077 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8078 single_10b_cdac_0.cdac_sw_1_2.x3.ck single_10b_cdac_0.cdac_sw_1_2.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8079 a_22697_35702# CF[3] single_10b_cdac_1.x4[3].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8080 single_10b_cdac_0.cdac_sw_8_1.x1.x5.A single_10b_cdac_0.cdac_sw_8_1.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8081 a_21680_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8082 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8083 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8084 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8085 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8086 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8087 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8088 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8089 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8090 VDREF SWP_IN[2] a_59372_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8091 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8092 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x8.A single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8093 single_10b_cdac_0.x4[3].x2.swn single_10b_cdac_0.x4[3].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8094 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8095 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8096 VSREF single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8097 single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8098 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8099 single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8100 VDREF single_10b_cdac_0.x4[3].x1.x4.A single_10b_cdac_0.x4[3].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8101 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8102 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8103 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8104 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8105 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8106 single_10b_cdac_0.x6[5].x3.ck single_10b_cdac_0.x6[5].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8107 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8108 single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.cdac_sw_4_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8109 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8110 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8111 VDREF single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8112 single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8113 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8114 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8115 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8116 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8117 VDREF single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8118 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8119 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8120 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8121 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8122 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8123 VDREF single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8124 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8125 single_10b_cdac_1.x3[0].x2.swn single_10b_cdac_1.x3[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8126 VSREF single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8127 single_10b_cdac_1.x4[3].x2.swn single_10b_cdac_1.x4[3].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8128 single_10b_cdac_0.cdac_sw_1_2.x3.ckb single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8129 VSREF single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8130 single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8131 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8132 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8133 a_55274_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8134 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8135 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8136 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8137 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x3.ck a_55274_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8138 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8139 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8140 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8141 VSREF single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8142 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8143 single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8144 VSREF single_10b_cdac_0.x4[2].x1.x9.A single_10b_cdac_0.x4[2].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8145 single_10b_cdac_1.cdac_sw_8_1.x1.x9.A single_10b_cdac_1.cdac_sw_8_1.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8146 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x3.Y single_10b_cdac_1.cdac_sw_1_2.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8147 single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8148 single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.cdac_sw_2_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8149 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8150 single_10b_cdac_1.x6[5].dac_out single_10b_cdac_1.x6[5].x3.ck a_15240_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8151 single_10b_cdac_1.cdac_sw_16_0.x1.x9.A single_10b_cdac_1.cdac_sw_16_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8152 VDREF single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8153 single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8154 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8155 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8156 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8157 single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8158 VSREF single_10b_cdac_1.x8[7].x1.x9.A single_10b_cdac_1.x8[7].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8159 single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8160 VDREF single_10b_cdac_1.x6[5].x1.x10.A single_10b_cdac_1.x6[5].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8161 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8162 single_10b_cdac_0.x4[3].x3.ck single_10b_cdac_0.x4[3].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8163 a_989_24944# single_10b_cdac_1.cdac_sw_16_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8164 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8165 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8166 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8167 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8168 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8169 single_10b_cdac_1.cdac_sw_2_0.x2.swp single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8170 single_10b_cdac_1.x6[4].x2.swn single_10b_cdac_1.x6[4].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8171 single_10b_cdac_1.x8[6].x3.ck single_10b_cdac_1.x8[6].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8172 VSREF single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8173 a_44150_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8174 VSREF single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8175 VSREF SWN_IN[4] a_14654_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8176 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8177 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x8.A single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8178 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8179 VDREF single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8180 single_10b_cdac_1.x3[0].x3.ck single_10b_cdac_1.x3[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8181 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8182 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8183 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8184 single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8185 VDREF single_10b_cdac_1.x3[0].x1.x7.A single_10b_cdac_1.x3[0].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8186 single_10b_cdac_1.cdac_sw_1_1.x1.x8.A single_10b_cdac_1.cdac_sw_1_1.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8187 single_10b_cdac_1.cdac_sw_8_1.x1.x5.A single_10b_cdac_1.cdac_sw_8_1.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8188 VCM single_10b_cdac_1.cdac_sw_4_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8189 a_10556_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8190 a_35954_34963# SWP_IN[9] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8191 single_10b_cdac_1.cdac_sw_1_1.x1.x7.A single_10b_cdac_1.cdac_sw_1_1.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8192 VSREF single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8193 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8194 VCM single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8195 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8196 VSREF CF[6] single_10b_cdac_0.x8[6].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8197 single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8198 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8199 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8200 VSREF single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8201 single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8202 single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8203 VDREF single_10b_cdac_0.x3[0].x1.x5.A single_10b_cdac_0.x3[0].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8204 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8205 single_10b_cdac_0.cdac_sw_1_1.x1.x7.A single_10b_cdac_0.cdac_sw_1_1.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8206 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8207 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8208 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8209 VDREF single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8210 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8211 VDREF SWP_IN[8] a_6458_34754# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8212 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8213 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8214 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8215 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8216 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8217 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8218 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8219 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8220 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8221 single_10b_cdac_1.x4[2].x2.swn single_10b_cdac_1.x4[2].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8222 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8223 single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8224 single_10b_cdac_0.cdac_sw_1_1.x1.x10.A single_10b_cdac_0.cdac_sw_1_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8225 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8226 VDREF single_10b_cdac_0.x3[1].x1.x11.A single_10b_cdac_0.x3[1].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8227 single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8228 single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8229 VSREF single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8230 single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8231 single_10b_cdac_1.cdac_sw_1_2.x2.swn single_10b_cdac_1.cdac_sw_1_2.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8232 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8233 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8234 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x10.A single_10b_cdac_1.cdac_sw_2_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8235 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8236 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8237 single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8238 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8239 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8240 VSREF CF[8] single_10b_cdac_1.x10[8].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8241 single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8242 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8243 single_10b_cdac_0.cdac_sw_8_0.x1.x9.A single_10b_cdac_0.cdac_sw_8_0.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8244 single_10b_cdac_1.x6[5].x3.ck single_10b_cdac_1.x6[5].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8245 single_10b_cdac_1.x6[4].x1.x4.A CF[4] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8246 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8247 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8248 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8249 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8250 VSREF single_10b_cdac_1.x6[4].x1.x5.A single_10b_cdac_1.x6[4].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8251 VCM single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8252 VSREF single_10b_cdac_0.x2[0].x1.x9.A single_10b_cdac_0.x2[0].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8253 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8254 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x3.ckb a_44150_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8255 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8256 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8257 single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8258 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8259 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8260 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8261 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8262 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8263 VSREF SWN_IN[2] a_8214_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8264 single_10b_cdac_1.cdac_sw_1_2.x3.ck single_10b_cdac_1.cdac_sw_1_2.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8265 a_47370_25722# SWN_IN[4] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8266 single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8267 VSREF single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8268 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8269 VDREF single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8270 single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8271 VSREF single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8272 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8273 single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8274 single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8275 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8276 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8277 a_44243_24080# single_10b_cdac_0.cdac_sw_8_0.x1.x3.Y VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8278 a_13776_25722# SWN_IN[4] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8279 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8280 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8281 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8282 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8283 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8284 VDREF single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8285 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8286 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8287 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8288 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8289 single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.cdac_sw_4_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8290 single_10b_cdac_1.x4[3].x3.ck single_10b_cdac_1.x4[3].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8291 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8292 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8293 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x8.A single_10b_cdac_1.cdac_sw_4_1.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8294 single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8295 VDREF single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8296 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8297 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8298 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8299 VDREF single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8300 VSREF single_10b_cdac_1.cdac_sw_1_2.x3.ckb single_10b_cdac_1.cdac_sw_1_2.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8301 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8302 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x11.A single_10b_cdac_1.cdac_sw_4_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8303 single_10b_cdac_1.cdac_sw_8_1.x1.x6.A single_10b_cdac_1.cdac_sw_8_1.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8304 VCM single_10b_cdac_1.cdac_sw_2_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[6] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8305 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8306 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8307 VSREF single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8308 single_10b_cdac_0.cdac_sw_2_1.x1.x10.A single_10b_cdac_0.cdac_sw_2_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8309 single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8310 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8311 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8312 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8313 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8314 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8315 VSREF single_10b_cdac_0.x10[8].x1.x11.A single_10b_cdac_0.x10[8].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8316 VDREF single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8317 single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.cdac_sw_8_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8318 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8319 VDREF single_10b_cdac_0.cdac_sw_4_0.x1.x9.A single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8320 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8321 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8322 single_10b_cdac_0.cdac_sw_1_2.x1.x10.A single_10b_cdac_0.cdac_sw_1_2.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8323 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8324 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8325 VSREF single_10b_cdac_0.x4[2].x1.x10.A single_10b_cdac_0.x4[2].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8326 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8327 single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8328 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8329 single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.cdac_sw_2_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8330 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8331 VDREF single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8332 a_16118_33146# single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8333 a_20216_25722# SWN_IN[6] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8334 VCM single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8335 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8336 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8337 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8338 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8339 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8340 single_10b_cdac_0.x10b_cap_array_0.SW[4] single_10b_cdac_0.cdac_sw_4_1.x3.ckb a_47370_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8341 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8342 single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8343 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8344 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8345 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8346 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8347 single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8348 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8349 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8350 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8351 VSREF single_10b_cdac_0.x8[7].x1.x9.A single_10b_cdac_0.x8[7].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8352 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8353 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x8.A single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8354 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8355 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8356 single_10b_cdac_0.x4[3].x2.swp single_10b_cdac_0.x4[3].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8357 VSREF single_10b_cdac_1.cdac_sw_8_1.x2.swp single_10b_cdac_1.cdac_sw_8_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8358 a_4116_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8359 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8360 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8361 VDREF single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8362 a_62592_26714# single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8363 single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8364 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8365 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8366 VSREF single_10b_cdac_1.x6[4].x1.x9.A single_10b_cdac_1.x6[4].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8367 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8368 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8369 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8370 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8371 single_10b_cdac_0.cdac_sw_1_1.x3.ck single_10b_cdac_0.cdac_sw_1_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8372 VSREF single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8373 single_10b_cdac_1.x2[0].x1.x4.A CF[1] a_4209_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8374 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8375 single_10b_cdac_0.cdac_sw_8_0.x2.swn single_10b_cdac_0.cdac_sw_8_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8376 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8377 single_10b_cdac_1.x6[5].x3.ck single_10b_cdac_1.x6[5].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8378 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8379 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8380 single_10b_cdac_1.cdac_sw_8_0.x1.x8.A single_10b_cdac_1.cdac_sw_8_0.x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8381 VSREF single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8382 VSREF single_10b_cdac_0.x6[5].x1.x9.A a_49851_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8383 a_32218_26714# single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8384 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8385 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x8.A single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8386 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8387 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8388 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x6.A single_10b_cdac_0.cdac_sw_1_2.x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8389 single_10b_cdac_0.x4[3].x2.swn single_10b_cdac_0.x4[3].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8390 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8391 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x11.A single_10b_cdac_1.cdac_sw_8_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8392 single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8393 VSREF single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8394 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8395 VDREF single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8396 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8397 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8398 VSREF single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8399 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8400 single_10b_cdac_0.cdac_sw_4_0.x1.x7.A single_10b_cdac_0.cdac_sw_4_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8401 VSREF single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8402 VSREF single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8403 a_40930_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8404 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8405 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8406 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8407 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8408 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8409 VDREF SWP_IN[2] a_25778_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8410 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8411 single_10b_cdac_0.x2[0].x1.x5.A single_10b_cdac_0.x2[0].x1.x8.A a_37803_24080# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8412 single_10b_cdac_1.x3[1].x3.ck single_10b_cdac_1.x3[1].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8413 single_10b_cdac_0.x6[4].dac_out single_10b_cdac_0.x6[4].x3.ck a_52054_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8414 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8415 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8416 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8417 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8418 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8419 single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.cdac_sw_2_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8420 VDREF single_10b_cdac_0.x3[0].x1.x9.A single_10b_cdac_0.x3[0].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8421 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8422 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8423 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8424 single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.cdac_sw_4_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8425 single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8426 VSREF single_10b_cdac_0.x6[5].x1.x6.A single_10b_cdac_0.x6[5].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8427 single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8428 single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x2[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8429 VDREF single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8430 single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8431 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8432 VSREF single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8433 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8434 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8435 single_10b_cdac_1.cdac_sw_4_1.x1.x6.A single_10b_cdac_1.cdac_sw_4_1.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8436 single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8437 VSREF single_10b_cdac_1.x8[7].x1.x9.A a_9817_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8438 single_10b_cdac_0.x10b_cap_array_0.SW[6] single_10b_cdac_0.cdac_sw_2_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8439 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8440 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8441 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8442 single_10b_cdac_1.x10b_cap_array_0.SW[5] single_10b_cdac_1.cdac_sw_4_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8443 VCM single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8444 single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8445 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8446 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8447 VSREF single_10b_cdac_1.x3[0].x1.x11.A single_10b_cdac_1.x3[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8448 VSREF single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8449 single_10b_cdac_0.x10b_cap_array_0.SW[5] single_10b_cdac_0.cdac_sw_4_0.x3.ckb a_50590_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8450 VSREF single_10b_cdac_0.x2[0].x1.x11.A single_10b_cdac_0.x2[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8451 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8452 single_10b_cdac_0.x8[6].x2.swn single_10b_cdac_0.x8[6].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8453 VDREF single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8454 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8455 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8456 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8457 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8458 VCP single_10b_cdac_1.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8459 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8460 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8461 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8462 VDREF CF[0] single_10b_cdac_1.x3[0].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8463 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8464 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8465 VSREF single_10b_cdac_0.x6[4].x1.x8.A single_10b_cdac_0.x6[4].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8466 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8467 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8468 a_56152_31002# single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8469 a_24900_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8470 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8471 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8472 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8473 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8474 VDREF single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8475 VSREF single_10b_cdac_1.x8[7].x1.x9.A single_10b_cdac_1.x8[7].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8476 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8477 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8478 VDREF single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8479 VSREF single_10b_cdac_1.x8[7].x1.x6.A single_10b_cdac_1.x8[7].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8480 VCM single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8481 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x9.A single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8482 single_10b_cdac_0.cdac_sw_1_0.x3.ck single_10b_cdac_0.cdac_sw_1_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8483 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8484 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8485 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8486 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8487 a_11434_25713# single_10b_cdac_1.cdac_sw_8_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8488 a_16257_35702# CF[5] single_10b_cdac_1.x6[5].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8489 single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x2[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8490 single_10b_cdac_0.cdac_sw_16_0.x1.x5.A single_10b_cdac_0.cdac_sw_16_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8491 VDREF single_10b_cdac_0.x4[3].x1.x10.A single_10b_cdac_0.x4[3].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8492 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8493 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8494 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8495 single_10b_cdac_1.cdac_sw_1_0.x1.x6.A single_10b_cdac_1.cdac_sw_1_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8496 a_59511_36566# single_10b_cdac_0.x4[2].x1.x8.A single_10b_cdac_0.x4[2].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8497 VSREF single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8498 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8499 single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8500 single_10b_cdac_0.x6[4].x3.ck single_10b_cdac_0.x6[4].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8501 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8502 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x8.A single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8503 VDREF single_10b_cdac_1.x8[7].x2.swp single_10b_cdac_1.x8[7].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8504 single_10b_cdac_0.x6[5].x2.swn single_10b_cdac_0.x6[5].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8505 VDREF single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8506 single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8507 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8508 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8509 single_10b_cdac_1.cdac_sw_1_0.x2.swn single_10b_cdac_1.cdac_sw_1_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8510 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8511 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8512 VCN single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8513 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8514 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8515 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8516 single_10b_cdac_0.cdac_sw_1_0.x1.x9.A single_10b_cdac_0.cdac_sw_1_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8517 single_10b_cdac_1.cdac_sw_8_1.x3.ckb single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8518 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8519 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x10.A single_10b_cdac_0.cdac_sw_4_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8520 VSREF single_10b_cdac_1.cdac_sw_2_0.x3.ckb single_10b_cdac_1.cdac_sw_2_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8521 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8522 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8523 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8524 VDREF single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8525 VSREF single_10b_cdac_1.x4[3].x1.x3.Y a_22697_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8526 VSREF single_10b_cdac_0.x3[0].x1.x9.A single_10b_cdac_0.x3[0].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8527 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8528 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8529 VDREF single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8530 single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8531 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8532 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8533 VDREF single_10b_cdac_0.x4[3].x3.ckb single_10b_cdac_0.x4[3].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8534 a_7336_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8535 single_10b_cdac_0.x2[0].x1.x4.A single_10b_cdac_0.x2[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8536 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8537 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8538 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8539 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8540 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8541 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8542 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8543 single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8544 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8545 single_10b_cdac_1.x8[7].x2.swn single_10b_cdac_1.x8[7].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8546 VSREF single_10b_cdac_0.x8[7].x1.x10.A single_10b_cdac_0.x8[7].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8547 single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.cdac_sw_4_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8548 single_10b_cdac_1.cdac_sw_2_1.x1.x11.A single_10b_cdac_1.cdac_sw_2_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8549 single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x2[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8550 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8551 VSREF single_10b_cdac_1.x4[2].x1.x11.A single_10b_cdac_1.x4[2].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8552 single_10b_cdac_0.x3[0].x2.swn single_10b_cdac_0.x3[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8553 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8554 VSREF SWN_IN[3] a_45028_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8555 VSREF single_10b_cdac_1.x4[3].x1.x7.A single_10b_cdac_1.x4[3].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8556 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8557 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8558 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8559 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8560 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8561 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x9.A single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8562 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8563 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8564 single_10b_cdac_0.x2[0].x3.ckb single_10b_cdac_0.x2[0].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8565 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8566 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8567 VSREF single_10b_cdac_0.x8[6].x1.x8.A single_10b_cdac_0.x8[6].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8568 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8569 single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.cdac_sw_4_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8570 VSREF single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8571 single_10b_cdac_0.x4[3].x1.x11.A single_10b_cdac_0.x4[3].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8572 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8573 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8574 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x9.A single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8575 a_53903_24944# single_10b_cdac_0.cdac_sw_2_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8576 VDREF single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8577 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8578 VCM single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[7] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8579 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8580 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8581 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8582 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8583 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8584 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8585 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8586 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8587 single_10b_cdac_1.x8[7].dac_out single_10b_cdac_1.x8[7].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8588 a_58494_32737# SWP_IN[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8589 VCM single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8590 single_10b_cdac_0.x3[0].x2.swn single_10b_cdac_0.x3[0].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8591 VDREF single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8592 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8593 single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8594 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8595 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8596 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8597 single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.cdac_sw_16_0.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8598 single_10b_cdac_1.cdac_sw_1_1.x1.x3.Y CF[8] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8599 VSREF SWN_IN[1] a_4994_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8600 single_10b_cdac_1.cdac_sw_1_0.x1.x5.A single_10b_cdac_1.cdac_sw_1_0.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8601 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8602 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8603 single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8604 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8605 single_10b_cdac_1.cdac_sw_2_1.x1.x3.Y CF[6] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8606 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8607 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8608 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8609 VSREF SWN_IN[0] a_1774_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8610 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8611 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8612 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8613 a_35368_25713# single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8614 a_38588_25713# single_10b_cdac_0.x2[0].x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8615 single_10b_cdac_0.cdac_sw_2_1.x3.ckb single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8616 VDREF CF[9] single_10b_cdac_1.cdac_sw_1_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8617 VSREF single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8618 VDREF single_10b_cdac_0.x4[2].x1.x5.A single_10b_cdac_0.x4[2].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8619 VCM single_10b_cdac_1.cdac_sw_16_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8620 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8621 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8622 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8623 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8624 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8625 VDREF single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8626 VSREF single_10b_cdac_1.x2[0].x2.swp single_10b_cdac_1.x2[0].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8627 single_10b_cdac_0.x3[1].x3.ck single_10b_cdac_0.x3[1].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8628 a_59372_31002# single_10b_cdac_0.x4[2].x3.ckb single_10b_cdac_0.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8629 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8630 VSREF single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8631 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8632 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8633 VDREF single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8634 single_10b_cdac_1.x8[6].x3.ck single_10b_cdac_1.x8[6].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8635 VDREF single_10b_cdac_0.x6[5].x1.x8.A single_10b_cdac_0.x6[5].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8636 VSREF single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8637 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8638 single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.cdac_sw_8_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8639 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8640 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8641 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8642 single_10b_cdac_1.cdac_sw_4_1.x1.x11.A single_10b_cdac_1.cdac_sw_4_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8643 VSREF single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8644 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8645 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8646 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8647 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8648 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8649 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8650 single_10b_cdac_1.x4[3].dac_out single_10b_cdac_1.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8651 single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8652 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8653 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8654 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8655 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8656 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8657 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8658 VDREF single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8659 single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8660 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8661 single_10b_cdac_1.cdac_sw_4_0.x2.swn single_10b_cdac_1.cdac_sw_4_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8662 single_10b_cdac_1.cdac_sw_1_2.x1.x5.A single_10b_cdac_1.cdac_sw_1_2.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8663 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x3.ck a_61714_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8664 VDREF SWP_IN[3] a_22558_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8665 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8666 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8667 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8668 VDREF single_10b_cdac_1.x8[7].x3.ckb single_10b_cdac_1.x8[7].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8669 single_10b_cdac_0.x6[5].x3.ck single_10b_cdac_0.x6[5].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8670 single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8671 VSREF single_10b_cdac_1.cdac_sw_8_1.x1.x9.A single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8672 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8673 VSREF single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8674 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8675 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8676 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8677 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8678 VCM single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8679 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8680 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8681 VSREF single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8682 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8683 single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8684 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8685 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8686 VSREF single_10b_cdac_1.x4[3].x1.x9.A single_10b_cdac_1.x4[3].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8687 single_10b_cdac_1.cdac_sw_1_2.x3.ck single_10b_cdac_1.cdac_sw_1_2.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8688 single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8689 single_10b_cdac_0.x4[2].x2.swn single_10b_cdac_0.x4[2].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8690 single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8691 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x8.A single_10b_cdac_0.cdac_sw_2_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8692 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8693 VDREF single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8694 VDREF SWP_IN[5] a_49712_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8695 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8696 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8697 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8698 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8699 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8700 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x10.A single_10b_cdac_0.cdac_sw_2_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8701 single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8702 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8703 single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8704 a_43411_36566# single_10b_cdac_0.x8[7].x1.x8.A single_10b_cdac_0.x8[7].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8705 VCN single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8706 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8707 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8708 VSREF SWN_IN[5] a_17874_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8709 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8710 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8711 single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8712 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8713 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8714 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8715 VSREF SWN_IN[2] a_8214_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8716 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8717 VSREF single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8718 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8719 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8720 VDREF single_10b_cdac_1.x6[4].x2.swp single_10b_cdac_1.x6[4].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8721 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8722 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8723 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8724 single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8725 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8726 VSREF single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8727 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8728 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x8.A single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8729 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8730 single_10b_cdac_0.x3[1].x2.swp single_10b_cdac_0.x3[1].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8731 VCM single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[6] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8732 single_10b_cdac_1.x2[0].x1.x11.A single_10b_cdac_1.x2[0].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8733 VSREF single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8734 a_8800_34645# SWP_IN[7] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8735 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8736 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8737 VCM single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8738 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8739 single_10b_cdac_1.cdac_sw_2_0.x1.x9.A single_10b_cdac_1.cdac_sw_2_0.x1.x7.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8740 single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8741 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8742 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8743 VCP single_10b_cdac_0.x3[1].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8744 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8745 single_10b_cdac_0.x8[6].x1.x5.A single_10b_cdac_0.x8[6].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8746 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8747 VCP single_10b_cdac_1.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8748 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8749 single_10b_cdac_0.cdac_sw_1_1.x2.swp single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8750 VDREF single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8751 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8752 single_10b_cdac_0.cdac_sw_1_0.x1.x11.A single_10b_cdac_0.cdac_sw_1_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8753 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8754 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8755 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8756 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8757 single_10b_cdac_0.cdac_sw_4_0.x1.x8.A single_10b_cdac_0.cdac_sw_4_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8758 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8759 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8760 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8761 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8762 single_10b_cdac_1.x10b_cap_array_0.SW[5] single_10b_cdac_1.cdac_sw_4_0.x3.ckb a_16996_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8763 VSREF single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8764 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x3.ckb a_40930_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8765 single_10b_cdac_0.cdac_sw_1_0.x2.swn single_10b_cdac_0.cdac_sw_1_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8766 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8767 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x8.A single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8768 single_10b_cdac_1.cdac_sw_8_1.x1.x10.A single_10b_cdac_1.cdac_sw_8_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8769 a_25778_31002# single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8770 VSREF SWN_IN[2] a_41808_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8771 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8772 VDREF single_10b_cdac_1.x8[7].x1.x11.A single_10b_cdac_1.x8[7].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8773 a_52054_34009# SWP_IN[4] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8774 single_10b_cdac_0.x6[5].x2.swp single_10b_cdac_0.x6[5].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8775 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8776 VDREF single_10b_cdac_1.x2[0].x1.x9.A single_10b_cdac_1.x2[0].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8777 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8778 single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8779 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8780 VSREF single_10b_cdac_1.x3[0].x1.x8.A single_10b_cdac_1.x3[0].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8781 VCM single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8782 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8783 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8784 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8785 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8786 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8787 VDREF single_10b_cdac_1.x3[1].x1.x9.A single_10b_cdac_1.x3[1].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8788 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8789 VCP single_10b_cdac_1.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8790 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8791 single_10b_cdac_0.cdac_sw_1_0.x3.ck single_10b_cdac_0.cdac_sw_1_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8792 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8793 a_62731_36566# single_10b_cdac_0.x3[1].x1.x8.A single_10b_cdac_0.x3[1].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8794 a_42394_34645# SWP_IN[7] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8795 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8796 a_10556_25722# SWN_IN[3] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8797 single_10b_cdac_0.cdac_sw_2_1.x3.ck single_10b_cdac_0.cdac_sw_2_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8798 single_10b_cdac_1.cdac_sw_1_1.x1.x4.A CF[8] a_26749_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8799 VCM single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8800 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8801 VDREF single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8802 single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8803 a_21680_32737# SWP_IN[3] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8804 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8805 a_49712_33146# single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8806 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8807 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8808 single_10b_cdac_1.cdac_sw_8_0.x1.x3.Y CF[3] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8809 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8810 single_10b_cdac_1.cdac_sw_4_1.x1.x5.A single_10b_cdac_1.cdac_sw_4_1.x1.x3.Y VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8811 VSREF single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8812 single_10b_cdac_0.x10b_cap_array_0.SW[2] single_10b_cdac_0.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8813 VDREF SWP_IN[1] a_62592_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8814 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8815 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8816 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8817 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8818 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8819 VDREF single_10b_cdac_1.cdac_sw_8_1.x1.x8.A single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8820 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8821 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8822 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8823 single_10b_cdac_0.cdac_sw_8_0.x1.x7.A single_10b_cdac_0.cdac_sw_8_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8824 VSREF single_10b_cdac_0.cdac_sw_1_0.x1.x8.A single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8825 VDREF single_10b_cdac_0.x6[5].x1.x11.A single_10b_cdac_0.x6[5].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8826 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8827 VSREF single_10b_cdac_0.cdac_sw_2_0.x2.swp single_10b_cdac_0.cdac_sw_2_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8828 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x9.A single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8829 VDREF single_10b_cdac_0.x8[7].x1.x5.A single_10b_cdac_0.x8[7].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8830 VSREF single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8831 single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8832 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8833 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8834 VDREF SWP_IN[1] a_28998_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8835 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8836 a_896_25722# SWN_IN[0] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8837 a_43272_34218# single_10b_cdac_0.x8[7].x3.ckb single_10b_cdac_0.x8[7].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8838 VSREF single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8839 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8840 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8841 VDREF SWP_IN[2] a_59372_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8842 single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8843 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8844 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8845 VSREF single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8846 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8847 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8848 VCP single_10b_cdac_1.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8849 single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8850 single_10b_cdac_0.cdac_sw_2_0.x1.x11.A single_10b_cdac_0.cdac_sw_2_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8851 single_10b_cdac_0.x10b_cap_array_0.SW[4] single_10b_cdac_0.cdac_sw_4_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8852 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8853 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8854 single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8855 VDREF single_10b_cdac_1.x6[4].x1.x6.A single_10b_cdac_1.x6[4].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8856 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8857 VSREF single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8858 single_10b_cdac_1.x2[0].x1.x8.A single_10b_cdac_1.x2[0].x1.x6.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8859 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x3.ckb a_44150_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8860 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8861 single_10b_cdac_0.cdac_sw_4_1.x1.x6.A single_10b_cdac_0.cdac_sw_4_1.x1.x4.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8862 VDREF single_10b_cdac_0.cdac_sw_1_0.x1.x8.A single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8863 single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8864 VSREF single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8865 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8866 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8867 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8868 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8869 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8870 single_10b_cdac_1.x2[0].x1.x7.A single_10b_cdac_1.x2[0].x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8871 single_10b_cdac_1.cdac_sw_16_0.x3.ckb single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8872 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x3.ck a_55274_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8873 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8874 single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.cdac_sw_2_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8875 single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8876 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8877 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8878 VSREF single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8879 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8880 VDREF CF[2] single_10b_cdac_1.x4[2].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8881 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8882 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x3.ck a_28120_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8883 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8884 single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8885 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8886 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8887 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8888 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8889 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8890 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8891 single_10b_cdac_1.cdac_sw_4_0.x3.ckb single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8892 a_48248_25713# single_10b_cdac_0.cdac_sw_4_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8893 VSREF single_10b_cdac_1.x4[2].x1.x8.A single_10b_cdac_1.x4[2].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8894 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8895 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8896 single_10b_cdac_0.cdac_sw_2_0.x3.ck single_10b_cdac_0.cdac_sw_2_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8897 VSREF single_10b_cdac_1.cdac_sw_4_0.x1.x9.A single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8898 VDREF single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8899 VDREF SWP_IN[2] a_25778_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8900 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x3.ck a_24900_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8901 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8902 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8903 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8904 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8905 VSREF single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8906 a_57030_25722# SWN_IN[7] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8907 single_10b_cdac_0.x8[7].x2.swn single_10b_cdac_0.x8[7].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8908 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8909 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8910 a_4209_24944# single_10b_cdac_1.x2[0].x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8911 VDREF single_10b_cdac_0.x6[5].x1.x10.A single_10b_cdac_0.x6[5].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8912 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x8.A single_10b_cdac_0.cdac_sw_8_1.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8913 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8914 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8915 VSREF single_10b_cdac_1.x10[8].x3.ckb single_10b_cdac_1.x10[8].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8916 single_10b_cdac_0.x8[6].x3.ck single_10b_cdac_0.x8[6].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8917 a_45028_25713# single_10b_cdac_0.cdac_sw_8_0.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8918 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8919 single_10b_cdac_1.x3[1].x2.swn single_10b_cdac_1.x3[1].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8920 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8921 VDREF single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8922 single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8923 single_10b_cdac_0.cdac_sw_1_0.x1.x6.A single_10b_cdac_0.cdac_sw_1_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8924 a_41808_25713# single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8925 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x10.A single_10b_cdac_1.cdac_sw_16_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8926 single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8927 single_10b_cdac_1.x6[4].x2.swn single_10b_cdac_1.x6[4].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8928 a_31340_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8929 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8930 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8931 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8932 single_10b_cdac_1.x10b_cap_array_0.SW[3] single_10b_cdac_1.cdac_sw_8_0.x3.ckb a_10556_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8933 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8934 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8935 single_10b_cdac_0.cdac_sw_1_0.x2.swn single_10b_cdac_0.cdac_sw_1_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8936 single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8937 single_10b_cdac_1.x8[6].x3.ckb single_10b_cdac_1.x8[6].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8938 VDREF single_10b_cdac_0.x10[8].x1.x7.A single_10b_cdac_0.x10[8].x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8939 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x11.A single_10b_cdac_1.cdac_sw_1_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8940 VSREF single_10b_cdac_1.x6[5].x1.x3.Y a_16257_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8941 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8942 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8943 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8944 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8945 VSREF single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8946 VDREF single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8947 VSREF single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8948 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8949 VDREF CF[3] single_10b_cdac_0.cdac_sw_8_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8950 VCP single_10b_cdac_1.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8951 VDREF single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8952 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8953 VCP single_10b_cdac_1.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8954 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x8.A single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8955 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8956 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8957 a_9817_35702# CF[7] single_10b_cdac_1.x8[7].x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8958 a_4994_25713# single_10b_cdac_1.x2[0].x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8959 single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8960 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8961 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8962 VDREF single_10b_cdac_1.x3[1].x1.x8.A single_10b_cdac_1.x3[1].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8963 a_1774_25713# single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8964 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8965 VDREF single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8966 VSREF single_10b_cdac_1.x6[4].x1.x11.A single_10b_cdac_1.x6[4].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8967 single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8968 single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.cdac_sw_2_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8969 single_10b_cdac_1.x10[8].x1.x11.A single_10b_cdac_1.x10[8].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8970 single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8971 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8972 single_10b_cdac_0.cdac_sw_2_1.x1.x11.A single_10b_cdac_0.cdac_sw_2_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8973 single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8974 VDREF single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8975 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x3.ckb a_896_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8976 VCN single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8977 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8978 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8979 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8980 VSREF single_10b_cdac_0.x4[3].x1.x7.A single_10b_cdac_0.x4[3].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8981 VSREF single_10b_cdac_0.x10[8].x1.x8.A single_10b_cdac_0.x10[8].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8982 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8983 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8984 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8985 single_10b_cdac_1.cdac_sw_4_0.x1.x7.A single_10b_cdac_1.cdac_sw_4_0.x1.x5.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8986 VDREF single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8987 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8988 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8989 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x3.ck a_64934_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8990 single_10b_cdac_1.x3[1].dac_out single_10b_cdac_1.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8991 single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.cdac_sw_4_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8992 a_47463_24944# single_10b_cdac_0.cdac_sw_4_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8993 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8994 single_10b_cdac_0.cdac_sw_1_1.x1.x4.A CF[8] a_60343_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8995 VDREF single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8996 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8997 single_10b_cdac_0.cdac_sw_4_0.x2.swp single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8998 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8999 single_10b_cdac_1.cdac_sw_4_0.x1.x10.A single_10b_cdac_1.cdac_sw_4_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9000 VSREF single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9001 single_10b_cdac_0.x3[0].dac_out single_10b_cdac_0.x3[0].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9002 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9003 single_10b_cdac_0.x4[2].x2.swn single_10b_cdac_0.x4[2].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9004 single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.cdac_sw_2_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9005 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9006 VDREF single_10b_cdac_1.x8[6].x1.x9.A single_10b_cdac_1.x8[6].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9007 single_10b_cdac_0.x10[8].x3.ck single_10b_cdac_0.x10[8].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9008 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9009 single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9010 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9011 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9012 single_10b_cdac_1.x8[7].x2.swn single_10b_cdac_1.x8[7].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9013 single_10b_cdac_1.cdac_sw_8_0.x1.x4.A CF[3] a_10649_24944# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9014 VSREF single_10b_cdac_0.x10[8].x1.x5.A single_10b_cdac_0.x10[8].x1.x7.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9015 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9016 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9017 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9018 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9019 a_61714_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9020 a_65812_26714# single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9021 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9022 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9023 single_10b_cdac_0.cdac_sw_2_1.x1.x3.Y CF[6] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9024 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9025 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9026 a_22697_36566# single_10b_cdac_1.x4[3].x1.x8.A single_10b_cdac_1.x4[3].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9027 VDREF CF[9] single_10b_cdac_0.cdac_sw_1_0.x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9028 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9029 VDREF single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9030 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9031 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9032 VSREF single_10b_cdac_0.cdac_sw_8_1.x2.swp single_10b_cdac_0.cdac_sw_8_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9033 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9034 single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9035 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9036 VSREF single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9037 VDREF single_10b_cdac_0.x4[2].x2.swp single_10b_cdac_0.x4[2].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9038 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9039 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9040 single_10b_cdac_0.cdac_sw_16_0.x3.ck single_10b_cdac_0.cdac_sw_16_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9041 VSREF single_10b_cdac_1.x3[0].x1.x10.A single_10b_cdac_1.x3[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9042 VSREF single_10b_cdac_0.cdac_sw_4_1.x3.ckb single_10b_cdac_0.cdac_sw_4_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9043 VDREF single_10b_cdac_0.x3[1].x1.x9.A single_10b_cdac_0.x3[1].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9044 single_10b_cdac_1.x10b_cap_array_0.SW[0] single_10b_cdac_1.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9045 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9046 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9047 single_10b_cdac_0.x6[5].x2.swn single_10b_cdac_0.x6[5].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9048 single_10b_cdac_0.x4[3].dac_out single_10b_cdac_0.x4[3].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9049 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9050 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9051 VSREF single_10b_cdac_1.cdac_sw_4_0.x2.swp single_10b_cdac_1.cdac_sw_4_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9052 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x9.A single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9053 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9054 single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.cdac_sw_8_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9055 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x10.A single_10b_cdac_1.cdac_sw_1_2.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9056 VCM single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9057 a_17874_25713# single_10b_cdac_1.cdac_sw_4_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9058 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9059 single_10b_cdac_1.x6[5].dac_out single_10b_cdac_1.x6[5].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9060 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9061 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9062 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9063 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9064 single_10b_cdac_0.cdac_sw_8_1.x1.x11.A single_10b_cdac_0.cdac_sw_8_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9065 VDREF single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9066 single_10b_cdac_1.x4[3].x2.swn single_10b_cdac_1.x4[3].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9067 single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9068 VDREF SWP_IN[5] a_16118_33146# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9069 single_10b_cdac_1.x10b_cap_array_0.SW[6] single_10b_cdac_1.cdac_sw_2_1.x3.ckb a_20216_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9070 VDREF single_10b_cdac_1.x3[0].x3.ckb single_10b_cdac_1.x3[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9071 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9072 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9073 VSREF single_10b_cdac_1.x8[6].x2.swp single_10b_cdac_1.x8[6].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9074 single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9075 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9076 single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.cdac_sw_8_1.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9077 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9078 single_10b_cdac_1.cdac_sw_1_0.x1.x8.A single_10b_cdac_1.cdac_sw_1_0.x1.x6.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9079 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9080 VDREF CF[7] single_10b_cdac_1.x8[7].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9081 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9082 single_10b_cdac_1.cdac_sw_8_0.x3.ckb single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9083 single_10b_cdac_0.x4[3].x3.ck single_10b_cdac_0.x4[3].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9084 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9085 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9086 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9087 VDREF single_10b_cdac_1.x3[0].x1.x9.A single_10b_cdac_1.x3[0].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9088 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9089 single_10b_cdac_0.x10b_cap_array_0.SW[3] single_10b_cdac_0.cdac_sw_8_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9090 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9091 VDREF single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9092 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9093 VSREF single_10b_cdac_1.x6[5].x1.x6.A single_10b_cdac_1.x6[5].x1.x8.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9094 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9095 single_10b_cdac_0.cdac_sw_8_1.x3.ck single_10b_cdac_0.cdac_sw_8_1.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9096 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x3.ckb a_4116_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9097 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9098 a_40930_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9099 single_10b_cdac_1.x10b_cap_array_0.SW[6] single_10b_cdac_1.cdac_sw_2_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9100 single_10b_cdac_1.cdac_sw_16_0.x1.x11.A single_10b_cdac_1.cdac_sw_16_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9101 single_10b_cdac_0.cdac_sw_1_0.x3.ckb single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9102 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9103 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9104 single_10b_cdac_0.cdac_sw_4_1.x2.swp single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9105 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9106 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9107 VSREF single_10b_cdac_0.x6[5].x1.x4.A single_10b_cdac_0.x6[5].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9108 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9109 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9110 single_10b_cdac_1.x8[6].x2.swn single_10b_cdac_1.x8[6].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9111 single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9112 a_16996_25722# SWN_IN[5] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9113 VSREF single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9114 VDREF single_10b_cdac_0.x6[4].x1.x11.A single_10b_cdac_0.x6[4].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9115 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9116 single_10b_cdac_1.x2[0].x2.swn single_10b_cdac_1.x2[0].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9117 VDREF SWP_IN[0] a_32218_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9118 single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9119 a_28120_30193# SWP_IN[1] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9120 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x11.A single_10b_cdac_1.cdac_sw_8_0.x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9121 VSREF single_10b_cdac_0.x8[6].x1.x10.A single_10b_cdac_0.x8[6].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9122 single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9123 single_10b_cdac_1.x10b_cap_array_0.SW[1] single_10b_cdac_1.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9124 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9125 VSREF single_10b_cdac_1.x3[1].x1.x11.A single_10b_cdac_1.x3[1].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9126 single_10b_cdac_1.cdac_sw_16_0.x3.ck single_10b_cdac_1.cdac_sw_16_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9127 VDREF single_10b_cdac_1.x4[3].x1.x5.A single_10b_cdac_1.x4[3].x1.x7.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9128 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9129 VCM single_10b_cdac_0.cdac_sw_4_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[4] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9130 VSREF single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9131 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9132 VDREF single_10b_cdac_0.x2[0].x2.swp single_10b_cdac_0.x2[0].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9133 VCM single_10b_cdac_1.x3[1].x2.swp single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9134 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9135 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9136 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9137 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9138 a_8214_25713# single_10b_cdac_1.cdac_sw_8_1.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9139 a_22558_31002# single_10b_cdac_1.x4[3].x3.ckb single_10b_cdac_1.x4[3].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9140 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9141 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9142 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9143 single_10b_cdac_1.cdac_sw_1_1.x2.swn single_10b_cdac_1.cdac_sw_1_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9144 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9145 VDREF single_10b_cdac_0.x6[4].x1.x3.Y single_10b_cdac_0.x6[4].x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9146 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9147 single_10b_cdac_1.cdac_sw_1_0.x2.swp single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9148 single_10b_cdac_0.x3[0].x1.x10.A single_10b_cdac_0.x3[0].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9149 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9150 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9151 single_10b_cdac_1.x6[5].x2.swn single_10b_cdac_1.x6[5].x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9152 single_10b_cdac_0.cdac_sw_2_1.x2.swp single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9153 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9154 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9155 VDREF single_10b_cdac_1.x8[6].x1.x8.A single_10b_cdac_1.x8[6].x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9156 single_10b_cdac_0.x6[5].dac_out single_10b_cdac_0.x6[5].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9157 a_40930_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9158 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9159 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9160 single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9161 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x8.A single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9162 single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.cdac_sw_16_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9163 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x10.A single_10b_cdac_1.cdac_sw_4_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9164 single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9165 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9166 single_10b_cdac_0.x8[6].x3.ckb single_10b_cdac_0.x8[6].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9167 a_28998_26714# single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9168 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9169 VDREF single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9170 VDREF single_10b_cdac_1.cdac_sw_1_1.x1.x9.A single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9171 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9172 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9173 VCM single_10b_cdac_1.cdac_sw_8_1.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9174 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9175 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9176 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9177 VDREF single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9178 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9179 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9180 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9181 VSREF single_10b_cdac_1.x4[2].x1.x8.A single_10b_cdac_1.x4[2].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9182 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9183 VDREF single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9184 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9185 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9186 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9187 single_10b_cdac_0.cdac_sw_2_0.x3.ckb single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9188 a_24314_25713# single_10b_cdac_1.cdac_sw_2_0.x3.ck single_10b_cdac_1.x10b_cap_array_0.SW[7] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9189 VSREF single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9190 VCM single_10b_cdac_1.x4[2].x2.swp single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9191 single_10b_cdac_1.x4[2].dac_out single_10b_cdac_1.x4[2].x3.ck a_24900_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9192 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9193 VSREF single_10b_cdac_1.cdac_sw_2_0.x1.x11.A single_10b_cdac_1.cdac_sw_2_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9194 single_10b_cdac_0.cdac_sw_16_0.x2.swp single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9195 single_10b_cdac_1.cdac_sw_1_2.x2.swn single_10b_cdac_1.cdac_sw_1_2.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9196 a_15240_34009# SWP_IN[5] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9197 single_10b_cdac_0.x3[0].x3.ck single_10b_cdac_0.x3[0].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9198 a_7336_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9199 VSREF SWN_IN[3] a_11434_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9200 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9201 single_10b_cdac_0.cdac_sw_8_1.x1.x10.A single_10b_cdac_0.cdac_sw_8_1.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9202 VDREF single_10b_cdac_1.x3[1].x1.x10.A single_10b_cdac_1.x3[1].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9203 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9204 VDREF SWP_IN[3] a_56152_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9205 single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9206 VCM single_10b_cdac_0.cdac_sw_4_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[5] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9207 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9208 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9209 VSREF single_10b_cdac_1.cdac_sw_1_0.x1.x10.A single_10b_cdac_1.cdac_sw_1_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9210 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9211 VCN single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9212 VCN single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9213 single_10b_cdac_0.cdac_sw_8_0.x1.x3.Y CF[3] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9214 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9215 single_10b_cdac_0.x2[0].x1.x6.A single_10b_cdac_0.x2[0].x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9216 VDREF single_10b_cdac_1.cdac_sw_2_1.x1.x10.A single_10b_cdac_1.cdac_sw_2_1.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9217 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9218 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9219 single_10b_cdac_1.x4[3].x1.x11.A single_10b_cdac_1.x4[3].x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9220 VDREF single_10b_cdac_1.x2[0].x3.ckb single_10b_cdac_1.x2[0].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9221 VSREF single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9222 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x3.ckb a_37710_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9223 single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9224 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9225 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9226 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9227 VCM single_10b_cdac_0.cdac_sw_8_1.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9228 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9229 VCM single_10b_cdac_1.cdac_sw_2_0.x2.swn single_10b_cdac_1.x10b_cap_array_0.SW[7] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9230 a_25778_31002# single_10b_cdac_1.x4[2].x3.ckb single_10b_cdac_1.x4[2].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9231 single_10b_cdac_0.x6[4].x3.ckb single_10b_cdac_0.x6[4].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9232 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9233 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9234 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9235 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9236 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9237 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9238 VSREF CF[3] single_10b_cdac_0.x4[3].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9239 a_36971_35702# CF[9] single_10b_cdac_0.cdac_sw_1_2.x1.x4.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9240 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9241 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9242 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9243 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9244 VDREF single_10b_cdac_0.x8[7].x2.swp single_10b_cdac_0.x8[7].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9245 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x3.ckb a_7336_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9246 VSREF single_10b_cdac_0.cdac_sw_16_0.x1.x11.A single_10b_cdac_0.cdac_sw_16_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9247 VSREF single_10b_cdac_1.cdac_sw_1_2.x2.swp single_10b_cdac_1.cdac_sw_1_2.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9248 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9249 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9250 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9251 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9252 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9253 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9254 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9255 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9256 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9257 VDREF single_10b_cdac_1.cdac_sw_1_2.x1.x7.A single_10b_cdac_1.cdac_sw_1_2.x1.x9.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9258 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9259 VCP single_10b_cdac_1.x4[3].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9260 VDREF single_10b_cdac_0.cdac_sw_2_0.x1.x8.A single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9261 single_10b_cdac_0.x3[0].x3.ckb single_10b_cdac_0.x3[0].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9262 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9263 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9264 single_10b_cdac_0.x6[5].dac_out single_10b_cdac_0.x6[5].x3.ck a_48834_34009# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9265 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9266 VDREF single_10b_cdac_0.cdac_sw_1_1.x3.ckb single_10b_cdac_0.cdac_sw_1_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9267 single_10b_cdac_0.x6[4].x1.x4.A CF[4] VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9268 single_10b_cdac_0.x10[8].x3.ckb single_10b_cdac_0.x10[8].x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9269 a_7336_25722# SWN_IN[2] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9270 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9271 VSREF single_10b_cdac_0.cdac_sw_1_0.x2.swp single_10b_cdac_0.cdac_sw_1_0.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9272 single_10b_cdac_0.cdac_sw_1_2.x1.x11.A single_10b_cdac_0.cdac_sw_1_2.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9273 VSREF single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9274 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9275 VDREF single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9276 VDREF single_10b_cdac_1.x6[5].x3.ckb single_10b_cdac_1.x6[5].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9277 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9278 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9279 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9280 VCN single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9281 VSREF single_10b_cdac_1.x6[4].x1.x8.A single_10b_cdac_1.x6[4].x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9282 single_10b_cdac_1.x10b_cap_array_0.SW[2] single_10b_cdac_1.cdac_sw_8_1.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9283 VDREF CF[2] single_10b_cdac_0.x4[2].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9284 VCN single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9285 single_10b_cdac_0.cdac_sw_2_1.x1.x9.A single_10b_cdac_0.cdac_sw_2_1.x1.x7.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9286 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9287 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9288 VDREF single_10b_cdac_1.x10[8].x2.swp single_10b_cdac_1.x10[8].x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9289 VSREF single_10b_cdac_1.cdac_sw_4_1.x2.swp single_10b_cdac_1.cdac_sw_4_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9290 a_26749_24944# single_10b_cdac_1.cdac_sw_1_1.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9291 VDREF SWP_IN[0] a_65812_26714# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9292 VCN single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9293 single_10b_cdac_0.x10b_cap_array_0.SW[1] single_10b_cdac_0.x2[0].x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9294 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9295 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9296 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9297 single_10b_cdac_1.cdac_sw_16_0.x2.swp single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9298 VDREF SWP_IN[2] a_59372_31002# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9299 VSREF single_10b_cdac_1.x3[1].x3.ckb single_10b_cdac_1.x3[1].x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9300 single_10b_cdac_0.x4[2].dac_out single_10b_cdac_0.x4[2].x3.ck a_58494_32737# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9301 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9302 single_10b_cdac_0.x10[8].x3.ck single_10b_cdac_0.x10[8].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9303 VDREF single_10b_cdac_0.cdac_sw_16_0.x1.x10.A single_10b_cdac_0.cdac_sw_16_0.x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9304 VCP single_10b_cdac_0.x6[4].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9305 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9306 single_10b_cdac_0.cdac_sw_2_0.x1.x6.A single_10b_cdac_0.cdac_sw_2_0.x1.x4.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9307 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9308 VDREF single_10b_cdac_0.x4[2].x1.x11.A single_10b_cdac_0.x4[2].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9309 single_10b_cdac_1.x3[0].dac_out single_10b_cdac_1.x3[0].x3.ck a_31340_30193# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9310 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9311 single_10b_cdac_0.cdac_sw_1_1.x3.ck single_10b_cdac_0.cdac_sw_1_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9312 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9313 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9314 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9315 VSREF single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9316 single_10b_cdac_0.cdac_sw_2_0.x2.swn single_10b_cdac_0.cdac_sw_2_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9317 single_10b_cdac_0.cdac_sw_1_1.x1.x11.A single_10b_cdac_0.cdac_sw_1_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9318 a_64934_30193# SWP_IN[0] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9319 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9320 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9321 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9322 VSREF SWN_IN[0] a_35368_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9323 VSREF SWN_IN[1] a_38588_25713# VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9324 single_10b_cdac_1.cdac_sw_1_1.x3.ckb single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9325 VDREF single_10b_cdac_1.x10[8].x1.x10.A single_10b_cdac_1.x10[8].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9326 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9327 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9328 VSREF single_10b_cdac_0.x8[6].x2.swp single_10b_cdac_0.x8[6].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9329 single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9330 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x11.A single_10b_cdac_0.cdac_sw_4_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9331 VSREF single_10b_cdac_0.x6[5].x1.x3.Y a_49851_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9332 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9333 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9334 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9335 single_10b_cdac_1.cdac_sw_8_0.x1.x10.A single_10b_cdac_1.cdac_sw_8_0.x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9336 VDREF single_10b_cdac_0.cdac_sw_1_2.x2.swp single_10b_cdac_0.cdac_sw_1_2.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9337 a_37710_25722# SWN_IN[1] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9338 VCM single_10b_cdac_0.x2[0].x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9339 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9340 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9341 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9342 VDREF single_10b_cdac_1.cdac_sw_1_1.x2.swp single_10b_cdac_1.cdac_sw_1_1.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9343 VDREF single_10b_cdac_1.cdac_sw_2_0.x1.x8.A single_10b_cdac_1.cdac_sw_2_0.x1.x5.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9344 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9345 VSREF single_10b_cdac_1.x8[6].x1.x11.A single_10b_cdac_1.x8[6].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9346 VSREF single_10b_cdac_1.cdac_sw_2_1.x2.swp single_10b_cdac_1.cdac_sw_2_1.x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9347 VCM single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9348 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9349 single_10b_cdac_1.x3[1].x3.ck single_10b_cdac_1.x3[1].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9350 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9351 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9352 single_10b_cdac_0.cdac_sw_16_0.x3.ckb single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9353 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9354 VSREF single_10b_cdac_0.cdac_sw_4_0.x1.x10.A single_10b_cdac_0.cdac_sw_4_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9355 VDREF single_10b_cdac_0.cdac_sw_1_2.x1.x9.A single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9356 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9357 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9358 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9359 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x2.swp VCM VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9360 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9361 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9362 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9363 single_10b_cdac_1.cdac_sw_8_0.x2.swn single_10b_cdac_1.cdac_sw_8_0.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9364 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9365 single_10b_cdac_1.x3[1].x2.swn single_10b_cdac_1.x3[1].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9366 single_10b_cdac_0.cdac_sw_1_0.x1.x10.A single_10b_cdac_0.cdac_sw_1_0.x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9367 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9368 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9369 VDREF single_10b_cdac_0.x3[0].x1.x11.A single_10b_cdac_0.x3[0].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9370 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9371 single_10b_cdac_0.cdac_sw_4_1.x1.x11.A single_10b_cdac_0.cdac_sw_4_1.x1.x9.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9372 VDREF single_10b_cdac_0.cdac_sw_1_1.x1.x9.A single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9373 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9374 VCP single_10b_cdac_0.x6[5].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9375 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9376 VSREF single_10b_cdac_0.x6[5].x1.x7.A single_10b_cdac_0.x6[5].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9377 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9378 VSREF single_10b_cdac_1.cdac_sw_1_1.x1.x10.A single_10b_cdac_1.cdac_sw_1_1.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9379 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9380 VCN single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9381 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9382 VCN single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9383 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9384 VSREF single_10b_cdac_1.x8[7].x1.x3.Y a_9817_36566# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9385 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9386 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9387 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9388 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9389 single_10b_cdac_0.cdac_sw_1_2.x2.swn single_10b_cdac_0.cdac_sw_1_2.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9390 single_10b_cdac_0.cdac_sw_8_0.x2.swp single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9391 VSREF single_10b_cdac_0.x6[4].x2.swp single_10b_cdac_0.x6[4].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9392 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9393 VDREF single_10b_cdac_1.cdac_sw_8_0.x1.x9.A single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9394 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9395 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9396 VCP single_10b_cdac_0.x8[6].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9397 VDREF single_10b_cdac_1.x6[5].x1.x4.A single_10b_cdac_1.x6[5].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9398 single_10b_cdac_0.x6[5].x3.ckb single_10b_cdac_0.x6[5].x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9399 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9400 VSREF single_10b_cdac_1.x6[4].x1.x10.A single_10b_cdac_1.x6[4].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9401 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9402 VCM single_10b_cdac_0.x3[0].x2.swp single_10b_cdac_0.x3[0].dac_out VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9403 single_10b_cdac_1.cdac_sw_4_1.x3.ck single_10b_cdac_1.cdac_sw_4_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9404 VSREF single_10b_cdac_0.x2[0].x1.x10.A single_10b_cdac_0.x2[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9405 single_10b_cdac_0.cdac_sw_4_0.x3.ckb single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9406 single_10b_cdac_1.x10[8].x3.ck single_10b_cdac_1.x10[8].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9407 VCN single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9408 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9409 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9410 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9411 VSREF single_10b_cdac_0.x6[4].x1.x9.A single_10b_cdac_0.x6[4].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9412 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9413 VDREF single_10b_cdac_1.cdac_sw_8_0.x2.swp single_10b_cdac_1.cdac_sw_8_0.x2.swn VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9414 single_10b_cdac_0.cdac_sw_8_1.x3.ckb single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9415 VSREF single_10b_cdac_0.x6[4].x1.x4.A single_10b_cdac_0.x6[4].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9416 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9417 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9418 VDREF single_10b_cdac_0.x8[6].x1.x9.A single_10b_cdac_0.x8[6].x1.x4.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9419 single_10b_cdac_1.x10[8].x3.ck single_10b_cdac_1.x10[8].x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9420 single_10b_cdac_1.cdac_sw_1_0.x1.x11.A single_10b_cdac_1.cdac_sw_1_0.x1.x9.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9421 VSREF single_10b_cdac_1.x8[7].x1.x7.A single_10b_cdac_1.x8[7].x1.x9.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9422 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9423 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9424 VDREF single_10b_cdac_1.x8[6].x1.x10.A single_10b_cdac_1.x8[6].x3.ckb VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9425 VDREF SWP_IN[8] a_40052_34754# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9426 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9427 a_16257_36566# single_10b_cdac_1.x6[5].x1.x8.A single_10b_cdac_1.x6[5].x1.x5.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9428 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9429 VSREF single_10b_cdac_1.x3[1].x1.x4.A single_10b_cdac_1.x3[1].x1.x6.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9430 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9431 VDREF single_10b_cdac_1.cdac_sw_4_1.x1.x8.A single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9432 VSREF single_10b_cdac_0.x10[8].x2.swp single_10b_cdac_0.x10[8].x2.swn VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9433 single_10b_cdac_1.x6[5].x2.swp single_10b_cdac_1.x6[5].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9434 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9435 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x11.A single_10b_cdac_0.cdac_sw_8_0.x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9436 single_10b_cdac_0.cdac_sw_2_1.x2.swn single_10b_cdac_0.cdac_sw_2_1.x2.swp VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9437 single_10b_cdac_0.x6[4].x2.swn single_10b_cdac_0.x6[4].x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9438 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9439 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9440 single_10b_cdac_0.x6[4].x1.x10.A single_10b_cdac_0.x6[4].x1.x8.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9441 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9442 VSREF single_10b_cdac_0.x4[2].x1.x9.A a_59511_35702# VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9443 VCN single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9444 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9445 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9446 VDREF single_10b_cdac_1.cdac_sw_4_1.x3.ckb single_10b_cdac_1.cdac_sw_4_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9447 VDREF single_10b_cdac_0.x8[6].x1.x6.A single_10b_cdac_0.x8[6].x1.x8.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9448 single_10b_cdac_0.x3[1].x3.ck single_10b_cdac_0.x3[1].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9449 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9450 single_10b_cdac_1.cdac_sw_1_0.x3.ck single_10b_cdac_1.cdac_sw_1_0.x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9451 VDREF single_10b_cdac_0.x4[3].x1.x9.A single_10b_cdac_0.x4[3].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9452 VSREF single_10b_cdac_1.x4[2].x1.x10.A single_10b_cdac_1.x4[2].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9453 VSREF CF[8] single_10b_cdac_0.x10[8].x1.x3.Y VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9454 single_10b_cdac_1.cdac_sw_2_1.x3.ck single_10b_cdac_1.cdac_sw_2_1.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9455 VSREF single_10b_cdac_0.cdac_sw_8_0.x1.x10.A single_10b_cdac_0.cdac_sw_8_0.x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9456 single_10b_cdac_0.x10b_cap_array_0.SW[0] single_10b_cdac_0.cdac_sw_16_0.x3.ckb a_34490_25722# VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9457 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9458 VDREF single_10b_cdac_1.x10[8].x1.x9.A single_10b_cdac_1.x10[8].x1.x11.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9459 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9460 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9461 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9462 single_10b_cdac_0.cdac_sw_1_2.x3.ck single_10b_cdac_0.cdac_sw_1_2.x3.ckb VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9463 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9464 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9465 VCN single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9466 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9467 single_10b_cdac_1.cdac_sw_8_1.x1.x3.Y CF[2] VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9468 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9469 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9470 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9471 single_10b_cdac_0.x10[8].x1.x10.A single_10b_cdac_0.x10[8].x1.x8.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9472 VCN single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9473 VCP single_10b_cdac_0.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9474 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9475 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9476 VCP single_10b_cdac_1.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9477 VCP single_10b_cdac_0.x8[7].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9478 single_10b_cdac_0.x3[1].dac_out single_10b_cdac_0.x3[1].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9479 VCP single_10b_cdac_0.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9480 single_10b_cdac_1.cdac_sw_8_0.x1.x7.A single_10b_cdac_1.cdac_sw_8_0.x1.x5.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9481 VDREF single_10b_cdac_1.x6[5].x1.x11.A single_10b_cdac_1.x6[5].x2.swp VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9482 VSREF single_10b_cdac_1.cdac_sw_16_0.x1.x8.A single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9483 single_10b_cdac_1.x3[0].x2.swp single_10b_cdac_1.x3[0].x1.x11.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9484 single_10b_cdac_0.cdac_sw_16_0.x2.swn single_10b_cdac_0.cdac_sw_16_0.x2.swp VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9485 single_10b_cdac_0.x8[7].dac_out single_10b_cdac_0.x8[7].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9486 VSREF single_10b_cdac_0.x8[7].x1.x11.A single_10b_cdac_0.x8[7].x2.swp VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9487 VCN single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9488 single_10b_cdac_1.x4[3].x2.swp single_10b_cdac_1.x4[3].x1.x11.A VDREF VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9489 VCN single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9490 VCP single_10b_cdac_1.x10[8].dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9491 VDREF single_10b_cdac_1.x10[8].x1.x4.A single_10b_cdac_1.x10[8].x1.x6.A VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9492 a_47370_25722# SWN_IN[4] VDREF VDREF sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X9493 single_10b_cdac_0.x6[5].x3.ck single_10b_cdac_0.x6[5].x3.ckb VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9494 VSREF single_10b_cdac_1.cdac_sw_1_0.x3.ckb single_10b_cdac_1.cdac_sw_1_0.x3.ck VSREF sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9495 VDREF CF[7] single_10b_cdac_0.x8[7].x1.x3.Y VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9496 VCP single_10b_cdac_1.cdac_sw_1_2.dac_out sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9497 VCN single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9498 VSREF single_10b_cdac_1.x2[0].x1.x10.A single_10b_cdac_1.x2[0].x3.ckb VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9499 single_10b_cdac_1.x6[4].dac_out single_10b_cdac_1.x6[4].x2.swn VCM VSREF sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9500 VDREF single_10b_cdac_1.cdac_sw_2_1.x3.ckb single_10b_cdac_1.cdac_sw_2_1.x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9501 single_10b_cdac_0.cdac_sw_8_0.x3.ckb single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VSREF VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9502 VSREF single_10b_cdac_0.x8[6].x1.x9.A single_10b_cdac_0.x8[6].x1.x11.A VSREF sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9503 VDREF single_10b_cdac_0.x3[1].x3.ckb single_10b_cdac_0.x3[1].x3.ck VDREF sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 VCN VSREF 0.797471p
C1 VCP VSREF 0.797471p
C2 SWN_IN[9] VSREF 35.5254f
C3 SWN_IN[8] VSREF 35.6574f
C4 SWP_IN[0] VSREF 86.4056f
C5 SWP_IN[1] VSREF 86.2736f
C6 SWN_IN[7] VSREF 39.0745f
C7 SWN_IN[6] VSREF 39.206497f
C8 SWN_IN[5] VSREF 45.9431f
C9 SWN_IN[4] VSREF 46.075104f
C10 SWN_IN[3] VSREF 57.810303f
C11 SWN_IN[2] VSREF 57.9423f
C12 SWP_IN[2] VSREF 57.9423f
C13 SWP_IN[3] VSREF 57.810303f
C14 SWP_IN[4] VSREF 46.075104f
C15 SWP_IN[5] VSREF 45.9431f
C16 SWP_IN[6] VSREF 39.206497f
C17 SWP_IN[7] VSREF 39.0745f
C18 SWN_IN[1] VSREF 86.2736f
C19 SWN_IN[0] VSREF 86.4056f
C20 SWP_IN[8] VSREF 35.6574f
C21 SWP_IN[9] VSREF 35.5254f
C22 VCM VSREF 0.473688p
C23 CF[0] VSREF 58.749306f
C24 CF[1] VSREF 58.749306f
C25 CF[2] VSREF 48.166103f
C26 CF[3] VSREF 48.166103f
C27 CF[4] VSREF 48.1086f
C28 CF[5] VSREF 48.1086f
C29 CF[6] VSREF 48.0511f
C30 CF[7] VSREF 48.0511f
C31 CF[8] VSREF 48.022396f
C32 CF[9] VSREF 48.022396f
C33 VDREF VSREF 1.71727p
C34 m1_49372_13869# VSREF 0.091357f $ **FLOATING
C35 m1_15778_13869# VSREF 0.091357f $ **FLOATING
C36 m1_51112_46803# VSREF 0.091357f $ **FLOATING
C37 m1_17518_46803# VSREF 0.091357f $ **FLOATING
C38 single_10b_cdac_0.cdac_sw_1_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C39 single_10b_cdac_0.cdac_sw_1_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C40 single_10b_cdac_0.cdac_sw_1_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C41 single_10b_cdac_0.cdac_sw_1_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C42 single_10b_cdac_0.cdac_sw_1_1.x1.x11.A VSREF 2.51762f $ **FLOATING
C43 single_10b_cdac_0.cdac_sw_1_1.x1.x7.A VSREF 0.615623f $ **FLOATING
C44 single_10b_cdac_0.cdac_sw_1_1.x1.x5.A VSREF 0.736451f $ **FLOATING
C45 single_10b_cdac_0.cdac_sw_1_1.x1.x3.Y VSREF 0.60393f $ **FLOATING
C46 single_10b_cdac_0.cdac_sw_2_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C47 single_10b_cdac_0.cdac_sw_2_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C48 single_10b_cdac_0.cdac_sw_2_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C49 single_10b_cdac_0.cdac_sw_2_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C50 single_10b_cdac_0.cdac_sw_2_1.x1.x11.A VSREF 2.51762f $ **FLOATING
C51 single_10b_cdac_0.cdac_sw_2_1.x1.x7.A VSREF 0.615623f $ **FLOATING
C52 single_10b_cdac_0.cdac_sw_2_1.x1.x5.A VSREF 0.736451f $ **FLOATING
C53 single_10b_cdac_0.cdac_sw_2_1.x1.x3.Y VSREF 0.60393f $ **FLOATING
C54 single_10b_cdac_0.cdac_sw_4_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C55 single_10b_cdac_0.cdac_sw_4_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C56 single_10b_cdac_0.cdac_sw_4_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C57 single_10b_cdac_0.cdac_sw_4_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C58 single_10b_cdac_0.cdac_sw_4_1.x1.x11.A VSREF 2.51762f $ **FLOATING
C59 single_10b_cdac_0.cdac_sw_4_1.x1.x7.A VSREF 0.615623f $ **FLOATING
C60 single_10b_cdac_0.cdac_sw_4_1.x1.x5.A VSREF 0.736451f $ **FLOATING
C61 single_10b_cdac_0.cdac_sw_4_1.x1.x3.Y VSREF 0.60393f $ **FLOATING
C62 single_10b_cdac_0.cdac_sw_8_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C63 single_10b_cdac_0.cdac_sw_8_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C64 single_10b_cdac_0.cdac_sw_8_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C65 single_10b_cdac_0.cdac_sw_8_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C66 single_10b_cdac_0.cdac_sw_8_1.x1.x11.A VSREF 2.51762f $ **FLOATING
C67 single_10b_cdac_0.cdac_sw_8_1.x1.x7.A VSREF 0.615623f $ **FLOATING
C68 single_10b_cdac_0.cdac_sw_8_1.x1.x5.A VSREF 0.736451f $ **FLOATING
C69 single_10b_cdac_0.cdac_sw_8_1.x1.x3.Y VSREF 0.60393f $ **FLOATING
C70 single_10b_cdac_0.x2[0].x1.x11.A VSREF 2.51762f $ **FLOATING
C71 single_10b_cdac_0.x2[0].x1.x7.A VSREF 0.615623f $ **FLOATING
C72 single_10b_cdac_0.x2[0].x1.x5.A VSREF 0.736451f $ **FLOATING
C73 single_10b_cdac_0.x2[0].x1.x3.Y VSREF 0.60393f $ **FLOATING
C74 single_10b_cdac_0.cdac_sw_16_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C75 single_10b_cdac_0.cdac_sw_16_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C76 single_10b_cdac_0.cdac_sw_16_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C77 single_10b_cdac_0.cdac_sw_16_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C78 single_10b_cdac_1.cdac_sw_1_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C79 single_10b_cdac_1.cdac_sw_1_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C80 single_10b_cdac_1.cdac_sw_1_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C81 single_10b_cdac_1.cdac_sw_1_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C82 single_10b_cdac_1.cdac_sw_1_1.x1.x11.A VSREF 2.51762f $ **FLOATING
C83 single_10b_cdac_1.cdac_sw_1_1.x1.x7.A VSREF 0.615623f $ **FLOATING
C84 single_10b_cdac_1.cdac_sw_1_1.x1.x5.A VSREF 0.736451f $ **FLOATING
C85 single_10b_cdac_1.cdac_sw_1_1.x1.x3.Y VSREF 0.60393f $ **FLOATING
C86 single_10b_cdac_1.cdac_sw_2_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C87 single_10b_cdac_1.cdac_sw_2_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C88 single_10b_cdac_1.cdac_sw_2_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C89 single_10b_cdac_1.cdac_sw_2_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C90 single_10b_cdac_1.cdac_sw_2_1.x1.x11.A VSREF 2.51762f $ **FLOATING
C91 single_10b_cdac_1.cdac_sw_2_1.x1.x7.A VSREF 0.615623f $ **FLOATING
C92 single_10b_cdac_1.cdac_sw_2_1.x1.x5.A VSREF 0.736451f $ **FLOATING
C93 single_10b_cdac_1.cdac_sw_2_1.x1.x3.Y VSREF 0.60393f $ **FLOATING
C94 single_10b_cdac_1.cdac_sw_4_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C95 single_10b_cdac_1.cdac_sw_4_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C96 single_10b_cdac_1.cdac_sw_4_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C97 single_10b_cdac_1.cdac_sw_4_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C98 single_10b_cdac_1.cdac_sw_4_1.x1.x11.A VSREF 2.51762f $ **FLOATING
C99 single_10b_cdac_1.cdac_sw_4_1.x1.x7.A VSREF 0.615623f $ **FLOATING
C100 single_10b_cdac_1.cdac_sw_4_1.x1.x5.A VSREF 0.736451f $ **FLOATING
C101 single_10b_cdac_1.cdac_sw_4_1.x1.x3.Y VSREF 0.60393f $ **FLOATING
C102 single_10b_cdac_1.cdac_sw_8_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C103 single_10b_cdac_1.cdac_sw_8_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C104 single_10b_cdac_1.cdac_sw_8_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C105 single_10b_cdac_1.cdac_sw_8_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C106 single_10b_cdac_1.cdac_sw_8_1.x1.x11.A VSREF 2.51762f $ **FLOATING
C107 single_10b_cdac_1.cdac_sw_8_1.x1.x7.A VSREF 0.615623f $ **FLOATING
C108 single_10b_cdac_1.cdac_sw_8_1.x1.x5.A VSREF 0.736451f $ **FLOATING
C109 single_10b_cdac_1.cdac_sw_8_1.x1.x3.Y VSREF 0.60393f $ **FLOATING
C110 single_10b_cdac_1.x2[0].x1.x11.A VSREF 2.51762f $ **FLOATING
C111 single_10b_cdac_1.x2[0].x1.x7.A VSREF 0.615623f $ **FLOATING
C112 single_10b_cdac_1.x2[0].x1.x5.A VSREF 0.736451f $ **FLOATING
C113 single_10b_cdac_1.x2[0].x1.x3.Y VSREF 0.60393f $ **FLOATING
C114 single_10b_cdac_1.cdac_sw_16_0.x1.x11.A VSREF 2.51762f $ **FLOATING
C115 single_10b_cdac_1.cdac_sw_16_0.x1.x7.A VSREF 0.615623f $ **FLOATING
C116 single_10b_cdac_1.cdac_sw_16_0.x1.x5.A VSREF 0.736451f $ **FLOATING
C117 single_10b_cdac_1.cdac_sw_16_0.x1.x3.Y VSREF 0.60393f $ **FLOATING
C118 single_10b_cdac_0.cdac_sw_1_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C119 single_10b_cdac_0.cdac_sw_1_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C120 single_10b_cdac_0.cdac_sw_1_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C121 single_10b_cdac_0.cdac_sw_1_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C122 single_10b_cdac_0.cdac_sw_1_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C123 single_10b_cdac_0.cdac_sw_1_1.x1.x10.A VSREF 2.51762f $ **FLOATING
C124 single_10b_cdac_0.cdac_sw_1_1.x1.x8.A VSREF 2.14748f $ **FLOATING
C125 single_10b_cdac_0.cdac_sw_1_1.x1.x6.A VSREF 0.615623f $ **FLOATING
C126 single_10b_cdac_0.cdac_sw_1_1.x1.x4.A VSREF 0.736451f $ **FLOATING
C127 single_10b_cdac_0.cdac_sw_1_1.x1.x9.A VSREF 2.26866f $ **FLOATING
C128 single_10b_cdac_0.cdac_sw_2_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C129 single_10b_cdac_0.cdac_sw_2_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C130 single_10b_cdac_0.cdac_sw_2_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C131 single_10b_cdac_0.cdac_sw_2_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C132 single_10b_cdac_0.cdac_sw_2_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C133 single_10b_cdac_0.cdac_sw_2_1.x1.x10.A VSREF 2.51762f $ **FLOATING
C134 single_10b_cdac_0.cdac_sw_2_1.x1.x8.A VSREF 2.14748f $ **FLOATING
C135 single_10b_cdac_0.cdac_sw_2_1.x1.x6.A VSREF 0.615623f $ **FLOATING
C136 single_10b_cdac_0.cdac_sw_2_1.x1.x4.A VSREF 0.736451f $ **FLOATING
C137 single_10b_cdac_0.cdac_sw_2_1.x1.x9.A VSREF 2.26866f $ **FLOATING
C138 single_10b_cdac_0.cdac_sw_4_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C139 single_10b_cdac_0.cdac_sw_4_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C140 single_10b_cdac_0.cdac_sw_4_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C141 single_10b_cdac_0.cdac_sw_4_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C142 single_10b_cdac_0.cdac_sw_4_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C143 single_10b_cdac_0.cdac_sw_4_1.x1.x10.A VSREF 2.51762f $ **FLOATING
C144 single_10b_cdac_0.cdac_sw_4_1.x1.x8.A VSREF 2.14748f $ **FLOATING
C145 single_10b_cdac_0.cdac_sw_4_1.x1.x6.A VSREF 0.615623f $ **FLOATING
C146 single_10b_cdac_0.cdac_sw_4_1.x1.x4.A VSREF 0.736451f $ **FLOATING
C147 single_10b_cdac_0.cdac_sw_4_1.x1.x9.A VSREF 2.26866f $ **FLOATING
C148 single_10b_cdac_0.cdac_sw_8_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C149 single_10b_cdac_0.cdac_sw_8_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C150 single_10b_cdac_0.cdac_sw_8_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C151 single_10b_cdac_0.cdac_sw_8_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C152 single_10b_cdac_0.cdac_sw_8_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C153 single_10b_cdac_0.cdac_sw_8_1.x1.x10.A VSREF 2.51762f $ **FLOATING
C154 single_10b_cdac_0.cdac_sw_8_1.x1.x8.A VSREF 2.14748f $ **FLOATING
C155 single_10b_cdac_0.cdac_sw_8_1.x1.x6.A VSREF 0.615623f $ **FLOATING
C156 single_10b_cdac_0.cdac_sw_8_1.x1.x4.A VSREF 0.736451f $ **FLOATING
C157 single_10b_cdac_0.cdac_sw_8_1.x1.x9.A VSREF 2.26866f $ **FLOATING
C158 single_10b_cdac_0.x2[0].x1.x10.A VSREF 2.51762f $ **FLOATING
C159 single_10b_cdac_0.x2[0].x1.x8.A VSREF 2.14748f $ **FLOATING
C160 single_10b_cdac_0.x2[0].x1.x6.A VSREF 0.615623f $ **FLOATING
C161 single_10b_cdac_0.x2[0].x1.x4.A VSREF 0.736451f $ **FLOATING
C162 single_10b_cdac_0.x2[0].x1.x9.A VSREF 2.26866f $ **FLOATING
C163 single_10b_cdac_0.cdac_sw_16_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C164 single_10b_cdac_0.cdac_sw_16_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C165 single_10b_cdac_0.cdac_sw_16_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C166 single_10b_cdac_0.cdac_sw_16_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C167 single_10b_cdac_0.cdac_sw_16_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C168 single_10b_cdac_1.cdac_sw_1_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C169 single_10b_cdac_1.cdac_sw_1_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C170 single_10b_cdac_1.cdac_sw_1_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C171 single_10b_cdac_1.cdac_sw_1_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C172 single_10b_cdac_1.cdac_sw_1_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C173 single_10b_cdac_1.cdac_sw_1_1.x1.x10.A VSREF 2.51762f $ **FLOATING
C174 single_10b_cdac_1.cdac_sw_1_1.x1.x8.A VSREF 2.14748f $ **FLOATING
C175 single_10b_cdac_1.cdac_sw_1_1.x1.x6.A VSREF 0.615623f $ **FLOATING
C176 single_10b_cdac_1.cdac_sw_1_1.x1.x4.A VSREF 0.736451f $ **FLOATING
C177 single_10b_cdac_1.cdac_sw_1_1.x1.x9.A VSREF 2.26866f $ **FLOATING
C178 single_10b_cdac_1.cdac_sw_2_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C179 single_10b_cdac_1.cdac_sw_2_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C180 single_10b_cdac_1.cdac_sw_2_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C181 single_10b_cdac_1.cdac_sw_2_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C182 single_10b_cdac_1.cdac_sw_2_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C183 single_10b_cdac_1.cdac_sw_2_1.x1.x10.A VSREF 2.51762f $ **FLOATING
C184 single_10b_cdac_1.cdac_sw_2_1.x1.x8.A VSREF 2.14748f $ **FLOATING
C185 single_10b_cdac_1.cdac_sw_2_1.x1.x6.A VSREF 0.615623f $ **FLOATING
C186 single_10b_cdac_1.cdac_sw_2_1.x1.x4.A VSREF 0.736451f $ **FLOATING
C187 single_10b_cdac_1.cdac_sw_2_1.x1.x9.A VSREF 2.26866f $ **FLOATING
C188 single_10b_cdac_1.cdac_sw_4_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C189 single_10b_cdac_1.cdac_sw_4_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C190 single_10b_cdac_1.cdac_sw_4_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C191 single_10b_cdac_1.cdac_sw_4_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C192 single_10b_cdac_1.cdac_sw_4_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C193 single_10b_cdac_1.cdac_sw_4_1.x1.x10.A VSREF 2.51762f $ **FLOATING
C194 single_10b_cdac_1.cdac_sw_4_1.x1.x8.A VSREF 2.14748f $ **FLOATING
C195 single_10b_cdac_1.cdac_sw_4_1.x1.x6.A VSREF 0.615623f $ **FLOATING
C196 single_10b_cdac_1.cdac_sw_4_1.x1.x4.A VSREF 0.736451f $ **FLOATING
C197 single_10b_cdac_1.cdac_sw_4_1.x1.x9.A VSREF 2.26866f $ **FLOATING
C198 single_10b_cdac_1.cdac_sw_8_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C199 single_10b_cdac_1.cdac_sw_8_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C200 single_10b_cdac_1.cdac_sw_8_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C201 single_10b_cdac_1.cdac_sw_8_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C202 single_10b_cdac_1.cdac_sw_8_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C203 single_10b_cdac_1.cdac_sw_8_1.x1.x10.A VSREF 2.51762f $ **FLOATING
C204 single_10b_cdac_1.cdac_sw_8_1.x1.x8.A VSREF 2.14748f $ **FLOATING
C205 single_10b_cdac_1.cdac_sw_8_1.x1.x6.A VSREF 0.615623f $ **FLOATING
C206 single_10b_cdac_1.cdac_sw_8_1.x1.x4.A VSREF 0.736451f $ **FLOATING
C207 single_10b_cdac_1.cdac_sw_8_1.x1.x9.A VSREF 2.26866f $ **FLOATING
C208 single_10b_cdac_1.x2[0].x1.x10.A VSREF 2.51762f $ **FLOATING
C209 single_10b_cdac_1.x2[0].x1.x8.A VSREF 2.14748f $ **FLOATING
C210 single_10b_cdac_1.x2[0].x1.x6.A VSREF 0.615623f $ **FLOATING
C211 single_10b_cdac_1.x2[0].x1.x4.A VSREF 0.736451f $ **FLOATING
C212 single_10b_cdac_1.x2[0].x1.x9.A VSREF 2.26866f $ **FLOATING
C213 single_10b_cdac_1.cdac_sw_16_0.x1.x10.A VSREF 2.51762f $ **FLOATING
C214 single_10b_cdac_1.cdac_sw_16_0.x1.x8.A VSREF 2.14748f $ **FLOATING
C215 single_10b_cdac_1.cdac_sw_16_0.x1.x6.A VSREF 0.615623f $ **FLOATING
C216 single_10b_cdac_1.cdac_sw_16_0.x1.x4.A VSREF 0.736451f $ **FLOATING
C217 single_10b_cdac_1.cdac_sw_16_0.x1.x9.A VSREF 2.26866f $ **FLOATING
C218 single_10b_cdac_0.cdac_sw_1_0.x2.swn VSREF 2.78825f $ **FLOATING
C219 single_10b_cdac_0.cdac_sw_1_0.x2.swp VSREF 4.63322f $ **FLOATING
C220 a_64348_25713# VSREF 0.295532f $ **FLOATING
C221 single_10b_cdac_0.cdac_sw_1_0.x3.ck VSREF 3.14422f $ **FLOATING
C222 single_10b_cdac_0.x10b_cap_array_0.SW[9] VSREF 0.499508p $ **FLOATING
C223 single_10b_cdac_0.cdac_sw_1_0.x3.ckb VSREF 5.12291f $ **FLOATING
C224 a_63470_25722# VSREF 0.588398f $ **FLOATING
C225 single_10b_cdac_0.cdac_sw_1_1.x2.swn VSREF 2.78825f $ **FLOATING
C226 single_10b_cdac_0.cdac_sw_1_1.x2.swp VSREF 4.63322f $ **FLOATING
C227 a_61128_25713# VSREF 0.295532f $ **FLOATING
C228 single_10b_cdac_0.cdac_sw_1_1.x3.ck VSREF 3.14422f $ **FLOATING
C229 single_10b_cdac_0.x10b_cap_array_0.SW[8] VSREF 0.259038p $ **FLOATING
C230 single_10b_cdac_0.cdac_sw_1_1.x3.ckb VSREF 5.12291f $ **FLOATING
C231 a_60250_25722# VSREF 0.588398f $ **FLOATING
C232 single_10b_cdac_0.cdac_sw_2_0.x2.swn VSREF 3.409f $ **FLOATING
C233 a_65812_26714# VSREF 16.1733f $ **FLOATING
C234 a_64934_30193# VSREF 8.6969f $ **FLOATING
C235 single_10b_cdac_0.x3[0].dac_out VSREF 52.5439f $ **FLOATING
C236 a_62592_26714# VSREF 16.1733f $ **FLOATING
C237 a_61714_30193# VSREF 8.6969f $ **FLOATING
C238 single_10b_cdac_0.cdac_sw_2_0.x2.swp VSREF 5.35635f $ **FLOATING
C239 a_57908_25713# VSREF 0.940559f $ **FLOATING
C240 single_10b_cdac_0.cdac_sw_2_0.x3.ck VSREF 3.76497f $ **FLOATING
C241 single_10b_cdac_0.x10b_cap_array_0.SW[7] VSREF 0.140663p $ **FLOATING
C242 single_10b_cdac_0.cdac_sw_2_0.x3.ckb VSREF 5.84648f $ **FLOATING
C243 a_57030_25722# VSREF 1.90105f $ **FLOATING
C244 single_10b_cdac_0.cdac_sw_2_1.x2.swn VSREF 3.409f $ **FLOATING
C245 single_10b_cdac_0.cdac_sw_2_1.x2.swp VSREF 5.35635f $ **FLOATING
C246 a_54688_25713# VSREF 0.940559f $ **FLOATING
C247 single_10b_cdac_0.cdac_sw_2_1.x3.ck VSREF 3.76497f $ **FLOATING
C248 single_10b_cdac_0.x10b_cap_array_0.SW[6] VSREF 80.502f $ **FLOATING
C249 single_10b_cdac_0.cdac_sw_2_1.x3.ckb VSREF 5.84648f $ **FLOATING
C250 a_53810_25722# VSREF 1.90105f $ **FLOATING
C251 single_10b_cdac_0.cdac_sw_4_0.x2.swn VSREF 4.65051f $ **FLOATING
C252 single_10b_cdac_0.cdac_sw_4_0.x2.swp VSREF 6.80262f $ **FLOATING
C253 a_51468_25713# VSREF 2.0817f $ **FLOATING
C254 single_10b_cdac_0.cdac_sw_4_0.x3.ck VSREF 5.00691f $ **FLOATING
C255 single_10b_cdac_0.x10b_cap_array_0.SW[5] VSREF 58.667103f $ **FLOATING
C256 single_10b_cdac_0.cdac_sw_4_0.x3.ckb VSREF 7.29232f $ **FLOATING
C257 a_50590_25722# VSREF 3.93995f $ **FLOATING
C258 single_10b_cdac_0.cdac_sw_4_1.x2.swn VSREF 4.65051f $ **FLOATING
C259 single_10b_cdac_0.cdac_sw_4_1.x2.swp VSREF 6.80262f $ **FLOATING
C260 a_48248_25713# VSREF 2.0817f $ **FLOATING
C261 single_10b_cdac_0.cdac_sw_4_1.x3.ck VSREF 5.00691f $ **FLOATING
C262 single_10b_cdac_0.x10b_cap_array_0.SW[4] VSREF 45.7835f $ **FLOATING
C263 single_10b_cdac_0.cdac_sw_4_1.x3.ckb VSREF 7.29232f $ **FLOATING
C264 a_47370_25722# VSREF 3.93995f $ **FLOATING
C265 single_10b_cdac_0.cdac_sw_8_0.x2.swn VSREF 7.13352f $ **FLOATING
C266 single_10b_cdac_0.cdac_sw_8_0.x2.swp VSREF 9.69516f $ **FLOATING
C267 a_45028_25713# VSREF 4.28676f $ **FLOATING
C268 single_10b_cdac_0.cdac_sw_8_0.x3.ck VSREF 7.49036f $ **FLOATING
C269 single_10b_cdac_0.x10b_cap_array_0.SW[3] VSREF 44.920498f $ **FLOATING
C270 single_10b_cdac_0.cdac_sw_8_0.x3.ckb VSREF 10.1849f $ **FLOATING
C271 a_44150_25722# VSREF 8.01774f $ **FLOATING
C272 single_10b_cdac_0.cdac_sw_8_1.x2.swn VSREF 7.13352f $ **FLOATING
C273 single_10b_cdac_0.cdac_sw_8_1.x2.swp VSREF 9.69516f $ **FLOATING
C274 a_41808_25713# VSREF 4.28676f $ **FLOATING
C275 single_10b_cdac_0.cdac_sw_8_1.x3.ck VSREF 7.49036f $ **FLOATING
C276 single_10b_cdac_0.x10b_cap_array_0.SW[2] VSREF 40.3181f $ **FLOATING
C277 single_10b_cdac_0.cdac_sw_8_1.x3.ckb VSREF 10.1849f $ **FLOATING
C278 a_40930_25722# VSREF 8.01774f $ **FLOATING
C279 single_10b_cdac_0.x3[1].dac_out VSREF 54.380604f $ **FLOATING
C280 single_10b_cdac_0.x2[0].x2.swn VSREF 12.0995f $ **FLOATING
C281 a_59372_31002# VSREF 8.01774f $ **FLOATING
C282 a_58494_32737# VSREF 4.28676f $ **FLOATING
C283 single_10b_cdac_0.x4[2].dac_out VSREF 40.3181f $ **FLOATING
C284 a_56152_31002# VSREF 8.01774f $ **FLOATING
C285 a_55274_32737# VSREF 4.28676f $ **FLOATING
C286 single_10b_cdac_0.x4[3].dac_out VSREF 44.920498f $ **FLOATING
C287 a_52932_33146# VSREF 3.93995f $ **FLOATING
C288 a_52054_34009# VSREF 2.0817f $ **FLOATING
C289 single_10b_cdac_0.x6[4].dac_out VSREF 45.7835f $ **FLOATING
C290 a_49712_33146# VSREF 3.93995f $ **FLOATING
C291 a_48834_34009# VSREF 2.0817f $ **FLOATING
C292 single_10b_cdac_0.x6[5].dac_out VSREF 58.667103f $ **FLOATING
C293 a_46492_34218# VSREF 1.90105f $ **FLOATING
C294 a_45614_34645# VSREF 0.940559f $ **FLOATING
C295 single_10b_cdac_0.x8[6].dac_out VSREF 80.502f $ **FLOATING
C296 a_43272_34218# VSREF 1.90105f $ **FLOATING
C297 a_42394_34645# VSREF 0.940559f $ **FLOATING
C298 single_10b_cdac_0.x2[0].x2.swp VSREF 15.4802f $ **FLOATING
C299 a_38588_25713# VSREF 8.6969f $ **FLOATING
C300 single_10b_cdac_0.x2[0].x3.ck VSREF 12.4572f $ **FLOATING
C301 single_10b_cdac_0.x10b_cap_array_0.SW[1] VSREF 54.380604f $ **FLOATING
C302 single_10b_cdac_0.x2[0].x3.ckb VSREF 15.9699f $ **FLOATING
C303 a_37710_25722# VSREF 16.1733f $ **FLOATING
C304 single_10b_cdac_0.cdac_sw_16_0.x2.swn VSREF 12.0995f $ **FLOATING
C305 single_10b_cdac_0.cdac_sw_16_0.x2.swp VSREF 15.4802f $ **FLOATING
C306 a_35368_25713# VSREF 8.6969f $ **FLOATING
C307 single_10b_cdac_0.cdac_sw_16_0.x3.ck VSREF 12.4572f $ **FLOATING
C308 single_10b_cdac_0.x10b_cap_array_0.SW[0] VSREF 52.5439f $ **FLOATING
C309 single_10b_cdac_0.cdac_sw_16_0.x3.ckb VSREF 15.9699f $ **FLOATING
C310 a_34490_25722# VSREF 16.1733f $ **FLOATING
C311 single_10b_cdac_1.cdac_sw_1_0.x2.swn VSREF 2.78825f $ **FLOATING
C312 single_10b_cdac_1.cdac_sw_1_0.x2.swp VSREF 4.63322f $ **FLOATING
C313 a_30754_25713# VSREF 0.295532f $ **FLOATING
C314 single_10b_cdac_1.cdac_sw_1_0.x3.ck VSREF 3.14422f $ **FLOATING
C315 single_10b_cdac_1.x10b_cap_array_0.SW[9] VSREF 0.499508p $ **FLOATING
C316 single_10b_cdac_1.cdac_sw_1_0.x3.ckb VSREF 5.12291f $ **FLOATING
C317 a_29876_25722# VSREF 0.588398f $ **FLOATING
C318 single_10b_cdac_1.cdac_sw_1_1.x2.swn VSREF 2.78825f $ **FLOATING
C319 single_10b_cdac_1.cdac_sw_1_1.x2.swp VSREF 4.63322f $ **FLOATING
C320 a_27534_25713# VSREF 0.295532f $ **FLOATING
C321 single_10b_cdac_1.cdac_sw_1_1.x3.ck VSREF 3.14422f $ **FLOATING
C322 single_10b_cdac_1.x10b_cap_array_0.SW[8] VSREF 0.259038p $ **FLOATING
C323 single_10b_cdac_1.cdac_sw_1_1.x3.ckb VSREF 5.12291f $ **FLOATING
C324 a_26656_25722# VSREF 0.588398f $ **FLOATING
C325 single_10b_cdac_1.cdac_sw_2_0.x2.swn VSREF 3.409f $ **FLOATING
C326 single_10b_cdac_0.x8[7].dac_out VSREF 0.140663p $ **FLOATING
C327 a_40052_34754# VSREF 0.588398f $ **FLOATING
C328 a_39174_34963# VSREF 0.295532f $ **FLOATING
C329 single_10b_cdac_0.x10[8].dac_out VSREF 0.259038p $ **FLOATING
C330 a_36832_34754# VSREF 0.588398f $ **FLOATING
C331 a_35954_34963# VSREF 0.295532f $ **FLOATING
C332 single_10b_cdac_0.cdac_sw_1_2.dac_out VSREF 0.499508p $ **FLOATING
C333 a_32218_26714# VSREF 16.1733f $ **FLOATING
C334 a_31340_30193# VSREF 8.6969f $ **FLOATING
C335 single_10b_cdac_1.x3[0].dac_out VSREF 52.5439f $ **FLOATING
C336 a_28998_26714# VSREF 16.1733f $ **FLOATING
C337 a_28120_30193# VSREF 8.6969f $ **FLOATING
C338 single_10b_cdac_1.cdac_sw_2_0.x2.swp VSREF 5.35635f $ **FLOATING
C339 a_24314_25713# VSREF 0.940559f $ **FLOATING
C340 single_10b_cdac_1.cdac_sw_2_0.x3.ck VSREF 3.76497f $ **FLOATING
C341 single_10b_cdac_1.x10b_cap_array_0.SW[7] VSREF 0.140663p $ **FLOATING
C342 single_10b_cdac_1.cdac_sw_2_0.x3.ckb VSREF 5.84648f $ **FLOATING
C343 a_23436_25722# VSREF 1.90105f $ **FLOATING
C344 single_10b_cdac_1.cdac_sw_2_1.x2.swn VSREF 3.409f $ **FLOATING
C345 single_10b_cdac_1.cdac_sw_2_1.x2.swp VSREF 5.35635f $ **FLOATING
C346 a_21094_25713# VSREF 0.940559f $ **FLOATING
C347 single_10b_cdac_1.cdac_sw_2_1.x3.ck VSREF 3.76497f $ **FLOATING
C348 single_10b_cdac_1.x10b_cap_array_0.SW[6] VSREF 80.502f $ **FLOATING
C349 single_10b_cdac_1.cdac_sw_2_1.x3.ckb VSREF 5.84648f $ **FLOATING
C350 a_20216_25722# VSREF 1.90105f $ **FLOATING
C351 single_10b_cdac_1.cdac_sw_4_0.x2.swn VSREF 4.65051f $ **FLOATING
C352 single_10b_cdac_1.cdac_sw_4_0.x2.swp VSREF 6.80262f $ **FLOATING
C353 a_17874_25713# VSREF 2.0817f $ **FLOATING
C354 single_10b_cdac_1.cdac_sw_4_0.x3.ck VSREF 5.00691f $ **FLOATING
C355 single_10b_cdac_1.x10b_cap_array_0.SW[5] VSREF 58.667103f $ **FLOATING
C356 single_10b_cdac_1.cdac_sw_4_0.x3.ckb VSREF 7.29232f $ **FLOATING
C357 a_16996_25722# VSREF 3.93995f $ **FLOATING
C358 single_10b_cdac_1.cdac_sw_4_1.x2.swn VSREF 4.65051f $ **FLOATING
C359 single_10b_cdac_1.cdac_sw_4_1.x2.swp VSREF 6.80262f $ **FLOATING
C360 a_14654_25713# VSREF 2.0817f $ **FLOATING
C361 single_10b_cdac_1.cdac_sw_4_1.x3.ck VSREF 5.00691f $ **FLOATING
C362 single_10b_cdac_1.x10b_cap_array_0.SW[4] VSREF 45.7835f $ **FLOATING
C363 single_10b_cdac_1.cdac_sw_4_1.x3.ckb VSREF 7.29232f $ **FLOATING
C364 a_13776_25722# VSREF 3.93995f $ **FLOATING
C365 single_10b_cdac_1.cdac_sw_8_0.x2.swn VSREF 7.13352f $ **FLOATING
C366 single_10b_cdac_1.cdac_sw_8_0.x2.swp VSREF 9.69516f $ **FLOATING
C367 a_11434_25713# VSREF 4.28676f $ **FLOATING
C368 single_10b_cdac_1.cdac_sw_8_0.x3.ck VSREF 7.49036f $ **FLOATING
C369 single_10b_cdac_1.x10b_cap_array_0.SW[3] VSREF 44.920498f $ **FLOATING
C370 single_10b_cdac_1.cdac_sw_8_0.x3.ckb VSREF 10.1849f $ **FLOATING
C371 a_10556_25722# VSREF 8.01774f $ **FLOATING
C372 single_10b_cdac_1.cdac_sw_8_1.x2.swn VSREF 7.13352f $ **FLOATING
C373 single_10b_cdac_1.cdac_sw_8_1.x2.swp VSREF 9.69516f $ **FLOATING
C374 a_8214_25713# VSREF 4.28676f $ **FLOATING
C375 single_10b_cdac_1.cdac_sw_8_1.x3.ck VSREF 7.49036f $ **FLOATING
C376 single_10b_cdac_1.x10b_cap_array_0.SW[2] VSREF 40.3181f $ **FLOATING
C377 single_10b_cdac_1.cdac_sw_8_1.x3.ckb VSREF 10.1849f $ **FLOATING
C378 a_7336_25722# VSREF 8.01774f $ **FLOATING
C379 single_10b_cdac_1.x3[1].dac_out VSREF 54.380604f $ **FLOATING
C380 single_10b_cdac_1.x2[0].x2.swn VSREF 12.0995f $ **FLOATING
C381 a_25778_31002# VSREF 8.01774f $ **FLOATING
C382 a_24900_32737# VSREF 4.28676f $ **FLOATING
C383 single_10b_cdac_1.x4[2].dac_out VSREF 40.3181f $ **FLOATING
C384 a_22558_31002# VSREF 8.01774f $ **FLOATING
C385 a_21680_32737# VSREF 4.28676f $ **FLOATING
C386 single_10b_cdac_1.x4[3].dac_out VSREF 44.920498f $ **FLOATING
C387 a_19338_33146# VSREF 3.93995f $ **FLOATING
C388 a_18460_34009# VSREF 2.0817f $ **FLOATING
C389 single_10b_cdac_1.x6[4].dac_out VSREF 45.7835f $ **FLOATING
C390 a_16118_33146# VSREF 3.93995f $ **FLOATING
C391 a_15240_34009# VSREF 2.0817f $ **FLOATING
C392 single_10b_cdac_1.x6[5].dac_out VSREF 58.667103f $ **FLOATING
C393 a_12898_34218# VSREF 1.90105f $ **FLOATING
C394 a_12020_34645# VSREF 0.940559f $ **FLOATING
C395 single_10b_cdac_1.x8[6].dac_out VSREF 80.502f $ **FLOATING
C396 a_9678_34218# VSREF 1.90105f $ **FLOATING
C397 a_8800_34645# VSREF 0.940559f $ **FLOATING
C398 single_10b_cdac_1.x2[0].x2.swp VSREF 15.4802f $ **FLOATING
C399 a_4994_25713# VSREF 8.6969f $ **FLOATING
C400 single_10b_cdac_1.x2[0].x3.ck VSREF 12.4572f $ **FLOATING
C401 single_10b_cdac_1.x10b_cap_array_0.SW[1] VSREF 54.380604f $ **FLOATING
C402 single_10b_cdac_1.x2[0].x3.ckb VSREF 15.9699f $ **FLOATING
C403 a_4116_25722# VSREF 16.1733f $ **FLOATING
C404 single_10b_cdac_1.cdac_sw_16_0.x2.swn VSREF 12.0995f $ **FLOATING
C405 single_10b_cdac_1.cdac_sw_16_0.x2.swp VSREF 15.4802f $ **FLOATING
C406 a_1774_25713# VSREF 8.6969f $ **FLOATING
C407 single_10b_cdac_1.cdac_sw_16_0.x3.ck VSREF 12.4572f $ **FLOATING
C408 single_10b_cdac_1.x10b_cap_array_0.SW[0] VSREF 52.5439f $ **FLOATING
C409 single_10b_cdac_1.cdac_sw_16_0.x3.ckb VSREF 15.9699f $ **FLOATING
C410 a_896_25722# VSREF 16.1733f $ **FLOATING
C411 single_10b_cdac_1.x8[7].dac_out VSREF 0.140663p $ **FLOATING
C412 a_6458_34754# VSREF 0.588398f $ **FLOATING
C413 a_5580_34963# VSREF 0.295532f $ **FLOATING
C414 single_10b_cdac_1.x10[8].dac_out VSREF 0.259038p $ **FLOATING
C415 a_3238_34754# VSREF 0.588398f $ **FLOATING
C416 a_2360_34963# VSREF 0.295532f $ **FLOATING
C417 single_10b_cdac_1.cdac_sw_1_2.dac_out VSREF 0.499508p $ **FLOATING
C418 single_10b_cdac_0.x3[0].x1.x4.A VSREF 0.736451f $ **FLOATING
C419 single_10b_cdac_0.x3[0].x3.ck VSREF 12.4572f $ **FLOATING
C420 single_10b_cdac_0.x3[0].x1.x6.A VSREF 0.615623f $ **FLOATING
C421 single_10b_cdac_0.x3[0].x1.x10.A VSREF 2.51762f $ **FLOATING
C422 single_10b_cdac_0.x3[0].x3.ckb VSREF 15.9699f $ **FLOATING
C423 single_10b_cdac_0.x3[1].x1.x4.A VSREF 0.736451f $ **FLOATING
C424 single_10b_cdac_0.x3[1].x3.ck VSREF 12.4572f $ **FLOATING
C425 single_10b_cdac_0.x3[1].x1.x6.A VSREF 0.615623f $ **FLOATING
C426 single_10b_cdac_0.x3[1].x1.x10.A VSREF 2.51762f $ **FLOATING
C427 single_10b_cdac_0.x3[1].x3.ckb VSREF 15.9699f $ **FLOATING
C428 single_10b_cdac_0.x4[2].x1.x4.A VSREF 0.736451f $ **FLOATING
C429 single_10b_cdac_0.x4[2].x3.ck VSREF 7.49036f $ **FLOATING
C430 single_10b_cdac_0.x4[2].x1.x6.A VSREF 0.615623f $ **FLOATING
C431 single_10b_cdac_0.x4[2].x1.x10.A VSREF 2.51762f $ **FLOATING
C432 single_10b_cdac_0.x4[2].x3.ckb VSREF 10.1849f $ **FLOATING
C433 single_10b_cdac_0.x4[3].x1.x4.A VSREF 0.736451f $ **FLOATING
C434 single_10b_cdac_0.x4[3].x3.ck VSREF 7.49036f $ **FLOATING
C435 single_10b_cdac_0.x4[3].x1.x6.A VSREF 0.615623f $ **FLOATING
C436 single_10b_cdac_0.x4[3].x1.x10.A VSREF 2.51762f $ **FLOATING
C437 single_10b_cdac_0.x4[3].x3.ckb VSREF 10.1849f $ **FLOATING
C438 single_10b_cdac_0.x6[4].x1.x4.A VSREF 0.736451f $ **FLOATING
C439 single_10b_cdac_0.x6[4].x3.ck VSREF 5.00691f $ **FLOATING
C440 single_10b_cdac_0.x6[4].x1.x6.A VSREF 0.615623f $ **FLOATING
C441 single_10b_cdac_0.x6[4].x1.x10.A VSREF 2.51762f $ **FLOATING
C442 single_10b_cdac_0.x6[4].x3.ckb VSREF 7.29232f $ **FLOATING
C443 single_10b_cdac_0.x6[5].x1.x4.A VSREF 0.736451f $ **FLOATING
C444 single_10b_cdac_0.x6[5].x3.ck VSREF 5.00691f $ **FLOATING
C445 single_10b_cdac_0.x6[5].x1.x6.A VSREF 0.615623f $ **FLOATING
C446 single_10b_cdac_0.x6[5].x1.x10.A VSREF 2.51762f $ **FLOATING
C447 single_10b_cdac_0.x6[5].x3.ckb VSREF 7.29232f $ **FLOATING
C448 single_10b_cdac_0.x8[6].x1.x4.A VSREF 0.736451f $ **FLOATING
C449 single_10b_cdac_0.x8[6].x3.ck VSREF 3.76497f $ **FLOATING
C450 single_10b_cdac_0.x8[6].x1.x6.A VSREF 0.615623f $ **FLOATING
C451 single_10b_cdac_0.x8[6].x1.x10.A VSREF 2.51762f $ **FLOATING
C452 single_10b_cdac_0.x8[6].x3.ckb VSREF 5.84648f $ **FLOATING
C453 single_10b_cdac_0.x8[7].x1.x4.A VSREF 0.736451f $ **FLOATING
C454 single_10b_cdac_0.x8[7].x3.ck VSREF 3.76497f $ **FLOATING
C455 single_10b_cdac_0.x8[7].x1.x6.A VSREF 0.615623f $ **FLOATING
C456 single_10b_cdac_0.x8[7].x1.x10.A VSREF 2.51762f $ **FLOATING
C457 single_10b_cdac_0.x8[7].x3.ckb VSREF 5.84648f $ **FLOATING
C458 single_10b_cdac_0.x10[8].x1.x4.A VSREF 0.736451f $ **FLOATING
C459 single_10b_cdac_0.x10[8].x3.ck VSREF 3.14422f $ **FLOATING
C460 single_10b_cdac_0.x10[8].x1.x6.A VSREF 0.615623f $ **FLOATING
C461 single_10b_cdac_0.x10[8].x1.x10.A VSREF 2.51762f $ **FLOATING
C462 single_10b_cdac_0.x10[8].x3.ckb VSREF 5.12291f $ **FLOATING
C463 single_10b_cdac_0.cdac_sw_1_2.x1.x4.A VSREF 0.736451f $ **FLOATING
C464 single_10b_cdac_0.cdac_sw_1_2.x3.ck VSREF 3.14422f $ **FLOATING
C465 single_10b_cdac_0.cdac_sw_1_2.x1.x6.A VSREF 0.615623f $ **FLOATING
C466 single_10b_cdac_0.cdac_sw_1_2.x1.x10.A VSREF 2.51762f $ **FLOATING
C467 single_10b_cdac_0.cdac_sw_1_2.x3.ckb VSREF 5.12291f $ **FLOATING
C468 single_10b_cdac_1.x3[0].x1.x4.A VSREF 0.736451f $ **FLOATING
C469 single_10b_cdac_1.x3[0].x3.ck VSREF 12.4572f $ **FLOATING
C470 single_10b_cdac_1.x3[0].x1.x6.A VSREF 0.615623f $ **FLOATING
C471 single_10b_cdac_1.x3[0].x1.x10.A VSREF 2.51762f $ **FLOATING
C472 single_10b_cdac_1.x3[0].x3.ckb VSREF 15.9699f $ **FLOATING
C473 single_10b_cdac_1.x3[1].x1.x4.A VSREF 0.736451f $ **FLOATING
C474 single_10b_cdac_1.x3[1].x3.ck VSREF 12.4572f $ **FLOATING
C475 single_10b_cdac_1.x3[1].x1.x6.A VSREF 0.615623f $ **FLOATING
C476 single_10b_cdac_1.x3[1].x1.x10.A VSREF 2.51762f $ **FLOATING
C477 single_10b_cdac_1.x3[1].x3.ckb VSREF 15.9699f $ **FLOATING
C478 single_10b_cdac_1.x4[2].x1.x4.A VSREF 0.736451f $ **FLOATING
C479 single_10b_cdac_1.x4[2].x3.ck VSREF 7.49036f $ **FLOATING
C480 single_10b_cdac_1.x4[2].x1.x6.A VSREF 0.615623f $ **FLOATING
C481 single_10b_cdac_1.x4[2].x1.x10.A VSREF 2.51762f $ **FLOATING
C482 single_10b_cdac_1.x4[2].x3.ckb VSREF 10.1849f $ **FLOATING
C483 single_10b_cdac_1.x4[3].x1.x4.A VSREF 0.736451f $ **FLOATING
C484 single_10b_cdac_1.x4[3].x3.ck VSREF 7.49036f $ **FLOATING
C485 single_10b_cdac_1.x4[3].x1.x6.A VSREF 0.615623f $ **FLOATING
C486 single_10b_cdac_1.x4[3].x1.x10.A VSREF 2.51762f $ **FLOATING
C487 single_10b_cdac_1.x4[3].x3.ckb VSREF 10.1849f $ **FLOATING
C488 single_10b_cdac_1.x6[4].x1.x4.A VSREF 0.736451f $ **FLOATING
C489 single_10b_cdac_1.x6[4].x3.ck VSREF 5.00691f $ **FLOATING
C490 single_10b_cdac_1.x6[4].x1.x6.A VSREF 0.615623f $ **FLOATING
C491 single_10b_cdac_1.x6[4].x1.x10.A VSREF 2.51762f $ **FLOATING
C492 single_10b_cdac_1.x6[4].x3.ckb VSREF 7.29232f $ **FLOATING
C493 single_10b_cdac_1.x6[5].x1.x4.A VSREF 0.736451f $ **FLOATING
C494 single_10b_cdac_1.x6[5].x3.ck VSREF 5.00691f $ **FLOATING
C495 single_10b_cdac_1.x6[5].x1.x6.A VSREF 0.615623f $ **FLOATING
C496 single_10b_cdac_1.x6[5].x1.x10.A VSREF 2.51762f $ **FLOATING
C497 single_10b_cdac_1.x6[5].x3.ckb VSREF 7.29232f $ **FLOATING
C498 single_10b_cdac_1.x8[6].x1.x4.A VSREF 0.736451f $ **FLOATING
C499 single_10b_cdac_1.x8[6].x3.ck VSREF 3.76497f $ **FLOATING
C500 single_10b_cdac_1.x8[6].x1.x6.A VSREF 0.615623f $ **FLOATING
C501 single_10b_cdac_1.x8[6].x1.x10.A VSREF 2.51762f $ **FLOATING
C502 single_10b_cdac_1.x8[6].x3.ckb VSREF 5.84648f $ **FLOATING
C503 single_10b_cdac_1.x8[7].x1.x4.A VSREF 0.736451f $ **FLOATING
C504 single_10b_cdac_1.x8[7].x3.ck VSREF 3.76497f $ **FLOATING
C505 single_10b_cdac_1.x8[7].x1.x6.A VSREF 0.615623f $ **FLOATING
C506 single_10b_cdac_1.x8[7].x1.x10.A VSREF 2.51762f $ **FLOATING
C507 single_10b_cdac_1.x8[7].x3.ckb VSREF 5.84648f $ **FLOATING
C508 single_10b_cdac_1.x10[8].x1.x4.A VSREF 0.736451f $ **FLOATING
C509 single_10b_cdac_1.x10[8].x3.ck VSREF 3.14422f $ **FLOATING
C510 single_10b_cdac_1.x10[8].x1.x6.A VSREF 0.615623f $ **FLOATING
C511 single_10b_cdac_1.x10[8].x1.x10.A VSREF 2.51762f $ **FLOATING
C512 single_10b_cdac_1.x10[8].x3.ckb VSREF 5.12291f $ **FLOATING
C513 single_10b_cdac_1.cdac_sw_1_2.x1.x4.A VSREF 0.736451f $ **FLOATING
C514 single_10b_cdac_1.cdac_sw_1_2.x3.ck VSREF 3.14422f $ **FLOATING
C515 single_10b_cdac_1.cdac_sw_1_2.x1.x6.A VSREF 0.615623f $ **FLOATING
C516 single_10b_cdac_1.cdac_sw_1_2.x1.x10.A VSREF 2.51762f $ **FLOATING
C517 single_10b_cdac_1.cdac_sw_1_2.x3.ckb VSREF 5.12291f $ **FLOATING
C518 single_10b_cdac_0.x3[0].x2.swn VSREF 12.0995f $ **FLOATING
C519 single_10b_cdac_0.x3[1].x2.swn VSREF 12.0995f $ **FLOATING
C520 single_10b_cdac_0.x4[2].x2.swn VSREF 7.13352f $ **FLOATING
C521 single_10b_cdac_0.x4[3].x2.swn VSREF 7.13352f $ **FLOATING
C522 single_10b_cdac_0.x6[4].x2.swn VSREF 4.65051f $ **FLOATING
C523 single_10b_cdac_0.x6[5].x2.swn VSREF 4.65051f $ **FLOATING
C524 single_10b_cdac_0.x8[6].x2.swn VSREF 3.409f $ **FLOATING
C525 single_10b_cdac_0.x8[7].x2.swn VSREF 3.409f $ **FLOATING
C526 single_10b_cdac_0.x10[8].x2.swn VSREF 2.78825f $ **FLOATING
C527 single_10b_cdac_0.cdac_sw_1_2.x2.swn VSREF 2.78825f $ **FLOATING
C528 single_10b_cdac_1.x3[0].x2.swn VSREF 12.0995f $ **FLOATING
C529 single_10b_cdac_1.x3[1].x2.swn VSREF 12.0995f $ **FLOATING
C530 single_10b_cdac_1.x4[2].x2.swn VSREF 7.13352f $ **FLOATING
C531 single_10b_cdac_1.x4[3].x2.swn VSREF 7.13352f $ **FLOATING
C532 single_10b_cdac_1.x6[4].x2.swn VSREF 4.65051f $ **FLOATING
C533 single_10b_cdac_1.x6[5].x2.swn VSREF 4.65051f $ **FLOATING
C534 single_10b_cdac_1.x8[6].x2.swn VSREF 3.409f $ **FLOATING
C535 single_10b_cdac_1.x8[7].x2.swn VSREF 3.409f $ **FLOATING
C536 single_10b_cdac_1.x10[8].x2.swn VSREF 2.78825f $ **FLOATING
C537 single_10b_cdac_1.cdac_sw_1_2.x2.swn VSREF 2.78825f $ **FLOATING
C538 single_10b_cdac_0.x3[0].x1.x3.Y VSREF 0.60393f $ **FLOATING
C539 single_10b_cdac_0.x3[0].x1.x8.A VSREF 2.14748f $ **FLOATING
C540 single_10b_cdac_0.x3[0].x1.x5.A VSREF 0.736451f $ **FLOATING
C541 single_10b_cdac_0.x3[0].x1.x7.A VSREF 0.615623f $ **FLOATING
C542 single_10b_cdac_0.x3[0].x1.x9.A VSREF 2.26866f $ **FLOATING
C543 single_10b_cdac_0.x3[0].x1.x11.A VSREF 2.51762f $ **FLOATING
C544 single_10b_cdac_0.x3[0].x2.swp VSREF 15.4802f $ **FLOATING
C545 single_10b_cdac_0.x3[1].x1.x3.Y VSREF 0.60393f $ **FLOATING
C546 single_10b_cdac_0.x3[1].x1.x8.A VSREF 2.14748f $ **FLOATING
C547 single_10b_cdac_0.x3[1].x1.x5.A VSREF 0.736451f $ **FLOATING
C548 single_10b_cdac_0.x3[1].x1.x7.A VSREF 0.615623f $ **FLOATING
C549 single_10b_cdac_0.x3[1].x1.x9.A VSREF 2.26866f $ **FLOATING
C550 single_10b_cdac_0.x3[1].x1.x11.A VSREF 2.51762f $ **FLOATING
C551 single_10b_cdac_0.x3[1].x2.swp VSREF 15.4802f $ **FLOATING
C552 single_10b_cdac_0.x4[2].x1.x3.Y VSREF 0.60393f $ **FLOATING
C553 single_10b_cdac_0.x4[2].x1.x8.A VSREF 2.14748f $ **FLOATING
C554 single_10b_cdac_0.x4[2].x1.x5.A VSREF 0.736451f $ **FLOATING
C555 single_10b_cdac_0.x4[2].x1.x7.A VSREF 0.615623f $ **FLOATING
C556 single_10b_cdac_0.x4[2].x1.x9.A VSREF 2.26866f $ **FLOATING
C557 single_10b_cdac_0.x4[2].x1.x11.A VSREF 2.51762f $ **FLOATING
C558 single_10b_cdac_0.x4[2].x2.swp VSREF 9.69516f $ **FLOATING
C559 single_10b_cdac_0.x4[3].x1.x3.Y VSREF 0.60393f $ **FLOATING
C560 single_10b_cdac_0.x4[3].x1.x8.A VSREF 2.14748f $ **FLOATING
C561 single_10b_cdac_0.x4[3].x1.x5.A VSREF 0.736451f $ **FLOATING
C562 single_10b_cdac_0.x4[3].x1.x7.A VSREF 0.615623f $ **FLOATING
C563 single_10b_cdac_0.x4[3].x1.x9.A VSREF 2.26866f $ **FLOATING
C564 single_10b_cdac_0.x4[3].x1.x11.A VSREF 2.51762f $ **FLOATING
C565 single_10b_cdac_0.x4[3].x2.swp VSREF 9.69516f $ **FLOATING
C566 single_10b_cdac_0.x6[4].x1.x3.Y VSREF 0.60393f $ **FLOATING
C567 single_10b_cdac_0.x6[4].x1.x8.A VSREF 2.14748f $ **FLOATING
C568 single_10b_cdac_0.x6[4].x1.x5.A VSREF 0.736451f $ **FLOATING
C569 single_10b_cdac_0.x6[4].x1.x7.A VSREF 0.615623f $ **FLOATING
C570 single_10b_cdac_0.x6[4].x1.x9.A VSREF 2.26866f $ **FLOATING
C571 single_10b_cdac_0.x6[4].x1.x11.A VSREF 2.51762f $ **FLOATING
C572 single_10b_cdac_0.x6[4].x2.swp VSREF 6.80262f $ **FLOATING
C573 single_10b_cdac_0.x6[5].x1.x3.Y VSREF 0.60393f $ **FLOATING
C574 single_10b_cdac_0.x6[5].x1.x8.A VSREF 2.14748f $ **FLOATING
C575 single_10b_cdac_0.x6[5].x1.x5.A VSREF 0.736451f $ **FLOATING
C576 single_10b_cdac_0.x6[5].x1.x7.A VSREF 0.615623f $ **FLOATING
C577 single_10b_cdac_0.x6[5].x1.x9.A VSREF 2.26866f $ **FLOATING
C578 single_10b_cdac_0.x6[5].x1.x11.A VSREF 2.51762f $ **FLOATING
C579 single_10b_cdac_0.x6[5].x2.swp VSREF 6.80262f $ **FLOATING
C580 single_10b_cdac_0.x8[6].x1.x3.Y VSREF 0.60393f $ **FLOATING
C581 single_10b_cdac_0.x8[6].x1.x8.A VSREF 2.14748f $ **FLOATING
C582 single_10b_cdac_0.x8[6].x1.x5.A VSREF 0.736451f $ **FLOATING
C583 single_10b_cdac_0.x8[6].x1.x7.A VSREF 0.615623f $ **FLOATING
C584 single_10b_cdac_0.x8[6].x1.x9.A VSREF 2.26866f $ **FLOATING
C585 single_10b_cdac_0.x8[6].x1.x11.A VSREF 2.51762f $ **FLOATING
C586 single_10b_cdac_0.x8[6].x2.swp VSREF 5.35635f $ **FLOATING
C587 single_10b_cdac_0.x8[7].x1.x3.Y VSREF 0.60393f $ **FLOATING
C588 single_10b_cdac_0.x8[7].x1.x8.A VSREF 2.14748f $ **FLOATING
C589 single_10b_cdac_0.x8[7].x1.x5.A VSREF 0.736451f $ **FLOATING
C590 single_10b_cdac_0.x8[7].x1.x7.A VSREF 0.615623f $ **FLOATING
C591 single_10b_cdac_0.x8[7].x1.x9.A VSREF 2.26866f $ **FLOATING
C592 single_10b_cdac_0.x8[7].x1.x11.A VSREF 2.51762f $ **FLOATING
C593 single_10b_cdac_0.x8[7].x2.swp VSREF 5.35635f $ **FLOATING
C594 single_10b_cdac_0.x10[8].x1.x3.Y VSREF 0.60393f $ **FLOATING
C595 single_10b_cdac_0.x10[8].x1.x8.A VSREF 2.14748f $ **FLOATING
C596 single_10b_cdac_0.x10[8].x1.x5.A VSREF 0.736451f $ **FLOATING
C597 single_10b_cdac_0.x10[8].x1.x7.A VSREF 0.615623f $ **FLOATING
C598 single_10b_cdac_0.x10[8].x1.x9.A VSREF 2.26866f $ **FLOATING
C599 single_10b_cdac_0.x10[8].x1.x11.A VSREF 2.51762f $ **FLOATING
C600 single_10b_cdac_0.x10[8].x2.swp VSREF 4.63322f $ **FLOATING
C601 single_10b_cdac_0.cdac_sw_1_2.x1.x3.Y VSREF 0.60393f $ **FLOATING
C602 single_10b_cdac_0.cdac_sw_1_2.x1.x8.A VSREF 2.14748f $ **FLOATING
C603 single_10b_cdac_0.cdac_sw_1_2.x1.x5.A VSREF 0.736451f $ **FLOATING
C604 single_10b_cdac_0.cdac_sw_1_2.x1.x7.A VSREF 0.615623f $ **FLOATING
C605 single_10b_cdac_0.cdac_sw_1_2.x1.x9.A VSREF 2.26866f $ **FLOATING
C606 single_10b_cdac_0.cdac_sw_1_2.x1.x11.A VSREF 2.51762f $ **FLOATING
C607 single_10b_cdac_0.cdac_sw_1_2.x2.swp VSREF 4.63322f $ **FLOATING
C608 single_10b_cdac_1.x3[0].x1.x3.Y VSREF 0.60393f $ **FLOATING
C609 single_10b_cdac_1.x3[0].x1.x8.A VSREF 2.14748f $ **FLOATING
C610 single_10b_cdac_1.x3[0].x1.x5.A VSREF 0.736451f $ **FLOATING
C611 single_10b_cdac_1.x3[0].x1.x7.A VSREF 0.615623f $ **FLOATING
C612 single_10b_cdac_1.x3[0].x1.x9.A VSREF 2.26866f $ **FLOATING
C613 single_10b_cdac_1.x3[0].x1.x11.A VSREF 2.51762f $ **FLOATING
C614 single_10b_cdac_1.x3[0].x2.swp VSREF 15.4802f $ **FLOATING
C615 single_10b_cdac_1.x3[1].x1.x3.Y VSREF 0.60393f $ **FLOATING
C616 single_10b_cdac_1.x3[1].x1.x8.A VSREF 2.14748f $ **FLOATING
C617 single_10b_cdac_1.x3[1].x1.x5.A VSREF 0.736451f $ **FLOATING
C618 single_10b_cdac_1.x3[1].x1.x7.A VSREF 0.615623f $ **FLOATING
C619 single_10b_cdac_1.x3[1].x1.x9.A VSREF 2.26866f $ **FLOATING
C620 single_10b_cdac_1.x3[1].x1.x11.A VSREF 2.51762f $ **FLOATING
C621 single_10b_cdac_1.x3[1].x2.swp VSREF 15.4802f $ **FLOATING
C622 single_10b_cdac_1.x4[2].x1.x3.Y VSREF 0.60393f $ **FLOATING
C623 single_10b_cdac_1.x4[2].x1.x8.A VSREF 2.14748f $ **FLOATING
C624 single_10b_cdac_1.x4[2].x1.x5.A VSREF 0.736451f $ **FLOATING
C625 single_10b_cdac_1.x4[2].x1.x7.A VSREF 0.615623f $ **FLOATING
C626 single_10b_cdac_1.x4[2].x1.x9.A VSREF 2.26866f $ **FLOATING
C627 single_10b_cdac_1.x4[2].x1.x11.A VSREF 2.51762f $ **FLOATING
C628 single_10b_cdac_1.x4[2].x2.swp VSREF 9.69516f $ **FLOATING
C629 single_10b_cdac_1.x4[3].x1.x3.Y VSREF 0.60393f $ **FLOATING
C630 single_10b_cdac_1.x4[3].x1.x8.A VSREF 2.14748f $ **FLOATING
C631 single_10b_cdac_1.x4[3].x1.x5.A VSREF 0.736451f $ **FLOATING
C632 single_10b_cdac_1.x4[3].x1.x7.A VSREF 0.615623f $ **FLOATING
C633 single_10b_cdac_1.x4[3].x1.x9.A VSREF 2.26866f $ **FLOATING
C634 single_10b_cdac_1.x4[3].x1.x11.A VSREF 2.51762f $ **FLOATING
C635 single_10b_cdac_1.x4[3].x2.swp VSREF 9.69516f $ **FLOATING
C636 single_10b_cdac_1.x6[4].x1.x3.Y VSREF 0.60393f $ **FLOATING
C637 single_10b_cdac_1.x6[4].x1.x8.A VSREF 2.14748f $ **FLOATING
C638 single_10b_cdac_1.x6[4].x1.x5.A VSREF 0.736451f $ **FLOATING
C639 single_10b_cdac_1.x6[4].x1.x7.A VSREF 0.615623f $ **FLOATING
C640 single_10b_cdac_1.x6[4].x1.x9.A VSREF 2.26866f $ **FLOATING
C641 single_10b_cdac_1.x6[4].x1.x11.A VSREF 2.51762f $ **FLOATING
C642 single_10b_cdac_1.x6[4].x2.swp VSREF 6.80262f $ **FLOATING
C643 single_10b_cdac_1.x6[5].x1.x3.Y VSREF 0.60393f $ **FLOATING
C644 single_10b_cdac_1.x6[5].x1.x8.A VSREF 2.14748f $ **FLOATING
C645 single_10b_cdac_1.x6[5].x1.x5.A VSREF 0.736451f $ **FLOATING
C646 single_10b_cdac_1.x6[5].x1.x7.A VSREF 0.615623f $ **FLOATING
C647 single_10b_cdac_1.x6[5].x1.x9.A VSREF 2.26866f $ **FLOATING
C648 single_10b_cdac_1.x6[5].x1.x11.A VSREF 2.51762f $ **FLOATING
C649 single_10b_cdac_1.x6[5].x2.swp VSREF 6.80262f $ **FLOATING
C650 single_10b_cdac_1.x8[6].x1.x3.Y VSREF 0.60393f $ **FLOATING
C651 single_10b_cdac_1.x8[6].x1.x8.A VSREF 2.14748f $ **FLOATING
C652 single_10b_cdac_1.x8[6].x1.x5.A VSREF 0.736451f $ **FLOATING
C653 single_10b_cdac_1.x8[6].x1.x7.A VSREF 0.615623f $ **FLOATING
C654 single_10b_cdac_1.x8[6].x1.x9.A VSREF 2.26866f $ **FLOATING
C655 single_10b_cdac_1.x8[6].x1.x11.A VSREF 2.51762f $ **FLOATING
C656 single_10b_cdac_1.x8[6].x2.swp VSREF 5.35635f $ **FLOATING
C657 single_10b_cdac_1.x8[7].x1.x3.Y VSREF 0.60393f $ **FLOATING
C658 single_10b_cdac_1.x8[7].x1.x8.A VSREF 2.14748f $ **FLOATING
C659 single_10b_cdac_1.x8[7].x1.x5.A VSREF 0.736451f $ **FLOATING
C660 single_10b_cdac_1.x8[7].x1.x7.A VSREF 0.615623f $ **FLOATING
C661 single_10b_cdac_1.x8[7].x1.x9.A VSREF 2.26866f $ **FLOATING
C662 single_10b_cdac_1.x8[7].x1.x11.A VSREF 2.51762f $ **FLOATING
C663 single_10b_cdac_1.x8[7].x2.swp VSREF 5.35635f $ **FLOATING
C664 single_10b_cdac_1.x10[8].x1.x3.Y VSREF 0.60393f $ **FLOATING
C665 single_10b_cdac_1.x10[8].x1.x8.A VSREF 2.14748f $ **FLOATING
C666 single_10b_cdac_1.x10[8].x1.x5.A VSREF 0.736451f $ **FLOATING
C667 single_10b_cdac_1.x10[8].x1.x7.A VSREF 0.615623f $ **FLOATING
C668 single_10b_cdac_1.x10[8].x1.x9.A VSREF 2.26866f $ **FLOATING
C669 single_10b_cdac_1.x10[8].x1.x11.A VSREF 2.51762f $ **FLOATING
C670 single_10b_cdac_1.x10[8].x2.swp VSREF 4.63322f $ **FLOATING
C671 single_10b_cdac_1.cdac_sw_1_2.x1.x3.Y VSREF 0.60393f $ **FLOATING
C672 single_10b_cdac_1.cdac_sw_1_2.x1.x8.A VSREF 2.14748f $ **FLOATING
C673 single_10b_cdac_1.cdac_sw_1_2.x1.x5.A VSREF 0.736451f $ **FLOATING
C674 single_10b_cdac_1.cdac_sw_1_2.x1.x7.A VSREF 0.615623f $ **FLOATING
C675 single_10b_cdac_1.cdac_sw_1_2.x1.x9.A VSREF 2.26866f $ **FLOATING
C676 single_10b_cdac_1.cdac_sw_1_2.x1.x11.A VSREF 2.51762f $ **FLOATING
C677 single_10b_cdac_1.cdac_sw_1_2.x2.swp VSREF 4.63322f $ **FLOATING
