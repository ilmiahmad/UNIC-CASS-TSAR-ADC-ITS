magic
tech sky130A
magscale 1 2
timestamp 1731350358
<< nwell >>
rect -95 -235 1374 331
rect 9241 -46 10564 331
rect 9241 -220 10200 -46
rect 10302 -220 10564 -46
rect 9241 -224 10213 -220
rect 10280 -224 10564 -220
rect 9241 -235 10564 -224
<< pwell >>
rect -96 388 11046 572
rect 10862 -292 11046 388
rect -96 -476 11046 -292
<< psubdiff >>
rect 5 518 57 544
rect 5 415 57 456
rect 10926 199 10978 249
rect 10926 -155 10978 -106
rect 5 -356 57 -319
rect 5 -449 57 -418
<< nsubdiff >>
rect 5 240 57 264
rect 5 -188 57 -164
rect 10399 249 10451 273
rect 10399 -179 10451 -155
<< psubdiffcont >>
rect 5 456 57 518
rect 10926 -106 10978 199
rect 5 -418 57 -356
<< nsubdiffcont >>
rect 5 -164 57 240
rect 10399 -155 10451 249
<< locali >>
rect 5 518 57 572
rect 5 388 57 456
rect 5 240 57 331
rect 10399 249 10451 331
rect 5 -235 57 -164
rect 10926 199 10978 249
rect 10926 -155 10978 -106
rect 10399 -235 10451 -155
rect 5 -356 57 -291
rect 5 -476 57 -418
<< viali >>
rect 5 456 57 518
rect 5 -164 57 240
rect 9856 -140 9896 -70
rect 10399 -155 10451 249
rect 10926 -106 10978 199
rect 10046 -276 10086 -236
rect 10186 -281 10220 -247
rect 5 -418 57 -356
<< metal1 >>
rect -66 544 178 640
rect 9820 544 10954 640
rect -1 518 63 544
rect -1 456 5 518
rect 57 456 63 518
rect -1 444 63 456
rect -1 240 63 252
rect -1 96 5 240
rect -66 0 5 96
rect -1 -164 5 0
rect 57 96 63 240
rect 10393 249 10457 261
rect 10393 96 10399 249
rect 57 0 178 96
rect 10263 0 10399 96
rect 57 -164 63 0
rect 9850 -70 9902 -58
rect 9840 -140 9850 -70
rect 9902 -140 9912 -70
rect 9850 -152 9902 -140
rect -1 -176 63 -164
rect 10393 -155 10399 0
rect 10451 -155 10457 249
rect 10393 -167 10457 -155
rect 10858 211 10954 544
rect 10858 199 10984 211
rect 10858 -106 10926 199
rect 10978 -106 10984 199
rect 10858 -118 10984 -106
rect 10030 -282 10040 -230
rect 10092 -282 10102 -230
rect 10164 -290 10174 -234
rect 10232 -290 10242 -234
rect -1 -356 63 -344
rect -1 -418 5 -356
rect 57 -418 63 -356
rect -1 -448 63 -418
rect 10858 -448 10954 -118
rect -66 -544 178 -448
rect 10276 -544 10954 -448
<< via1 >>
rect 9850 -140 9856 -70
rect 9856 -140 9896 -70
rect 9896 -140 9902 -70
rect 10040 -236 10092 -230
rect 10040 -276 10046 -236
rect 10046 -276 10086 -236
rect 10086 -276 10092 -236
rect 10040 -282 10092 -276
rect 10174 -247 10232 -234
rect 10174 -281 10186 -247
rect 10186 -281 10220 -247
rect 10220 -281 10232 -247
rect 10174 -290 10232 -281
<< metal2 >>
rect -182 399 216 451
rect 5297 400 5306 456
rect 5362 400 5371 456
rect -179 277 449 327
rect 1936 231 1996 240
rect 1936 162 1996 171
rect 3874 231 3934 240
rect 3874 162 3934 171
rect 452 129 512 138
rect 452 60 512 69
rect 2386 129 2446 138
rect 2386 60 2446 69
rect 4316 129 4376 138
rect 4316 60 4376 69
rect 281 24 341 33
rect 281 -45 341 -36
rect 2213 24 2273 33
rect 2213 -45 2273 -36
rect 4145 27 4205 36
rect 4145 -42 4205 -33
rect 1770 -76 1830 -67
rect 1770 -145 1830 -136
rect 3702 -75 3762 -66
rect 3702 -144 3762 -135
rect 4829 -231 4879 325
rect 5806 231 5866 240
rect 5806 162 5866 171
rect 7738 231 7798 240
rect 7738 162 7798 171
rect 9670 231 9730 240
rect 9670 162 9730 171
rect 6248 129 6308 138
rect 6248 60 6308 69
rect 8180 129 8240 138
rect 8180 60 8240 69
rect 6076 27 6136 36
rect 6076 -42 6136 -33
rect 8014 27 8074 36
rect 8014 -42 8074 -33
rect 9851 -60 9901 -58
rect 5634 -75 5694 -66
rect 5634 -144 5694 -135
rect 7564 -75 7624 -66
rect 7564 -144 7624 -135
rect 9498 -75 9558 -66
rect 9498 -144 9558 -135
rect 9850 -70 9902 -60
rect 9850 -150 9902 -140
rect 9851 -181 9901 -150
rect 9699 -231 9901 -181
rect 10040 -230 10092 -224
rect 5304 -299 5364 -290
rect 5304 -368 5364 -359
rect 10040 -872 10092 -282
rect 10174 -234 10274 -224
rect 10232 -290 10274 -234
rect 10174 -300 10274 -290
rect 10222 -864 10274 -300
<< via2 >>
rect 5306 400 5362 456
rect 1936 171 1996 231
rect 3874 171 3934 231
rect 452 69 512 129
rect 2386 69 2446 129
rect 4316 69 4376 129
rect 281 -36 341 24
rect 2213 -36 2273 24
rect 4145 -33 4205 27
rect 1770 -136 1830 -76
rect 3702 -135 3762 -75
rect 5806 171 5866 231
rect 7738 171 7798 231
rect 9670 171 9730 231
rect 6248 69 6308 129
rect 8180 69 8240 129
rect 6076 -33 6136 27
rect 8014 -33 8074 27
rect 5634 -135 5694 -75
rect 7564 -135 7624 -75
rect 9498 -135 9558 -75
rect 5304 -359 5364 -299
<< metal3 >>
rect 281 29 341 956
rect 1936 236 1996 956
rect 1931 231 2001 236
rect 1931 171 1936 231
rect 1996 171 2001 231
rect 1931 166 2001 171
rect 447 129 517 134
rect 447 69 452 129
rect 512 69 517 129
rect 447 64 517 69
rect 276 24 346 29
rect 276 -36 281 24
rect 341 -36 346 24
rect 276 -41 346 -36
rect 452 -873 512 64
rect 2213 29 2273 956
rect 3874 236 3934 956
rect 3869 231 3939 236
rect 3869 171 3874 231
rect 3934 171 3939 231
rect 3869 166 3939 171
rect 2381 129 2451 134
rect 2381 69 2386 129
rect 2446 69 2451 129
rect 2381 64 2451 69
rect 2208 24 2278 29
rect 2208 -36 2213 24
rect 2273 -36 2278 24
rect 2208 -41 2278 -36
rect 1765 -76 1835 -71
rect 1765 -136 1770 -76
rect 1830 -136 1835 -76
rect 1765 -141 1835 -136
rect 1770 -873 1830 -141
rect 2386 -873 2446 64
rect 4145 32 4205 956
rect 5301 456 5367 461
rect 5301 400 5306 456
rect 5362 400 5367 456
rect 5301 395 5367 400
rect 4311 129 4381 134
rect 4311 69 4316 129
rect 4376 69 4381 129
rect 4311 64 4381 69
rect 4140 27 4210 32
rect 4140 -33 4145 27
rect 4205 -33 4210 27
rect 4140 -38 4210 -33
rect 3697 -75 3767 -70
rect 3697 -135 3702 -75
rect 3762 -135 3767 -75
rect 3697 -140 3767 -135
rect 3702 -873 3762 -140
rect 4316 -873 4376 64
rect 5304 -294 5364 395
rect 5806 236 5866 956
rect 5801 231 5871 236
rect 5801 171 5806 231
rect 5866 171 5871 231
rect 5801 166 5871 171
rect 6076 32 6136 956
rect 7738 236 7798 956
rect 7733 231 7803 236
rect 7733 171 7738 231
rect 7798 171 7803 231
rect 7733 166 7803 171
rect 6243 129 6313 134
rect 6243 69 6248 129
rect 6308 69 6313 129
rect 6243 64 6313 69
rect 6071 27 6141 32
rect 6071 -33 6076 27
rect 6136 -33 6141 27
rect 6071 -38 6141 -33
rect 5629 -75 5699 -70
rect 5629 -135 5634 -75
rect 5694 -135 5699 -75
rect 5629 -140 5699 -135
rect 5299 -299 5369 -294
rect 5299 -359 5304 -299
rect 5364 -359 5369 -299
rect 5299 -364 5369 -359
rect 5634 -873 5694 -140
rect 6248 -873 6308 64
rect 8014 32 8074 956
rect 9670 236 9730 956
rect 9665 231 9735 236
rect 9665 171 9670 231
rect 9730 171 9735 231
rect 9665 166 9735 171
rect 8175 129 8245 134
rect 8175 69 8180 129
rect 8240 69 8245 129
rect 8175 64 8245 69
rect 8009 27 8079 32
rect 8009 -33 8014 27
rect 8074 -33 8079 27
rect 8009 -38 8079 -33
rect 7559 -75 7629 -70
rect 7559 -135 7564 -75
rect 7624 -135 7629 -75
rect 7559 -140 7629 -135
rect 7564 -873 7624 -140
rect 8180 -873 8240 64
rect 9493 -75 9563 -70
rect 9493 -135 9498 -75
rect 9558 -135 9563 -75
rect 9493 -140 9563 -135
rect 9498 -872 9558 -140
use and_latch  and_latch_0
timestamp 1731349849
transform -1 0 29994 0 1 -16
box 19662 -528 20198 112
use flip_flop_5_latch  flip_flop_5_latch_0
timestamp 1731349849
transform 1 0 342 0 -1 -974
box -205 -1614 9531 -974
use flip_flop_5_latch  flip_flop_5_latch_1
timestamp 1731349849
transform -1 0 9668 0 1 1070
box -205 -1614 9531 -974
<< labels >>
flabel metal2 10250 -850 10250 -850 0 FreeSans 800 0 0 0 FINAL
port 0 nsew
flabel metal2 10066 -754 10066 -754 0 FreeSans 800 0 0 0 CLKS
port 1 nsew
flabel metal1 -54 -504 -54 -504 0 FreeSans 800 0 0 0 VSSD
port 2 nsew
flabel metal1 -54 48 -54 48 0 FreeSans 800 0 0 0 VDDD
port 3 nsew
flabel metal2 -164 424 -164 424 0 FreeSans 800 0 0 0 EN
port 4 nsew
flabel metal2 -170 290 -170 290 0 FreeSans 800 0 0 0 CK
port 5 nsew
flabel metal3 1962 930 1968 930 0 FreeSans 800 0 0 0 DOUT[1]
port 8 nsew
flabel metal3 2248 718 2254 718 0 FreeSans 800 0 0 0 DOUT[2]
port 9 nsew
flabel metal3 3904 936 3910 936 0 FreeSans 800 0 0 0 DOUT[3]
port 10 nsew
flabel metal3 4176 714 4182 714 0 FreeSans 800 0 0 0 DOUT[4]
port 11 nsew
flabel metal3 5834 930 5840 930 0 FreeSans 800 0 0 0 DOUT[5]
port 12 nsew
flabel metal3 6110 712 6116 712 0 FreeSans 800 0 0 0 DOUT[6]
port 13 nsew
flabel metal3 7758 918 7764 918 0 FreeSans 800 0 0 0 DOUT[7]
port 14 nsew
flabel metal3 8044 714 8050 714 0 FreeSans 800 0 0 0 DOUT[8]
port 15 nsew
flabel metal3 9696 922 9702 922 0 FreeSans 800 0 0 0 DOUT[9]
port 16 nsew
flabel metal3 1802 -828 1802 -828 0 FreeSans 800 0 0 0 SWP[0]
port 17 nsew
flabel metal3 474 -846 474 -846 0 FreeSans 800 0 0 0 SWP[1]
port 18 nsew
flabel metal3 3736 -832 3736 -832 0 FreeSans 800 0 0 0 SWP[2]
port 19 nsew
flabel metal3 2412 -836 2412 -836 0 FreeSans 800 0 0 0 SWP[3]
port 20 nsew
flabel metal3 5666 -848 5666 -848 0 FreeSans 800 0 0 0 SWP[4]
port 21 nsew
flabel metal3 4342 -834 4342 -834 0 FreeSans 800 0 0 0 SWP[5]
port 22 nsew
flabel metal3 7598 -848 7598 -848 0 FreeSans 800 0 0 0 SWP[6]
port 23 nsew
flabel metal3 6278 -838 6278 -838 0 FreeSans 800 0 0 0 SWP[7]
port 24 nsew
flabel metal3 9528 -846 9528 -846 0 FreeSans 800 0 0 0 SWP[8]
port 25 nsew
flabel metal3 8212 -852 8212 -838 0 FreeSans 800 0 0 0 SWP[9]
port 26 nsew
flabel metal3 314 924 314 938 0 FreeSans 800 0 0 0 DOUT[0]
port 27 nsew
flabel metal1 -28 598 -28 598 0 FreeSans 800 0 0 0 VSSD
port 28 nsew
<< end >>
