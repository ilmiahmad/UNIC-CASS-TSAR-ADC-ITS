* PEX produced on Jum 08 Nov 2024 03:54:37  CST using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from sar.ext - technology: sky130A

.subckt sar CKO DOUT[0] DOUT[1] DOUT[2] DOUT[3] DOUT[4] DOUT[5] DOUT[6] DOUT[7] DOUT[8]
+ DOUT[9] CLKS CLKSB CLK EN VSSD VDDD CF[0] CF[1] CF[2] CF[3] CF[4] CF[5] CF[6] CF[7]
+ CF[8] CF[9] SWP[9] SWP[8] SWP[7] SWP[6] SWP[5] SWP[4] SWP[3] SWP[2] SWP[1] SWP[0]
+ SWN[9] SWN[8] SWN[7] SWN[6] SWN[5] SWN[4] SWN[3] SWN[2] SWN[1] SWN[0] COMP_P COMP_N
X0 VDDD.t1069 a_7068_n1029.t4 a_7243_n1055.t2 VDDD.t1068 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_n1085_3923.t2 a_n1709_3557.t2 a_n1193_3557.t2 VDDD.t1133 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2 a_n4691_n10054.t2 a_n4909_n9650.t4 VDDD.t724 VDDD.t723 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3 VSSD.t1111 CLKS.t16 a_n2715_n9662.t0 VSSD.t1053 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_5624_n5650.t1 a_5911_n5372.t4 VDDD.t228 VDDD.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X5 a_3236_3557.t2 a_2155_3557.t2 a_2889_3799.t3 VDDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6 a_4679_n663.t2 CLKS.t17 VDDD.t545 VDDD.t544 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X7 a_8520_n9662.t2 cdac_ctrl_0.x2.X.t16 VSSD.t936 VSSD.t897 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X8 out_latch_0.FINAL.t15 a_n784_n1599.t6 VDDD.t672 VDDD.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VSSD.t421 a_8160_n5482.t2 a_8121_n5356.t0 VSSD.t420 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 a_855_n1331.t1 CLK.t0 VDDD.t694 VDDD.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 VSSD.t54 a_7274_2691.t3 auto_sampling_0.x21.D.t1 VSSD.t53 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VSSD.t245 a_n10393_n10028.t6 cdac_ctrl_0.x2.X.t0 VSSD.t193 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_6779_n9484.t1 a_6333_n9484.t2 a_6683_n9484.t1 VSSD.t443 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X14 a_n8555_n9242.t3 a_n8773_n9484.t4 VDDD.t382 VDDD.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X15 VDDD.t763 a_4452_n5387.t4 a_4383_n5258.t2 VDDD.t762 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X16 a_2830_n5624.t0 a_2451_n5258.t4 a_2758_n5624.t0 VSSD.t52 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 VDDD.t1078 a_4713_n4702.t4 a_4888_n4776.t1 VDDD.t1077 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_n480_n9650.t0 a_n1395_n10022.t2 a_n827_n10054.t0 VSSD.t775 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X19 DOUT[0].t3 a_n172_n5650.t3 VDDD.t811 VDDD.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VSSD.t1163 a_n454_2691.t3 auto_sampling_0.x22.A.t1 VSSD.t1162 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_1011_n5080.t0 a_n66_n5074.t2 a_849_n4702.t0 VDDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 a_995_n9118.t0 a_371_n9484.t2 a_887_n9484.t0 VDDD.t1402 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X23 a_n1193_3557.t0 a_n1543_3557.t2 a_n1288_3557.t0 VDDD.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X24 VSSD.t735 a_n305_n9510.t3 a_n371_n9484.t1 VSSD.t137 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_n2869_n10028.t2 CLKS.t18 VDDD.t547 VDDD.t546 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 a_n8665_n9118.t2 CLKS.t19 VDDD.t631 VDDD.t630 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X27 a_1626_n1029.t1 CLKS.t20 VSSD.t1110 VSSD.t1109 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X28 a_3397_3083.t0 a_2320_2717.t2 a_3235_2717.t1 VDDD.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 VDDD.t1059 EN.t0 a_4597_n5258.t0 VDDD.t1058 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X30 VSSD.t392 a_8583_n1331.t2 a_8544_n1457.t0 VSSD.t391 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 VSSD.t342 a_1479_3531.t3 a_1413_3557.t0 VSSD.t341 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X32 a_5311_n1055.t2 CLKS.t21 VDDD.t633 VDDD.t632 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X33 a_8615_n9650.t1 a_8099_n10022.t2 a_8520_n9662.t0 VSSD.t23 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X34 a_7843_n5372.t0 a_8121_n5356.t2 a_8077_n5258.t1 VDDD.t1284 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X35 a_n975_3799.t2 a_n1193_3557.t4 VSSD.t844 VSSD.t843 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X36 VSSD.t559 CLK.t1 a_2155_3557.t1 VSSD.t558 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X37 a_6754_n4702.t0 a_5564_n5074.t2 a_6645_n4702.t1 VSSD.t490 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X38 CF[5].t3 a_9175_n1055.t3 VDDD.t1230 VDDD.t1229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X39 a_8466_2717.t1 a_7950_2717.t2 a_8371_2717.t0 VSSD.t923 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X40 VSSD.t5 CF[4].t4 a_n1561_n10022.t0 VSSD.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X41 VDDD.t918 CF[8].t4 a_6167_n10022.t1 VDDD.t917 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X42 CF[3].t3 a_6047_n1599.t3 VDDD.t1076 VDDD.t1075 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X43 a_4969_n9242.t1 a_4751_n9484.t4 VDDD.t1228 VDDD.t1227 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X44 VDDD.t1127 a_502_n5106.t4 a_392_n5080.t2 VDDD.t1126 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X45 VSSD.t216 a_1447_n1055.t3 a_1381_n1029.t0 VSSD.t215 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X46 VDDD.t1101 a_1024_n4776.t3 a_1011_n5080.t1 VDDD.t1100 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X47 a_n937_n10028.t2 CLKS.t22 VDDD.t635 VDDD.t634 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X48 a_5425_n9650.t0 a_4235_n10022.t2 a_5316_n9650.t0 VSSD.t149 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X49 a_6947_n5258.t0 a_6189_n5356.t2 a_6384_n5387.t1 VDDD.t1191 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X50 a_n1097_3557.t0 a_n1543_3557.t3 a_n1193_3557.t1 VSSD.t238 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X51 a_2889_3799.t0 a_2671_3557.t4 VDDD.t351 VDDD.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X52 a_n4691_n10054.t3 a_n4909_n9650.t5 VSSD.t835 VSSD.t834 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X53 VDDD.t1061 EN.t1 a_3692_n5650.t0 VDDD.t1060 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X54 VDDD.t283 CF[9].t4 a_8099_n10022.t0 VDDD.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X55 a_n628_3557.t1 a_n1543_3557.t4 a_n975_3799.t0 VSSD.t239 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X56 a_8752_n4776.t2 a_8577_n4702.t4 a_8931_n4714.t1 VSSD.t242 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X57 VSSD.t105 SWP[4].t4 a_5015_n5258.t0 VSSD.t104 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X58 a_5343_3531.t0 EN.t2 VDDD.t1063 VDDD.t1062 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X59 CLKS.t4 auto_sampling_0.x24.A.t8 VSSD.t211 VSSD.t210 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X60 VDDD.t419 a_2888_2959.t4 a_2778_3083.t1 VDDD.t418 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X61 a_n8868_n9662.t3 cdac_ctrl_0.x2.X.t17 VDDD.t1184 VDDD.t1183 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X62 VDDD.t1242 a_4888_n4776.t3 DOUT[5].t3 VDDD.t1241 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X63 a_7068_n1029.t0 a_5987_n1029.t2 a_6721_n787.t3 VDDD.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X64 auto_sampling_0.x21.Q.t3 a_9206_2691.t3 VDDD.t404 VDDD.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X65 VSSD.t827 EN.t3 a_4864_2717.t0 VSSD.t826 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X66 a_815_n663.t2 CLKS.t23 VDDD.t637 VDDD.t636 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X67 VDDD.t226 auto_sampling_0.x24.A.t9 CLKS.t5 VDDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X68 a_6440_3557.t3 auto_sampling_0.x5.D.t4 VDDD.t817 VDDD.t816 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X69 a_n6841_n9484.t2 a_n7357_n9484.t2 a_n6936_n9484.t1 VSSD.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X70 a_8230_n5106.t2 a_8012_n4702.t4 VSSD.t477 VSSD.t476 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X71 VSSD.t1108 CLKS.t24 a_2505_n1207.t1 VSSD.t1107 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X72 VDDD.t809 a_4969_n10054.t4 a_4859_n10028.t1 VDDD.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X73 a_n6733_n9118.t0 a_n7357_n9484.t3 a_n6841_n9484.t1 VDDD.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X74 a_2520_n5387.t1 a_2364_n5482.t2 a_2665_n5258.t2 VDDD.t628 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X75 a_n2715_n9662.t1 a_n2759_n10054.t4 a_n2881_n9650.t1 VSSD.t142 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X76 CF[9].t1 a_1447_n1055.t4 VSSD.t218 VSSD.t217 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X77 a_n6167_n9650.t1 a_n7357_n10022.t2 a_n6276_n9650.t3 VSSD.t520 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X78 a_6945_n9662.t0 a_6901_n10054.t4 a_6779_n9650.t0 VSSD.t505 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X79 a_2478_n4714.t1 a_2434_n5106.t4 a_2312_n4702.t0 VSSD.t197 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X80 VSSD.t873 a_n6101_n9724.t3 SWN[1].t1 VSSD.t684 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X81 a_4667_n1029.t0 a_4221_n1029.t2 a_4571_n1029.t1 VSSD.t757 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X82 a_9180_n9484.t1 a_8099_n9484.t2 a_8833_n9242.t1 VDDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X83 VDDD.t798 a_n4691_n9242.t4 a_n4801_n9118.t0 VDDD.t797 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X84 a_9487_n5472.t0 out_latch_0.FINAL.t16 a_9661_n5596.t0 VSSD.t759 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X85 VSSD.t1137 a_3379_n1055.t3 CF[8].t1 VSSD.t1136 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X86 a_6047_n1599.t1 a_6334_n1441.t4 VDDD.t800 VDDD.t799 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X87 VDDD.t1222 SWP[8].t4 a_8879_n5258.t1 VDDD.t1221 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X88 a_7275_3531.t1 a_7100_3557.t4 a_7454_3557.t1 VSSD.t99 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X89 VDDD.t677 a_5311_n1055.t3 a_5298_n663.t0 VDDD.t676 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X90 VDDD.t244 a_n2237_n9510.t3 a_n2250_n9118.t0 VDDD.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X91 VSSD.t780 a_3411_3531.t3 auto_sampling_0.x3.D.t1 VSSD.t779 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X92 a_6645_n4702.t2 a_5730_n5074.t2 a_6298_n5106.t2 VSSD.t576 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X93 VSSD.t496 a_855_n1331.t2 a_816_n1457.t0 VSSD.t495 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X94 a_n4182_n9118.t0 a_n5259_n9484.t2 a_n4344_n9484.t1 VDDD.t593 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X95 a_4401_n9484.t0 a_4235_n9484.t2 VSSD.t739 VSSD.t436 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X96 CF[8].t2 a_3379_n1055.t4 VDDD.t1366 VDDD.t1365 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X97 a_7100_3557.t3 a_6019_3557.t2 a_6753_3799.t2 VDDD.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X98 a_847_3923.t0 EN.t4 VDDD.t1065 VDDD.t1064 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X99 a_6738_n1573.t0 a_6651_n1331.t2 a_6334_n1441.t0 VDDD.t697 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X100 a_4806_n1573.t3 a_4680_n1457.t2 a_4402_n1441.t1 VSSD.t995 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X101 a_5316_n9650.t2 a_4401_n10022.t2 a_4969_n10054.t2 VSSD.t534 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X102 VDDD.t551 a_n480_n9484.t4 a_n305_n9510.t0 VDDD.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X103 VSSD.t1106 CLKS.t25 a_n4647_n9662.t1 VSSD.t1047 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X104 a_380_n4702.t0 a_n66_n5074.t3 a_284_n4702.t0 VSSD.t563 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X105 a_9302_n1573.t0 a_8583_n1331.t3 a_8739_n1599.t1 VSSD.t393 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X106 SWN[5].t1 a_1627_n9724.t3 VSSD.t958 VSSD.t585 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X107 a_644_3557.t2 auto_sampling_0.x7.Q.t4 VSSD.t583 VSSD.t582 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X108 VSSD.t448 CF[5].t4 a_371_n10022.t0 VSSD.t447 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X109 VSSD.t1115 CKO.t4 a_3632_n5074.t0 VSSD.t1114 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X110 a_4888_n4776.t0 EN.t5 VDDD.t176 VDDD.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X111 SWP[7].t1 a_5491_n9510.t3 VSSD.t565 VSSD.t564 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X112 VDDD.t609 a_1304_3557.t4 a_1479_3531.t1 VDDD.t608 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X113 a_4603_3557.t1 a_4087_3557.t2 a_4508_3557.t0 VSSD.t675 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X114 a_n8208_n9650.t0 a_n9123_n10022.t2 a_n8555_n10054.t1 VSSD.t787 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X115 a_2787_n1331.t1 CLK.t2 VDDD.t826 VDDD.t825 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X116 VDDD.t575 a_5343_3531.t3 a_5330_3923.t1 VDDD.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X117 a_n7191_n10022.t0 a_n7357_n10022.t3 VSSD.t522 VSSD.t521 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 a_n4169_n9724.t2 CLKS.t26 VDDD.t514 VDDD.t513 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X119 VDDD.t828 CLK.t3 a_4055_n1029.t1 VDDD.t827 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X120 VSSD.t136 a_n8033_n9510.t3 a_n8099_n9484.t1 VSSD.t7 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X121 cdac_ctrl_0.x1.X.t7 a_n10393_n9484.t6 VSSD.t192 VSSD.t191 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X122 a_5730_n5074.t0 a_5564_n5074.t3 VSSD.t492 VSSD.t491 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 a_n2237_n9724.t0 a_n2412_n9650.t4 a_n2058_n9662.t0 VSSD.t380 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X124 a_n2250_n10028.t1 a_n3327_n10022.t2 a_n2412_n9650.t1 VDDD.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X125 a_9175_n1055.t1 CLKS.t27 VDDD.t516 VDDD.t515 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X126 a_8077_n5258.t0 a_7556_n5650.t3 VDDD.t150 VDDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X127 a_2888_2959.t1 a_2670_2717.t4 VSSD.t929 VSSD.t928 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X128 a_3558_n1029.t1 CLKS.t28 VSSD.t1105 VSSD.t1104 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X129 a_1272_n1029.t0 a_191_n1029.t2 a_925_n787.t0 VDDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X130 auto_sampling_0.x15.D.t3 a_3410_2691.t3 VDDD.t1030 VDDD.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X131 a_n628_3557.t3 a_n1709_3557.t3 a_n975_3799.t1 VDDD.t589 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X132 a_9031_2717.t3 a_8116_2717.t2 a_8684_2959.t3 VSSD.t337 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X133 a_9355_n9510.t0 a_9180_n9484.t4 a_9534_n9484.t0 VSSD.t519 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X134 SWP[7].t3 a_5491_n9510.t4 VDDD.t700 VDDD.t699 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X135 a_5316_n9650.t1 a_4235_n10022.t3 a_4969_n10054.t0 VDDD.t497 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X136 a_5491_n9510.t2 CLKS.t29 VDDD.t1269 VDDD.t1268 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X137 cdac_ctrl_0.x1.X.t15 a_n10393_n9484.t7 VDDD.t212 VDDD.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X138 a_6753_3799.t3 a_6535_3557.t4 VDDD.t683 VDDD.t682 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X139 a_7357_n9650.t1 a_6167_n10022.t2 a_7248_n9650.t1 VSSD.t200 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X140 SWN[9].t3 a_9355_n9724.t3 VDDD.t118 VDDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X141 a_1479_3531.t2 a_1304_3557.t5 a_1658_3557.t1 VSSD.t504 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X142 a_8833_n10054.t3 a_8615_n9650.t4 VDDD.t1108 VDDD.t1107 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X143 a_2943_n1599.t1 a_2787_n1331.t2 a_3088_n1573.t0 VDDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X144 a_n6623_n10054.t0 a_n6841_n9650.t4 VSSD.t984 VSSD.t404 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X145 VDDD.t178 EN.t6 a_5624_n5650.t0 VDDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 a_9207_3531.t0 EN.t7 VDDD.t180 VDDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X147 DOUT[5].t2 a_4888_n4776.t4 VDDD.t1244 VDDD.t1243 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X148 a_4677_n1207.t1 a_4115_n1599.t3 VSSD.t966 VSSD.t965 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X149 a_772_n1573.t1 a_251_n1599.t3 VDDD.t1143 VDDD.t1142 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X150 VDDD.t1271 CLKS.t30 a_3088_n1573.t2 VDDD.t1270 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X151 a_1614_n9118.t0 a_537_n9484.t2 a_1452_n9484.t2 VDDD.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X152 a_4402_n1441.t3 a_4719_n1331.t2 a_4677_n1207.t0 VSSD.t972 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X153 VDDD.t534 CF[5].t5 a_9302_n1573.t3 VDDD.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X154 VDDD.t1399 a_n454_2691.t4 a_n467_3083.t0 VDDD.t1398 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X155 VSSD.t636 a_n172_n5650.t4 DOUT[0].t1 VSSD.t635 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X156 VDDD.t33 a_3559_n9510.t3 a_3546_n9118.t1 VDDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X157 a_n8773_n9484.t0 a_n9289_n9484.t2 a_n8868_n9484.t0 VSSD.t116 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X158 a_1574_n1573.t3 a_855_n1331.t3 a_1011_n1599.t3 VSSD.t497 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X159 VDDD.t942 a_8752_n4776.t3 a_8739_n5080.t0 VDDD.t941 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X160 CF[8].t3 a_3379_n1055.t5 VSSD.t1139 VSSD.t1138 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X161 a_n8099_n9650.t0 a_n9289_n10022.t2 a_n8208_n9650.t3 VSSD.t630 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X162 a_6721_n787.t0 a_6503_n1029.t4 VSSD.t40 VSSD.t39 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X163 VDDD.t1338 a_1105_n9242.t4 a_995_n9118.t2 VDDD.t1337 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X164 VSSD.t165 EN.t8 a_546_n4714.t0 VSSD.t164 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X165 VDDD.t1232 a_9175_n1055.t4 a_9162_n663.t0 VDDD.t1231 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X166 a_1321_n1207.t1 a_942_n1573.t4 a_1249_n1207.t0 VSSD.t712 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X167 VDDD.t1057 a_6298_n5106.t4 a_6188_n5080.t2 VDDD.t1056 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X168 VSSD.t752 a_8752_n4776.t4 DOUT[9].t1 VSSD.t751 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X169 VSSD.t1 CF[4].t5 a_7370_n1573.t1 VSSD.t0 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X170 a_n2759_n9242.t2 a_n2977_n9484.t4 VSSD.t63 VSSD.t34 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X171 SWP[1].t1 a_n6101_n9510.t3 VSSD.t348 VSSD.t288 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X172 VDDD.t1379 a_n6623_n9242.t4 a_n6733_n9118.t2 VDDD.t1378 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X173 a_2665_n5258.t1 a_2451_n5258.t5 VDDD.t47 VDDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X174 a_5670_n9662.t1 CLKS.t31 VSSD.t1103 VSSD.t1039 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X175 a_1203_n4714.t1 EN.t9 VSSD.t167 VSSD.t166 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X176 a_8723_n10028.t0 a_8099_n10022.t3 a_8615_n9650.t0 VDDD.t947 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X177 VSSD.t101 a_7275_3531.t3 auto_sampling_0.x11.D.t1 VSSD.t100 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X178 VDDD.t398 a_n4169_n9510.t3 a_n4182_n9118.t1 VDDD.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X179 a_3379_n1055.t2 CLKS.t32 VDDD.t1273 VDDD.t1272 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X180 VSSD.t230 CF[7].t4 a_4235_n9484.t0 VSSD.t229 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X181 VSSD.t144 a_7556_n5650.t4 DOUT[8].t1 VSSD.t143 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X182 a_3546_n10028.t1 a_2469_n10022.t2 a_3384_n9650.t3 VDDD.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X183 VSSD.t892 a_n453_3531.t3 auto_sampling_0.x7.Q.t0 VSSD.t891 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X184 VDDD.t316 a_n6101_n9724.t4 a_n6114_n10028.t1 VDDD.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X185 a_n2412_n9650.t2 a_n3493_n10022.t2 a_n2759_n10054.t2 VDDD.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X186 CLKS.t6 auto_sampling_0.x24.A.t10 VSSD.t213 VSSD.t212 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X187 a_n1085_3923.t0 EN.t10 VDDD.t182 VDDD.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X188 VDDD.t441 a_8583_n1331.t4 a_8544_n1457.t1 VDDD.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X189 a_n305_n9510.t1 a_n480_n9484.t5 a_n126_n9484.t0 VSSD.t273 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X190 a_6333_n9484.t1 a_6167_n9484.t2 VSSD.t997 VSSD.t202 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X191 a_1627_n9724.t2 CLKS.t33 VDDD.t1275 VDDD.t1274 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X192 VSSD.t869 a_1024_n4776.t4 a_958_n4702.t0 VSSD.t868 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X193 a_7243_n1055.t1 a_7068_n1029.t5 a_7422_n1029.t0 VSSD.t833 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X194 a_3235_2717.t0 a_2320_2717.t3 a_2888_2959.t0 VSSD.t362 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X195 a_1627_n9510.t2 a_1452_n9484.t4 a_1806_n9484.t1 VSSD.t68 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X196 SWP[1].t3 a_n6101_n9510.t4 VDDD.t862 VDDD.t861 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X197 a_7248_n9650.t3 a_6333_n10022.t2 a_6901_n10054.t1 VSSD.t744 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X198 a_7230_n663.t1 a_6153_n1029.t2 a_7068_n1029.t2 VDDD.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X199 a_792_n9662.t2 cdac_ctrl_0.x2.X.t18 VSSD.t937 VSSD.t899 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X200 a_n3072_n9484.t1 cdac_ctrl_0.x1.X.t16 VSSD.t31 VSSD.t30 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X201 VDDD.t720 a_1760_n5650.t3 DOUT[2].t3 VDDD.t719 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X202 a_8467_3557.t0 a_7951_3557.t2 a_8372_3557.t0 VSSD.t1005 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X203 VDDD.t526 a_9207_3531.t3 a_9194_3923.t0 VDDD.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X204 a_3181_n1207.t1 CLKS.t34 VSSD.t1102 VSSD.t1101 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X205 SWN[6].t1 a_3559_n9724.t3 VSSD.t620 VSSD.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X206 VSSD.t194 a_n10393_n9484.t8 cdac_ctrl_0.x1.X.t6 VSSD.t193 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X207 a_2451_n5258.t3 a_2325_n5356.t2 a_2047_n5372.t0 VSSD.t1178 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X208 VSSD.t1117 CKO.t5 a_5564_n5074.t0 VSSD.t1116 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X209 VSSD.t789 a_2183_n1599.t3 CF[1].t1 VSSD.t788 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X210 VDDD.t1137 a_n6276_n9650.t4 a_n6101_n9724.t1 VDDD.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X211 a_2451_n5258.t1 a_2364_n5482.t3 a_2047_n5372.t2 VDDD.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X212 a_733_n5258.t2 a_519_n5258.t4 VDDD.t994 VDDD.t993 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X213 a_6080_n4702.t0 a_5564_n5074.t4 a_5985_n4714.t0 VSSD.t604 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X214 a_8711_n9650.t1 a_8265_n10022.t2 a_8615_n9650.t2 VSSD.t69 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X215 a_n454_2691.t0 EN.t11 VDDD.t304 VDDD.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X216 a_n5004_n9662.t3 cdac_ctrl_0.x2.X.t19 VDDD.t1186 VDDD.t1185 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X217 a_n3327_n10022.t1 a_n3493_n10022.t3 VDDD.t592 VDDD.t591 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X218 VDDD.t142 a_1105_n10054.t4 a_995_n10028.t0 VDDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X219 a_2819_n9484.t2 a_2303_n9484.t2 a_2724_n9484.t3 VSSD.t190 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X220 a_n4169_n9724.t0 a_n4344_n9650.t4 a_n3990_n9662.t0 VSSD.t560 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X221 a_n975_3799.t3 a_n1193_3557.t5 VDDD.t689 VDDD.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X222 a_390_n5624.t0 a_n172_n5650.t5 VSSD.t638 VSSD.t637 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X223 a_2364_n5482.t0 CKO.t6 VDDD.t1341 VDDD.t1340 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X224 a_n5922_n9484.t0 CLKS.t35 VSSD.t1100 VSSD.t1078 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X225 VDDD.t83 CF[1].t4 a_1574_n1573.t1 VDDD.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X226 a_7208_2717.t0 a_6018_2717.t2 a_7099_2717.t3 VSSD.t17 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X227 a_887_n9650.t3 a_371_n10022.t2 a_792_n9662.t1 VSSD.t112 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X228 a_115_n5372.t0 a_393_n5356.t2 a_349_n5258.t0 VDDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X229 VDDD.t186 a_n10393_n9484.t9 cdac_ctrl_0.x1.X.t14 VDDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X230 VSSD.t1099 CLKS.t36 a_1149_n9662.t1 VSSD.t1030 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X231 a_7262_3923.t1 a_6185_3557.t2 a_7100_3557.t1 VDDD.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X232 VSSD.t275 EN.t12 a_150_n5624.t0 VSSD.t274 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X233 VSSD.t277 EN.t13 a_4865_3557.t0 VSSD.t276 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X234 a_3083_n5258.t0 a_2325_n5356.t3 a_2520_n5387.t3 VDDD.t1422 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X235 VDDD.t268 a_n10393_n10028.t7 cdac_ctrl_0.x2.X.t1 VDDD.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X236 VDDD.t1181 a_6721_n787.t4 a_6611_n663.t0 VDDD.t1180 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X237 VSSD.t312 a_1024_n4776.t5 DOUT[1].t1 VSSD.t311 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X238 VSSD.t128 a_n2237_n9724.t3 a_n2303_n9650.t0 VSSD.t127 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X239 a_n8033_n9510.t2 CLKS.t37 VDDD.t785 VDDD.t784 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X240 VSSD.t645 CLK.t4 a_2123_n1029.t0 VSSD.t644 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X241 a_n2881_n9650.t0 a_n3327_n10022.t3 a_n2977_n9650.t0 VSSD.t335 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X242 SWN[0].t3 a_n8033_n9724.t3 VDDD.t600 VDDD.t599 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X243 a_4875_n1599.t0 a_4719_n1331.t3 a_5020_n1573.t0 VDDD.t1263 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X244 VDDD.t132 CF[6].t4 a_2303_n9484.t0 VDDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X245 a_6630_2717.t1 a_6184_2717.t2 a_6534_2717.t2 VSSD.t6 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X246 a_8265_n10022.t0 a_8099_n10022.t4 VSSD.t762 VSSD.t24 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 a_n371_n9484.t0 a_n1561_n9484.t2 a_n480_n9484.t1 VSSD.t285 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X248 VDDD.t597 a_855_n1331.t4 a_816_n1457.t1 VDDD.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X249 a_7453_2717.t0 EN.t14 VSSD.t279 VSSD.t278 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X250 a_3088_n1573.t1 a_2874_n1573.t4 VDDD.t641 VDDD.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X251 a_3546_n9118.t0 a_2469_n9484.t2 a_3384_n9484.t0 VDDD.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X252 a_3559_n9724.t0 a_3384_n9650.t4 a_3738_n9662.t0 VSSD.t465 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X253 a_n10393_n10028.t0 COMP_N.t0 VDDD.t287 VDDD.t286 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X254 a_9289_n9484.t0 a_8099_n9484.t3 a_9180_n9484.t2 VSSD.t22 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X255 a_3081_n9662.t0 a_3037_n10054.t4 a_2915_n9650.t0 VSSD.t538 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X256 a_1434_n663.t1 a_357_n1029.t2 a_1272_n1029.t2 VDDD.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X257 a_n5004_n9662.t2 cdac_ctrl_0.x2.X.t20 VSSD.t812 VSSD.t536 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X258 a_2047_n5372.t3 a_2364_n5482.t4 a_2322_n5624.t1 VSSD.t919 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X259 VSSD.t685 a_n6101_n9510.t5 SWP[1].t0 VSSD.t684 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X260 VDDD.t647 a_6753_3799.t4 a_6643_3923.t1 VDDD.t646 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X261 a_6651_n1331.t0 CLK.t5 VSSD.t647 VSSD.t646 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X262 a_n932_2717.t1 a_n976_2959.t4 a_n1098_2717.t1 VSSD.t550 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X263 a_3253_n1207.t0 a_2874_n1573.t5 a_3181_n1207.t0 VSSD.t761 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X264 VSSD.t1003 a_1011_n1599.t4 a_942_n1573.t2 VSSD.t1002 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X265 VSSD.t1165 a_n454_2691.t5 a_n520_2717.t0 VSSD.t1164 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X266 DOUT[8].t0 a_7556_n5650.t5 VSSD.t146 VSSD.t145 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X267 VDDD.t1250 a_4115_n1599.t4 CF[2].t3 VDDD.t1249 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X268 a_3135_n4714.t0 EN.t15 VSSD.t281 VSSD.t280 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X269 a_n3072_n9484.t2 cdac_ctrl_0.x1.X.t17 VDDD.t236 VDDD.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X270 a_4252_2717.t0 a_4086_2717.t2 VSSD.t442 VSSD.t441 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X271 VSSD.t524 CF[8].t5 a_6167_n9484.t0 VSSD.t523 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X272 a_4571_n1029.t0 a_4221_n1029.t3 a_4476_n1029.t0 VDDD.t943 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X273 a_6188_n5080.t1 a_5564_n5074.t5 a_6080_n4702.t1 VDDD.t756 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X274 a_n7854_n9662.t1 CLKS.t38 VSSD.t1098 VSSD.t1026 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X275 a_8626_n5624.t0 a_8247_n5258.t4 a_8554_n5624.t1 VSSD.t43 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X276 VDDD.t749 a_n6101_n9510.t6 SWP[1].t2 VDDD.t748 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X277 a_9175_n1055.t2 a_9000_n1029.t4 a_9354_n1029.t1 VSSD.t1160 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X278 a_2889_3799.t1 a_2671_3557.t5 VSSD.t316 VSSD.t315 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X279 a_2888_2959.t2 a_2670_2717.t5 VDDD.t1167 VDDD.t1166 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X280 a_1466_3923.t1 a_389_3557.t2 a_1304_3557.t0 VDDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X281 VSSD.t655 CF[3].t4 a_n3493_n9484.t0 VSSD.t654 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X282 VDDD.t1004 auto_sampling_0.x23.A.t4 auto_sampling_0.x24.A.t6 VDDD.t1003 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X283 a_4859_n10028.t2 CLKS.t39 VDDD.t614 VDDD.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X284 SWP[5].t1 a_1627_n9510.t3 VSSD.t586 VSSD.t585 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X285 a_9032_3557.t2 a_8117_3557.t2 a_8685_3799.t1 VSSD.t592 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X286 VDDD.t937 a_5343_3531.t4 auto_sampling_0.x5.D.t3 VDDD.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X287 a_4969_n9242.t0 a_4751_n9484.t5 VSSD.t957 VSSD.t678 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X288 a_5985_n4714.t2 SWP[7].t4 VSSD.t980 VSSD.t979 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X289 a_8266_n1441.t3 a_8544_n1457.t2 a_8500_n1573.t0 VDDD.t840 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X290 a_6791_n9118.t2 CLKS.t40 VDDD.t616 VDDD.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X291 VDDD.t541 a_8833_n9242.t4 a_8723_n9118.t1 VDDD.t540 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X292 a_4252_2717.t1 a_4086_2717.t3 VDDD.t511 VDDD.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X293 a_4383_n5258.t0 a_4257_n5356.t2 a_3979_n5372.t2 VSSD.t784 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X294 a_738_2717.t3 a_388_2717.t2 a_643_2717.t3 VDDD.t747 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X295 VSSD.t1097 CLKS.t41 a_n8511_n9484.t1 VSSD.t1071 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X296 a_2216_n4702.t3 a_1866_n5074.t2 a_2121_n4714.t3 VDDD.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X297 a_6791_n9118.t1 a_6167_n9484.t3 a_6683_n9484.t3 VDDD.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X298 a_4603_3557.t2 a_4253_3557.t2 a_4508_3557.t3 VDDD.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X299 a_349_n5258.t1 a_n172_n5650.t6 VDDD.t813 VDDD.t812 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X300 a_1657_2717.t0 EN.t16 VSSD.t283 VSSD.t282 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X301 a_4296_n5482.t1 CKO.t7 VDDD.t1435 VDDD.t1434 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X302 a_2505_n1207.t0 a_2470_n1441.t4 a_2183_n1599.t0 VSSD.t199 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X303 a_3037_n10054.t0 a_2819_n9650.t4 VDDD.t194 VDDD.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X304 SWP[5].t3 a_1627_n9510.t4 VDDD.t1012 VDDD.t1011 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X305 VSSD.t480 a_8752_n4776.t5 a_8686_n4702.t0 VSSD.t479 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X306 VDDD.t618 CLKS.t42 a_4115_n1599.t0 VDDD.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X307 a_7177_n1029.t0 a_5987_n1029.t3 a_7068_n1029.t1 VSSD.t328 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X308 a_8520_n9662.t3 cdac_ctrl_0.x2.X.t21 VDDD.t1038 VDDD.t1037 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X309 a_4256_n5080.t0 EN.t17 VDDD.t894 VDDD.t893 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X310 VDDD.t946 out_latch_0.FINAL.t17 a_9487_n5472.t1 VDDD.t945 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X311 a_846_3083.t2 a_222_2717.t2 a_738_2717.t0 VDDD.t772 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X312 VSSD.t1096 CLKS.t43 a_3081_n9662.t1 VSSD.t1022 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X313 VSSD.t1095 CLKS.t44 a_n783_n9662.t1 VSSD.t1020 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X314 VSSD.t547 a_n784_n1599.t7 out_latch_0.FINAL.t7 VSSD.t546 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X315 a_3590_3557.t0 EN.t18 VSSD.t725 VSSD.t724 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X316 VDDD.t289 a_n8208_n9484.t4 a_n8033_n9510.t0 VDDD.t288 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X317 a_3235_2717.t3 a_2154_2717.t2 a_2888_2959.t3 VDDD.t1375 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X318 a_4711_3923.t1 a_4087_3557.t3 a_4603_3557.t0 VDDD.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X319 a_8697_n1029.t0 a_8653_n787.t4 a_8531_n1029.t0 VSSD.t1143 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X320 a_8108_n4702.t1 a_7662_n5074.t2 a_8012_n4702.t1 VSSD.t577 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X321 a_8728_2717.t1 a_8684_2959.t4 a_8562_2717.t1 VSSD.t981 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X322 VSSD.t649 CLK.t6 a_4055_n1029.t0 VSSD.t648 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X323 a_n1194_2717.t3 a_n1710_2717.t2 a_n1289_2717.t3 VSSD.t398 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X324 a_6820_n4776.t1 a_6645_n4702.t4 a_6999_n4714.t1 VSSD.t343 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X325 VDDD.t1294 a_2781_n4702.t4 a_2956_n4776.t1 VDDD.t1293 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X326 VSSD.t674 CF[2].t4 a_n5425_n10022.t0 VSSD.t673 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X327 VDDD.t692 a_9180_n9650.t4 a_9355_n9724.t0 VDDD.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X328 VDDD.t361 a_4875_n1599.t4 a_4806_n1573.t1 VDDD.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X329 VDDD.t1437 CKO.t8 a_3632_n5074.t1 VDDD.t1436 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X330 a_1000_2717.t1 a_956_2959.t4 a_834_2717.t0 VSSD.t672 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X331 a_887_n9650.t0 a_537_n10022.t2 a_792_n9662.t0 VDDD.t564 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X332 VDDD.t737 a_n2412_n9650.t5 a_n2237_n9724.t1 VDDD.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X333 a_588_n5387.t1 a_432_n5482.t2 a_733_n5258.t1 VDDD.t1094 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X334 VSSD.t562 a_6651_n1331.t3 a_6612_n1457.t0 VSSD.t561 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X335 VDDD.t553 a_1479_3531.t4 auto_sampling_0.x2.D.t3 VDDD.t552 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X336 a_2857_n787.t1 a_2639_n1029.t4 VSSD.t718 VSSD.t717 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X337 a_5911_n5372.t2 a_6189_n5356.t3 a_6145_n5258.t0 VDDD.t1192 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X338 a_3236_3557.t0 a_2321_3557.t2 a_2889_3799.t2 VSSD.t399 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X339 VDDD.t1178 a_432_n5482.t3 a_393_n5356.t0 VDDD.t1177 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X340 a_5730_n5074.t1 a_5564_n5074.t6 VDDD.t758 VDDD.t757 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X341 a_8371_2717.t2 auto_sampling_0.x21.D.t4 VSSD.t118 VSSD.t117 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X342 a_6683_n9650.t2 a_6333_n10022.t3 a_6588_n9662.t1 VDDD.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X343 a_n4813_n9484.t0 a_n5259_n9484.t3 a_n4909_n9484.t1 VSSD.t614 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X344 a_8583_n1331.t0 CLK.t7 VSSD.t651 VSSD.t650 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X345 a_n2977_n9650.t1 a_n3327_n10022.t4 a_n3072_n9662.t0 VDDD.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X346 VSSD.t412 a_2943_n1599.t4 a_2874_n1573.t0 VSSD.t411 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X347 a_8435_n1029.t1 a_8085_n1029.t2 a_8340_n1029.t0 VDDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X348 a_8265_n10022.t1 a_8099_n10022.t5 VDDD.t949 VDDD.t948 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X349 a_388_2717.t0 a_222_2717.t3 VSSD.t347 VSSD.t346 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X350 a_6588_n9484.t0 cdac_ctrl_0.x1.X.t18 VSSD.t228 VSSD.t227 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X351 a_n4909_n9650.t1 a_n5425_n10022.t2 a_n5004_n9662.t0 VSSD.t711 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X352 a_2639_n1029.t1 a_2123_n1029.t2 a_2544_n1029.t2 VSSD.t629 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X353 a_707_n1029.t3 a_357_n1029.t3 a_612_n1029.t3 VDDD.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X354 a_6384_n5387.t0 a_6189_n5356.t4 a_6694_n5624.t0 VSSD.t938 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X355 VDDD.t563 a_3384_n9484.t4 a_3559_n9510.t0 VDDD.t562 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X356 a_2758_n5624.t1 EN.t19 VSSD.t727 VSSD.t726 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X357 a_7068_n1029.t3 a_6153_n1029.t3 a_6721_n787.t2 VSSD.t539 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X358 a_6752_2959.t2 a_6534_2717.t4 VDDD.t16 VDDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X359 a_n3327_n9484.t0 a_n3493_n9484.t2 VSSD.t978 VSSD.t59 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X360 a_4253_3557.t1 a_4087_3557.t4 VDDD.t857 VDDD.t856 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X361 a_n3072_n9662.t3 cdac_ctrl_0.x2.X.t22 VDDD.t1040 VDDD.t1039 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X362 a_n9123_n9484.t1 a_n9289_n9484.t3 VDDD.t126 VDDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X363 a_5342_2691.t0 EN.t20 VDDD.t896 VDDD.t895 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X364 VDDD.t528 a_9207_3531.t4 auto_sampling_0.x11.Q.t3 VDDD.t527 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X365 a_7209_3557.t1 a_6019_3557.t3 a_7100_3557.t0 VSSD.t317 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X366 VDDD.t371 a_n305_n9724.t3 a_n318_n10028.t1 VDDD.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X367 VSSD.t454 a_4296_n5482.t2 a_4257_n5356.t1 VSSD.t453 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X368 VDDD.t803 a_2956_n4776.t3 DOUT[3].t3 VDDD.t802 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X369 a_8543_n663.t0 a_7919_n1029.t2 a_8435_n1029.t2 VDDD.t504 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X370 VSSD.t499 a_9355_n9510.t3 a_9289_n9484.t1 VSSD.t498 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X371 VSSD.t115 a_5342_2691.t3 a_5276_2717.t1 VSSD.t114 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X372 a_6439_2717.t2 auto_sampling_0.x16.D.t4 VDDD.t1343 VDDD.t1342 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X373 a_388_2717.t1 a_222_2717.t4 VDDD.t395 VDDD.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X374 a_2915_n9484.t1 a_2469_n9484.t3 a_2819_n9484.t0 VSSD.t444 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X375 a_815_n663.t0 a_191_n1029.t3 a_707_n1029.t0 VDDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X376 a_n783_n9662.t0 a_n827_n10054.t4 a_n949_n9650.t1 VSSD.t272 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X377 SWP[6].t1 a_3559_n9510.t4 VSSD.t42 VSSD.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X378 a_6901_n9242.t2 a_6683_n9484.t4 VSSD.t841 VSSD.t840 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X379 a_2724_n9484.t1 cdac_ctrl_0.x1.X.t19 VDDD.t238 VDDD.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X380 a_n8665_n10028.t0 a_n9289_n10022.t3 a_n8773_n9650.t0 VDDD.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X381 a_7917_n4714.t1 SWP[9].t4 VDDD.t959 VDDD.t958 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X382 auto_sampling_0.x24.A.t7 auto_sampling_0.x23.A.t5 VSSD.t793 VSSD.t792 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X383 a_8467_3557.t2 a_8117_3557.t3 a_8372_3557.t3 VDDD.t1363 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X384 a_6807_n1599.t1 a_6612_n1457.t2 a_7117_n1207.t0 VSSD.t740 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X385 a_983_n9650.t1 a_537_n10022.t3 a_887_n9650.t1 VSSD.t591 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X386 VSSD.t1094 CLKS.t45 a_8697_n1029.t1 VSSD.t1093 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X387 a_707_n1029.t1 a_191_n1029.t4 a_612_n1029.t2 VSSD.t324 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X388 a_4148_n4702.t2 a_3798_n5074.t2 a_4053_n4714.t3 VDDD.t792 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X389 a_n4801_n9118.t2 CLKS.t46 VDDD.t900 VDDD.t899 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X390 a_n1289_2717.t1 auto_sampling_0.x12.D.t2 VDDD.t506 VDDD.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X391 VDDD.t910 a_n305_n9510.t4 a_n318_n9118.t1 VDDD.t909 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X392 VSSD.t220 a_1447_n1055.t5 CF[9].t0 VSSD.t219 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X393 a_826_n5624.t0 EN.t21 VSSD.t729 VSSD.t728 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X394 a_2890_n4702.t0 a_1700_n5074.t2 a_2781_n4702.t1 VSSD.t1112 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X395 auto_sampling_0.x23.A.t1 auto_sampling_0.x22.A.t4 VSSD.t507 VSSD.t506 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X396 a_2932_2717.t1 a_2888_2959.t5 a_2766_2717.t1 VSSD.t367 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X397 a_n6733_n10028.t0 CLKS.t47 VDDD.t902 VDDD.t901 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X398 DOUT[9].t0 a_8752_n4776.t6 VSSD.t482 VSSD.t481 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X399 auto_sampling_0.x11.D.t3 a_7275_3531.t4 VDDD.t104 VDDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X400 a_4437_n1207.t1 a_4402_n1441.t4 a_4115_n1599.t2 VSSD.t996 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X401 CF[1].t3 a_2183_n1599.t4 VDDD.t1332 VDDD.t1331 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X402 SWP[6].t3 a_3559_n9510.t5 VDDD.t35 VDDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X403 a_6631_3557.t0 a_6185_3557.t3 a_6535_3557.t0 VSSD.t445 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X404 a_n949_n9650.t0 a_n1395_n10022.t3 a_n1045_n9650.t0 VSSD.t590 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X405 a_n2250_n9118.t1 a_n3327_n9484.t2 a_n2412_n9484.t0 VDDD.t1225 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X406 a_7099_2717.t2 a_6018_2717.t3 a_6752_2959.t0 VDDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X407 a_7454_3557.t0 EN.t22 VSSD.t731 VSSD.t730 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X408 a_n6841_n9484.t0 a_n7191_n9484.t2 a_n6936_n9484.t0 VDDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X409 a_846_3083.t0 EN.t23 VDDD.t1415 VDDD.t1414 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X410 a_8575_3923.t1 a_7951_3557.t3 a_8467_3557.t1 VDDD.t1330 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X411 a_2575_2717.t1 auto_sampling_0.x14.D.t4 VSSD.t968 VSSD.t967 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X412 VDDD.t385 a_n10393_n10028.t8 cdac_ctrl_0.x2.X.t2 VDDD.t384 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X413 a_792_n9484.t3 cdac_ctrl_0.x1.X.t20 VDDD.t417 VDDD.t416 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X414 a_6651_n1331.t1 CLK.t8 VDDD.t830 VDDD.t829 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X415 VDDD.t602 a_9355_n9510.t4 a_9342_n9118.t0 VDDD.t601 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X416 a_2639_n1029.t3 a_2289_n1029.t2 a_2544_n1029.t3 VDDD.t1339 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X417 a_n274_3557.t0 EN.t24 VSSD.t1172 VSSD.t1171 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X418 a_4476_n1029.t1 CF[8].t6 VSSD.t526 VSSD.t525 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X419 a_4751_n9484.t2 a_4401_n9484.t2 a_4656_n9484.t1 VDDD.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X420 VDDD.t1258 a_1303_2717.t4 a_1478_2691.t2 VDDD.t1257 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X421 VSSD.t259 COMP_N.t1 a_n10393_n10028.t1 VSSD.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X422 VDDD.t157 a_5342_2691.t4 a_5329_3083.t1 VDDD.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X423 a_7422_n1029.t1 CLKS.t48 VSSD.t1092 VSSD.t1091 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X424 a_n5259_n10022.t0 a_n5425_n10022.t3 VSSD.t425 VSSD.t424 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X425 VSSD.t960 a_1627_n9724.t4 SWN[5].t0 VSSD.t959 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X426 a_537_n10022.t0 a_371_n10022.t3 VSSD.t113 VSSD.t28 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X427 a_1806_n9484.t0 CLKS.t49 VSSD.t1090 VSSD.t1061 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X428 a_3798_n5074.t0 a_3632_n5074.t2 VSSD.t932 VSSD.t931 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X429 a_4253_3557.t0 a_4087_3557.t5 VSSD.t677 VSSD.t676 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X430 a_4366_n5106.t1 a_4148_n4702.t4 VSSD.t302 VSSD.t301 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X431 a_n1395_n9484.t1 a_n1561_n9484.t3 VDDD.t761 VDDD.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X432 cdac_ctrl_0.x2.X.t3 a_n10393_n10028.t9 VDDD.t387 VDDD.t386 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X433 VSSD.t82 CF[1].t5 a_n7357_n10022.t0 VSSD.t81 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X434 VDDD.t1234 a_6807_n1599.t4 a_6738_n1573.t3 VDDD.t1233 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X435 VDDD.t1439 CKO.t9 a_5564_n5074.t1 VDDD.t1438 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X436 a_8118_n5624.t0 a_7556_n5650.t6 VSSD.t148 VSSD.t147 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X437 VSSD.t850 a_7243_n1055.t3 a_7177_n1029.t1 VSSD.t849 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X438 a_2747_n663.t0 a_2123_n1029.t3 a_2639_n1029.t2 VDDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X439 VSSD.t802 a_1627_n9510.t5 a_1561_n9484.t1 VSSD.t801 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X440 a_4789_n787.t2 a_4571_n1029.t4 VSSD.t196 VSSD.t195 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X441 a_5316_n9484.t1 a_4235_n9484.t3 a_4969_n9242.t2 VDDD.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X442 VSSD.t1174 EN.t25 a_6342_n4714.t0 VSSD.t1173 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X443 VDDD.t1149 a_2364_n5482.t5 a_2325_n5356.t1 VDDD.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X444 a_2183_n1599.t1 a_2470_n1441.t5 VDDD.t222 VDDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X445 SWN[2].t1 a_n4169_n9724.t3 VSSD.t686 VSSD.t502 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X446 a_6408_n1029.t3 CF[7].t5 VDDD.t240 VDDD.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X447 SWN[6].t3 a_3559_n9724.t4 VDDD.t771 VDDD.t770 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X448 auto_sampling_0.x16.D.t1 a_5342_2691.t5 VSSD.t153 VSSD.t152 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X449 VDDD.t864 a_n4169_n9724.t4 SWN[2].t3 VDDD.t863 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X450 SWN[4].t3 a_n305_n9724.t4 VDDD.t147 VDDD.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X451 a_n6101_n9510.t1 a_n6276_n9484.t4 a_n5922_n9484.t1 VSSD.t756 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X452 a_2781_n4702.t2 a_1866_n5074.t3 a_2434_n5106.t1 VSSD.t450 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X453 VDDD.t256 a_5316_n9484.t4 a_5491_n9510.t0 VDDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X454 VSSD.t821 CLK.t9 a_n1710_2717.t0 VSSD.t820 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X455 a_389_3557.t0 a_223_3557.t2 VDDD.t974 VDDD.t973 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X456 a_898_n5624.t1 a_519_n5258.t5 a_826_n5624.t1 VSSD.t783 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X457 CF[0].t1 a_251_n1599.t4 VSSD.t911 VSSD.t910 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X458 auto_sampling_0.x2.D.t2 a_1479_3531.t5 VDDD.t555 VDDD.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X459 a_2874_n1573.t2 a_2787_n1331.t3 a_2470_n1441.t0 VDDD.t363 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X460 a_9206_2691.t0 EN.t26 VDDD.t1417 VDDD.t1416 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X461 a_150_n5624.t1 a_115_n5372.t4 a_n172_n5650.t0 VSSD.t628 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X462 a_1658_3557.t0 EN.t27 VSSD.t1176 VSSD.t1175 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X463 VSSD.t1089 CLKS.t50 a_8301_n1207.t1 VSSD.t1088 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X464 VSSD.t356 a_9206_2691.t4 a_9140_2717.t0 VSSD.t355 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X465 a_1303_2717.t2 a_222_2717.t5 a_956_2959.t3 VDDD.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X466 a_2779_3923.t1 a_2155_3557.t3 a_2671_3557.t0 VDDD.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X467 a_8316_n5387.t3 a_8160_n5482.t3 a_8461_n5258.t2 VDDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X468 a_n8511_n9662.t0 a_n8555_n10054.t4 a_n8677_n9650.t1 VSSD.t320 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X469 CF[6].t1 a_7243_n1055.t4 VSSD.t848 VSSD.t847 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X470 a_2121_n4714.t0 SWP[3].t4 VSSD.t45 VSSD.t44 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X471 a_8274_n4714.t1 a_8230_n5106.t4 a_8108_n4702.t0 VSSD.t108 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X472 a_4789_n787.t3 a_4571_n1029.t5 VDDD.t214 VDDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X473 a_1024_n4776.t2 EN.t28 VDDD.t1419 VDDD.t1418 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X474 a_n4344_n9650.t3 a_n5259_n10022.t2 a_n4691_n10054.t1 VSSD.t615 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X475 a_538_n1441.t0 a_816_n1457.t2 a_772_n1573.t0 VDDD.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X476 a_4847_n9484.t0 a_4401_n9484.t3 a_4751_n9484.t3 VSSD.t935 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X477 VDDD.t1014 a_1627_n9510.t6 a_1614_n9118.t1 VDDD.t1013 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X478 a_1105_n10054.t0 a_887_n9650.t4 VDDD.t595 VDDD.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X479 VDDD.t1048 CLK.t10 a_7919_n1029.t1 VDDD.t1047 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X480 VDDD.t165 a_2520_n5387.t4 a_2451_n5258.t0 VDDD.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X481 VDDD.t1050 CLK.t11 a_n1710_2717.t1 VDDD.t1049 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X482 a_4213_n5258.t0 a_3692_n5650.t3 VDDD.t839 VDDD.t838 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X483 CLKS.t12 auto_sampling_0.x24.A.t11 VDDD.t1429 VDDD.t1428 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X484 a_3506_n1573.t3 a_2748_n1457.t2 a_2943_n1599.t3 VDDD.t842 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X485 a_8879_n5258.t3 a_8160_n5482.t4 a_8316_n5387.t2 VSSD.t422 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X486 a_n6733_n9118.t1 CLKS.t51 VDDD.t904 VDDD.t903 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X487 a_6752_2959.t1 a_6534_2717.t5 VSSD.t19 VSSD.t18 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X488 a_8729_3557.t1 a_8685_3799.t4 a_8563_3557.t1 VSSD.t126 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X489 VDDD.t1212 a_1272_n1029.t4 a_1447_n1055.t0 VDDD.t1211 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X490 VDDD.t200 EN.t29 a_2665_n5258.t0 VDDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X491 VDDD.t679 a_5311_n1055.t4 CF[7].t3 VDDD.t678 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X492 a_6683_n9650.t0 a_6167_n10022.t3 a_6588_n9662.t0 VSSD.t201 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X493 VSSD.t1145 a_2520_n5387.t5 a_2451_n5258.t2 VSSD.t1144 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X494 CF[2].t2 a_4115_n1599.t5 VDDD.t1252 VDDD.t1251 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X495 a_3037_n9242.t1 a_2819_n9484.t4 VDDD.t260 VDDD.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X496 a_6439_2717.t1 auto_sampling_0.x16.D.t5 VSSD.t1119 VSSD.t1118 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X497 VSSD.t579 a_3559_n9724.t5 a_3493_n9650.t0 VSSD.t578 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X498 VDDD.t1426 a_6651_n1331.t4 a_6612_n1457.t1 VDDD.t1425 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X499 a_3493_n9650.t1 a_2303_n10022.t2 a_3384_n9650.t1 VSSD.t839 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X500 VDDD.t712 a_5491_n9724.t3 a_5478_n10028.t0 VDDD.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X501 a_1001_3557.t1 a_957_3799.t4 a_835_3557.t0 VSSD.t573 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X502 a_9180_n9650.t0 a_8099_n10022.t6 a_8833_n10054.t0 VDDD.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X503 a_n8046_n10028.t1 a_n9123_n10022.t3 a_n8208_n9650.t1 VDDD.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X504 VDDD.t604 a_3384_n9650.t5 a_3559_n9724.t1 VDDD.t603 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X505 a_8583_n1331.t1 CLK.t12 VDDD.t1052 VDDD.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X506 cdac_ctrl_0.x2.X.t4 a_n10393_n10028.t10 VSSD.t339 VSSD.t170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X507 a_n1140_n9484.t1 cdac_ctrl_0.x1.X.t21 VSSD.t364 VSSD.t363 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X508 a_6153_n1029.t1 a_5987_n1029.t4 VDDD.t368 VDDD.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X509 a_969_n1029.t0 a_925_n787.t4 a_803_n1029.t0 VSSD.t807 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X510 VDDD.t406 a_9206_2691.t5 a_9193_3083.t0 VDDD.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X511 a_n2759_n10054.t0 a_n2977_n9650.t4 VSSD.t35 VSSD.t34 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X512 VDDD.t202 EN.t30 a_1760_n5650.t0 VDDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X513 auto_sampling_0.x12.D.t1 auto_sampling_0.x11.Q.t4 VDDD.t324 VDDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X514 a_8372_3557.t1 auto_sampling_0.x11.D.t4 VSSD.t332 VSSD.t331 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X515 a_n8033_n9724.t1 a_n8208_n9650.t4 a_n7854_n9662.t0 VSSD.t531 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X516 a_8723_n10028.t2 CLKS.t52 VDDD.t906 VDDD.t905 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X517 DOUT[1].t3 a_1024_n4776.t6 VDDD.t347 VDDD.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X518 a_n4344_n9484.t3 a_n5425_n9484.t2 a_n4691_n9242.t3 VDDD.t1157 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X519 a_2670_2717.t2 a_2154_2717.t3 a_2575_2717.t3 VSSD.t395 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X520 a_8543_n663.t2 CLKS.t53 VDDD.t908 VDDD.t907 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X521 VSSD.t1153 SWP[2].t4 a_3083_n5258.t2 VSSD.t1152 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X522 VDDD.t674 a_n976_2959.t5 a_n1086_3083.t2 VDDD.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X523 a_389_3557.t1 a_223_3557.t3 VSSD.t774 VSSD.t773 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X524 VDDD.t204 EN.t31 a_733_n5258.t0 VDDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X525 a_3410_2691.t2 EN.t32 VDDD.t206 VDDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X526 a_9354_n1029.t0 CLKS.t54 VSSD.t1087 VSSD.t1086 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X527 VDDD.t159 a_5342_2691.t6 auto_sampling_0.x16.D.t3 VDDD.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X528 a_n519_3557.t0 a_n1709_3557.t4 a_n628_3557.t2 VSSD.t832 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X529 a_3738_n9484.t1 CLKS.t55 VSSD.t1085 VSSD.t1058 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X530 a_n8033_n9724.t2 CLKS.t56 VDDD.t499 VDDD.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X531 auto_sampling_0.x24.A.t0 auto_sampling_0.x23.A.t6 VSSD.t120 VSSD.t119 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X532 a_6298_n5106.t1 a_6080_n4702.t4 VSSD.t488 VSSD.t487 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X533 a_n4801_n9118.t1 a_n5425_n9484.t3 a_n4909_n9484.t3 VDDD.t1158 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X534 VDDD.t854 CF[2].t5 a_n5425_n10022.t1 VDDD.t853 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X535 a_n4235_n9650.t1 a_n5425_n10022.t4 a_n4344_n9650.t0 VSSD.t426 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X536 VSSD.t187 EN.t33 a_1000_2717.t0 VSSD.t186 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X537 VSSD.t76 a_n4169_n9724.t5 SWN[2].t0 VSSD.t75 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X538 a_2735_n1029.t0 a_2289_n1029.t3 a_2639_n1029.t0 VSSD.t556 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X539 VSSD.t545 CF[2].t6 a_3506_n1573.t1 VSSD.t544 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X540 VSSD.t189 EN.t34 a_8274_n4714.t0 VSSD.t188 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X541 a_7261_3083.t0 a_6184_2717.t3 a_7099_2717.t0 VDDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X542 auto_sampling_0.x21.Q.t1 a_9206_2691.t6 VSSD.t358 VSSD.t357 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X543 a_4115_n1599.t1 a_4402_n1441.t5 VDDD.t1296 VDDD.t1295 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X544 VSSD.t748 a_5343_3531.t5 a_5277_3557.t1 VSSD.t747 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X545 a_n1045_n9650.t3 a_n1561_n10022.t2 a_n1140_n9662.t1 VSSD.t284 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X546 a_8739_n1599.t0 a_8583_n1331.t5 a_8884_n1573.t0 VDDD.t1328 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X547 a_n2759_n10054.t1 a_n2977_n9650.t5 VDDD.t28 VDDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X548 VSSD.t138 a_n305_n9724.t5 a_n371_n9650.t1 VSSD.t137 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X549 a_n784_n1599.t2 CF[0].t4 VSSD.t376 VSSD.t375 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X550 a_8575_3923.t0 EN.t35 VDDD.t777 VDDD.t776 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X551 a_n784_n1599.t3 CF[0].t5 VSSD.t378 VSSD.t377 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X552 a_7410_n9118.t1 a_6333_n9484.t3 a_7248_n9484.t3 VDDD.t934 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X553 VSSD.t107 a_9355_n9724.t4 SWN[9].t1 VSSD.t106 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X554 a_2874_n1573.t3 a_2748_n1457.t3 a_2470_n1441.t2 VSSD.t659 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X555 VSSD.t549 a_n784_n1599.t8 out_latch_0.FINAL.t6 VSSD.t548 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X556 a_n6276_n9650.t2 a_n7357_n10022.t4 a_n6623_n10054.t3 VDDD.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X557 a_3384_n9650.t2 a_2469_n10022.t3 a_3037_n10054.t3 VSSD.t589 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X558 a_2289_n1029.t0 a_2123_n1029.t4 VSSD.t37 VSSD.t36 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X559 a_2933_3557.t1 a_2889_3799.t4 a_2767_3557.t0 VSSD.t319 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X560 CF[5].t1 a_9175_n1055.t5 VSSD.t291 VSSD.t290 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X561 a_803_n1029.t1 a_357_n1029.t4 a_707_n1029.t2 VSSD.t865 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X562 a_n937_n10028.t0 a_n1561_n10022.t3 a_n1045_n9650.t2 VDDD.t307 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X563 a_4053_n4714.t1 SWP[5].t4 VSSD.t634 VSSD.t633 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X564 VSSD.t1189 CKO.t10 a_1700_n5074.t0 VSSD.t1188 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X565 a_4859_n9118.t1 CLKS.t57 VDDD.t501 VDDD.t500 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X566 a_2956_n4776.t0 EN.t36 VDDD.t779 VDDD.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X567 a_2469_n9484.t1 a_2303_n9484.t3 VDDD.t210 VDDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X568 a_n6276_n9650.t0 a_n7191_n10022.t2 a_n6623_n10054.t2 VSSD.t889 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X569 VDDD.t130 auto_sampling_0.x23.A.t7 auto_sampling_0.x24.A.t1 VDDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X570 VDDD.t815 a_n172_n5650.t7 DOUT[0].t2 VDDD.t814 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X571 a_9342_n10028.t1 a_8265_n10022.t3 a_9180_n9650.t3 VDDD.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X572 a_n8208_n9650.t2 a_n9289_n10022.t4 a_n8555_n10054.t3 VDDD.t921 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X573 a_8461_n5258.t1 a_8247_n5258.t5 VDDD.t39 VDDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X574 a_2576_3557.t1 auto_sampling_0.x2.D.t4 VSSD.t786 VSSD.t785 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X575 VDDD.t561 a_6752_2959.t4 a_6642_3083.t2 VDDD.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X576 VSSD.t600 a_n6101_n9510.t7 a_n6167_n9484.t1 VSSD.t286 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X577 a_7423_n9724.t2 CLKS.t58 VDDD.t503 VDDD.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X578 VDDD.t1106 a_5136_n1029.t4 a_5311_n1055.t0 VDDD.t1105 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X579 VDDD.t322 a_9175_n1055.t6 CF[5].t2 VDDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X580 a_1304_3557.t2 a_223_3557.t4 a_957_3799.t2 VDDD.t1456 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X581 a_2747_n663.t2 CLKS.t59 VDDD.t1301 VDDD.t1300 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X582 a_6145_n5258.t1 a_5624_n5650.t3 VDDD.t306 VDDD.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X583 a_5438_n1573.t1 a_4680_n1457.t3 a_4875_n1599.t3 VDDD.t985 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X584 VDDD.t49 a_1478_2691.t3 auto_sampling_0.x14.D.t2 VDDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X585 VDDD.t620 auto_sampling_0.x22.A.t5 auto_sampling_0.x23.A.t3 VDDD.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X586 VDDD.t536 CF[5].t6 a_371_n10022.t1 VDDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X587 a_7423_n9510.t1 a_7248_n9484.t4 a_7602_n9484.t0 VSSD.t584 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X588 VSSD.t606 a_4452_n5387.t5 a_4383_n5258.t1 VSSD.t605 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X589 a_4476_n1029.t2 CF[8].t7 VDDD.t643 VDDD.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X590 VDDD.t521 a_7556_n5650.t7 DOUT[8].t3 VDDD.t520 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X591 a_n9123_n10022.t0 a_n9289_n10022.t5 VDDD.t923 VDDD.t922 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X592 a_1465_3083.t1 a_388_2717.t3 a_1303_2717.t0 VDDD.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X593 a_1760_n5650.t1 a_2047_n5372.t4 VDDD.t1194 VDDD.t1193 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X594 auto_sampling_0.x15.D.t1 a_3410_2691.t4 VSSD.t809 VSSD.t808 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X595 a_n480_n9484.t2 a_n1395_n9484.t2 a_n827_n9242.t3 VSSD.t775 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X596 a_8247_n5258.t2 a_8121_n5356.t3 a_7843_n5372.t1 VSSD.t141 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X597 a_4713_n4702.t1 a_3632_n5074.t3 a_4366_n5106.t0 VDDD.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X598 VSSD.t383 a_7979_n1599.t3 CF[4].t0 VSSD.t382 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X599 VSSD.t1183 auto_sampling_0.x24.A.t12 CLKS.t13 VSSD.t1182 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X600 VSSD.t622 EN.t37 a_n931_3557.t0 VSSD.t621 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X601 a_n6936_n9662.t2 cdac_ctrl_0.x2.X.t23 VDDD.t1042 VDDD.t1041 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X602 a_6534_2717.t0 a_6018_2717.t4 a_6439_2717.t0 VSSD.t321 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X603 a_1011_n1599.t2 a_855_n1331.t5 a_1156_n1573.t0 VDDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X604 VDDD.t961 a_5168_3557.t4 a_5343_3531.t1 VDDD.t960 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X605 a_1149_n9484.t0 a_1105_n9242.t5 a_983_n9484.t1 VSSD.t133 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X606 a_2779_3923.t0 EN.t38 VDDD.t781 VDDD.t780 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X607 VSSD.t542 COMP_P.t0 a_n10393_n9484.t0 VSSD.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X608 a_2364_n5482.t1 CKO.t11 VSSD.t1156 VSSD.t1155 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X609 VDDD.t408 a_9206_2691.t7 auto_sampling_0.x21.Q.t2 VDDD.t407 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X610 a_8615_n9484.t2 a_8099_n9484.t4 a_8520_n9484.t1 VSSD.t23 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X611 DOUT[3].t2 a_2956_n4776.t4 VDDD.t413 VDDD.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X612 a_4401_n10022.t0 a_4235_n10022.t4 VSSD.t437 VSSD.t436 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X613 a_2745_n1207.t1 a_2183_n1599.t5 VSSD.t971 VSSD.t970 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X614 a_n6276_n9484.t1 a_n7357_n9484.t4 a_n6623_n9242.t0 VDDD.t805 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X615 auto_sampling_0.x5.D.t1 a_5343_3531.t6 VSSD.t750 VSSD.t749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X616 VSSD.t1179 a_1627_n9510.t7 SWP[5].t0 VSSD.t959 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X617 a_8160_n5482.t1 CKO.t12 VDDD.t1391 VDDD.t1390 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X618 a_2470_n1441.t1 a_2787_n1331.t4 a_2745_n1207.t0 VSSD.t794 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X619 VDDD.t1 CF[4].t6 a_7370_n1573.t2 VDDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X620 a_4602_2717.t2 a_4252_2717.t2 a_4507_2717.t1 VDDD.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X621 a_5425_n9484.t0 a_4235_n9484.t4 a_5316_n9484.t0 VSSD.t149 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X622 a_957_3799.t0 a_739_3557.t4 VDDD.t331 VDDD.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X623 VDDD.t291 a_6820_n4776.t3 a_6807_n5080.t0 VDDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X624 VDDD.t1054 CLK.t13 a_191_n1029.t1 VDDD.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X625 auto_sampling_0.x7.Q.t1 a_n453_3531.t4 VSSD.t894 VSSD.t893 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X626 VSSD.t222 a_9207_3531.t5 a_9141_3557.t1 VSSD.t221 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X627 VDDD.t666 COMP_P.t1 a_n10393_n9484.t1 VDDD.t665 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X628 VDDD.t746 a_n2759_n10054.t5 a_n2869_n10028.t1 VDDD.t745 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X629 VDDD.t1008 a_9355_n9724.t5 SWN[9].t2 VDDD.t1007 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X630 a_4969_n10054.t3 a_4751_n9650.t4 VSSD.t679 VSSD.t678 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X631 VDDD.t892 a_4366_n5106.t4 a_4256_n5080.t2 VDDD.t891 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X632 a_3411_3531.t0 EN.t39 VDDD.t783 VDDD.t782 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X633 VSSD.t263 a_6820_n4776.t4 DOUT[7].t1 VSSD.t262 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X634 VSSD.t657 CF[3].t5 a_5438_n1573.t2 VSSD.t656 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X635 SWP[2].t1 a_n4169_n9510.t4 VSSD.t503 VSSD.t502 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X636 DOUT[4].t1 a_3692_n5650.t4 VSSD.t662 VSSD.t661 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X637 VSSD.t8 a_n8033_n9724.t4 a_n8099_n9650.t1 VSSD.t7 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X638 VDDD.t1424 a_1627_n9510.t8 SWP[5].t2 VDDD.t1423 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X639 VSSD.t624 EN.t40 a_7878_n5624.t0 VSSD.t623 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X640 auto_sampling_0.x21.D.t3 a_7274_2691.t4 VDDD.t53 VDDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X641 a_n8868_n9484.t2 cdac_ctrl_0.x1.X.t22 VSSD.t366 VSSD.t365 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X642 a_n2977_n9650.t3 a_n3493_n10022.t4 a_n3072_n9662.t1 VSSD.t58 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X643 a_4710_3083.t1 a_4086_2717.t4 a_4602_2717.t1 VDDD.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X644 VSSD.t124 CF[6].t5 a_2303_n9484.t1 VSSD.t123 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X645 a_2324_n5080.t1 a_1700_n5074.t3 a_2216_n4702.t0 VDDD.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X646 a_813_n1207.t1 a_251_n1599.t5 VSSD.t913 VSSD.t912 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X647 VDDD.t285 CF[9].t5 a_8099_n9484.t1 VDDD.t284 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X648 out_latch_0.FINAL.t5 a_n784_n1599.t9 VSSD.t852 VSSD.t851 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 VDDD.t687 a_n4691_n10054.t4 a_n4801_n10028.t0 VDDD.t686 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X650 a_519_n5258.t2 a_432_n5482.t4 a_115_n5372.t2 VDDD.t1179 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X651 a_8884_n1573.t1 a_8670_n1573.t4 VDDD.t329 VDDD.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X652 a_5311_n1055.t1 a_5136_n1029.t5 a_5490_n1029.t0 VSSD.t872 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X653 a_9342_n9118.t1 a_8265_n9484.t2 a_9180_n9484.t3 VDDD.t858 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X654 a_9355_n9724.t1 a_9180_n9650.t5 a_9534_n9662.t0 VSSD.t519 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X655 a_n6167_n9484.t0 a_n7357_n9484.t5 a_n6276_n9484.t0 VSSD.t520 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X656 a_8685_3799.t3 a_8467_3557.t4 VDDD.t421 VDDD.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X657 a_6753_3799.t0 a_6535_3557.t5 VSSD.t360 VSSD.t359 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X658 VDDD.t1368 a_3379_n1055.t6 a_3366_n663.t0 VDDD.t1367 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X659 VSSD.t1084 CLKS.t60 a_573_n1207.t1 VSSD.t1083 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X660 SWP[2].t3 a_n4169_n9510.t5 VDDD.t1336 VDDD.t1335 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X661 VDDD.t1431 auto_sampling_0.x24.A.t13 CLKS.t14 VDDD.t1430 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X662 VSSD.t1158 CKO.t13 a_n232_n5074.t0 VSSD.t1157 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X663 a_4402_n1441.t2 a_4680_n1457.t4 a_4636_n1573.t0 VDDD.t986 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X664 a_7843_n5372.t3 a_8160_n5482.t5 a_8118_n5624.t1 VSSD.t423 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X665 a_546_n4714.t1 a_502_n5106.t5 a_380_n4702.t1 VSSD.t888 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X666 VDDD.t1240 a_9000_n1029.t5 a_9175_n1055.t0 VDDD.t1239 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X667 VSSD.t261 COMP_N.t2 a_n10393_n10028.t2 VSSD.t260 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X668 a_5168_3557.t0 a_4087_3557.t6 a_4821_3799.t0 VDDD.t1348 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X669 a_6611_n663.t2 CLKS.t61 VDDD.t1303 VDDD.t1302 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X670 a_6503_n1029.t2 a_5987_n1029.t5 a_6408_n1029.t0 VSSD.t329 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X671 VDDD.t1246 a_n8033_n9510.t4 a_n8046_n9118.t1 VDDD.t1245 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X672 a_3798_n5074.t1 a_3632_n5074.t4 VDDD.t426 VDDD.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X673 a_3384_n9650.t0 a_2303_n10022.t3 a_3037_n10054.t2 VDDD.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X674 a_6622_n5624.t0 EN.t41 VSSD.t267 VSSD.t266 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X675 a_n976_2959.t1 a_n1194_2717.t4 VSSD.t459 VSSD.t458 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X676 VDDD.t112 SWP[4].t5 a_5015_n5258.t1 VDDD.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X677 a_432_n5482.t1 CKO.t14 VDDD.t1393 VDDD.t1392 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X678 a_5316_n9484.t3 a_4401_n9484.t4 a_4969_n9242.t3 VSSD.t534 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X679 a_3313_n1029.t1 a_2123_n1029.t5 a_3204_n1029.t2 VSSD.t38 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X680 a_2671_3557.t1 a_2155_3557.t4 a_2576_3557.t0 VSSD.t535 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X681 VDDD.t1130 a_n453_3531.t5 a_n466_3923.t1 VDDD.t1129 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X682 a_4452_n5387.t0 a_4257_n5356.t3 a_4762_n5624.t0 VSSD.t704 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X683 DOUT[8].t2 a_7556_n5650.t8 VDDD.t523 VDDD.t522 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X684 VDDD.t988 a_3411_3531.t4 a_3398_3923.t0 VDDD.t987 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X685 a_6791_n10028.t2 CLKS.t62 VDDD.t1305 VDDD.t1304 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X686 a_7099_2717.t1 a_6184_2717.t4 a_6752_2959.t3 VSSD.t57 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X687 a_n318_n10028.t0 a_n1395_n10022.t4 a_n480_n9650.t1 VDDD.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X688 a_n8208_n9484.t3 a_n9123_n9484.t2 a_n8555_n9242.t1 VSSD.t787 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X689 a_1151_n5258.t1 a_393_n5356.t3 a_588_n5387.t3 VDDD.t208 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X690 CLKSB.t1 CLKS.t63 VDDD.t1307 VDDD.t1306 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X691 SWN[8].t1 a_7423_n9724.t3 VSSD.t1150 VSSD.t733 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X692 a_n1098_2717.t0 a_n1544_2717.t2 a_n1194_2717.t1 VSSD.t916 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X693 SWN[4].t1 a_n305_n9724.t6 VSSD.t140 VSSD.t139 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X694 a_6588_n9484.t1 cdac_ctrl_0.x1.X.t23 VDDD.t98 VDDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X695 auto_sampling_0.x14.D.t3 a_1478_2691.t4 VDDD.t51 VDDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X696 VSSD.t269 EN.t42 a_1001_3557.t0 VSSD.t268 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X697 cdac_ctrl_0.x1.X.t5 a_n10393_n9484.t10 VSSD.t171 VSSD.t170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X698 a_n6101_n9510.t0 CLKS.t64 VDDD.t493 VDDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X699 a_n629_2717.t1 a_n1544_2717.t3 a_n976_2959.t0 VSSD.t379 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X700 VSSD.t231 CF[7].t6 a_4235_n10022.t0 VSSD.t229 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X701 VSSD.t1082 CLKS.t65 a_6945_n9484.t1 VSSD.t1045 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X702 VDDD.t976 CF[0].t6 a_n9289_n9484.t1 VDDD.t975 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X703 a_4859_n10028.t0 a_4235_n10022.t5 a_4751_n9650.t0 VDDD.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X704 a_1412_2717.t1 a_222_2717.t6 a_1303_2717.t3 VSSD.t669 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X705 auto_sampling_0.x11.Q.t1 a_9207_3531.t6 VSSD.t224 VSSD.t223 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X706 a_8466_2717.t2 a_8116_2717.t3 a_8371_2717.t1 VDDD.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X707 a_4296_n5482.t0 CKO.t15 VSSD.t72 VSSD.t71 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X708 a_n305_n9724.t0 a_n480_n9650.t4 a_n126_n9662.t0 VSSD.t273 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X709 a_995_n10028.t1 a_371_n10022.t4 a_887_n9650.t2 VDDD.t750 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X710 a_6333_n10022.t0 a_6167_n10022.t4 VSSD.t203 VSSD.t202 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X711 a_4821_3799.t3 a_4603_3557.t4 VDDD.t704 VDDD.t703 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X712 a_1156_n1573.t1 a_942_n1573.t5 VDDD.t880 VDDD.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X713 a_8301_n1207.t0 a_8266_n1441.t4 a_7979_n1599.t0 VSSD.t1161 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X714 a_1627_n9724.t0 a_1452_n9650.t4 a_1806_n9662.t0 VSSD.t68 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X715 a_6807_n5080.t1 a_5730_n5074.t3 a_6645_n4702.t3 VDDD.t1400 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X716 a_7357_n9484.t1 a_6167_n9484.t4 a_7248_n9484.t0 VSSD.t200 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X717 a_n3072_n9662.t2 cdac_ctrl_0.x2.X.t24 VSSD.t813 VSSD.t30 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X718 a_6791_n10028.t0 a_6167_n10022.t5 a_6683_n9650.t1 VDDD.t1173 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X719 cdac_ctrl_0.x1.X.t13 a_n10393_n9484.t11 VDDD.t188 VDDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X720 DOUT[7].t0 a_6820_n4776.t5 VSSD.t265 VSSD.t264 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X721 a_7275_3531.t0 EN.t43 VDDD.t293 VDDD.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X722 VSSD.t1113 a_n4169_n9510.t6 SWP[2].t0 VSSD.t75 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X723 a_2434_n5106.t3 a_2216_n4702.t4 VDDD.t1016 VDDD.t1015 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X724 cdac_ctrl_0.x2.X.t5 a_n10393_n10028.t11 VDDD.t389 VDDD.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X725 a_n318_n9118.t0 a_n1395_n9484.t3 a_n480_n9484.t0 VDDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X726 a_4719_n1331.t0 CLK.t14 VSSD.t823 VSSD.t822 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X727 VDDD.t77 a_n4169_n9724.t6 a_n4182_n10028.t1 VDDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X728 a_8574_3083.t1 a_7950_2717.t3 a_8466_2717.t0 VDDD.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X729 a_6901_n10054.t2 a_6683_n9650.t4 VSSD.t941 VSSD.t840 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X730 a_9661_n4742.t1 CLKS.t66 VSSD.t1081 VSSD.t1080 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X731 a_644_3557.t3 auto_sampling_0.x7.Q.t5 VDDD.t730 VDDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X732 a_2724_n9484.t0 cdac_ctrl_0.x1.X.t24 VSSD.t98 VSSD.t97 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X733 DOUT[6].t1 a_5624_n5650.t4 VSSD.t903 VSSD.t902 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X734 VDDD.t1262 a_2183_n1599.t6 CF[1].t2 VDDD.t1261 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X735 VSSD.t1185 auto_sampling_0.x24.A.t14 CLKS.t15 VSSD.t1184 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X736 a_n4647_n9484.t0 a_n4691_n9242.t5 a_n4813_n9484.t1 VSSD.t464 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X737 a_n453_3531.t0 EN.t44 VDDD.t295 VDDD.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X738 a_8877_n9484.t0 a_8833_n9242.t5 a_8711_n9484.t1 VSSD.t452 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X739 a_n1140_n9484.t2 cdac_ctrl_0.x1.X.t25 VDDD.t100 VDDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X740 a_4256_n5080.t1 a_3632_n5074.t5 a_4148_n4702.t0 VDDD.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X741 a_3204_n1029.t1 a_2289_n1029.t4 a_2857_n787.t0 VSSD.t557 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X742 a_n5922_n9662.t1 CLKS.t67 VSSD.t1079 VSSD.t1078 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X743 a_2819_n9484.t1 a_2469_n9484.t4 a_2724_n9484.t2 VDDD.t790 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X744 a_6694_n5624.t1 a_6315_n5258.t4 a_6622_n5624.t1 VSSD.t767 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X745 VSSD.t1140 a_9355_n9510.t5 SWP[9].t1 VSSD.t106 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X746 VDDD.t1350 a_n4169_n9510.t7 SWP[2].t2 VDDD.t1349 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X747 VSSD.t340 a_n10393_n10028.t12 cdac_ctrl_0.x2.X.t6 VSSD.t172 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X748 VDDD.t696 a_n4344_n9650.t5 a_n4169_n9724.t1 VDDD.t695 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X749 a_n8099_n9484.t0 a_n9289_n9484.t4 a_n8208_n9484.t1 VSSD.t630 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X750 VDDD.t391 a_n10393_n10028.t13 cdac_ctrl_0.x2.X.t7 VDDD.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X751 VSSD.t934 a_432_n5482.t5 a_393_n5356.t1 VSSD.t933 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X752 a_n453_3531.t1 a_n628_3557.t4 a_n274_3557.t1 VSSD.t1147 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X753 a_n1395_n10022.t0 a_n1561_n10022.t4 VDDD.t309 VDDD.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X754 VSSD.t567 a_5491_n9510.t5 a_5425_n9484.t1 VSSD.t566 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X755 a_n8773_n9650.t3 a_n9123_n10022.t4 a_n8868_n9662.t1 VDDD.t998 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X756 a_n10393_n10028.t3 COMP_N.t3 VSSD.t419 VSSD.t418 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X757 CLKS.t7 auto_sampling_0.x24.A.t15 VDDD.t470 VDDD.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X758 a_502_n5106.t2 a_284_n4702.t4 VDDD.t878 VDDD.t877 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X759 a_3037_n9242.t0 a_2819_n9484.t5 VSSD.t607 VSSD.t178 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X760 a_5298_n663.t1 a_4221_n1029.t4 a_5136_n1029.t0 VDDD.t944 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X761 a_6334_n1441.t1 a_6612_n1457.t3 a_6568_n1573.t0 VDDD.t1095 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X762 VDDD.t612 a_6901_n9242.t4 a_6791_n9118.t0 VDDD.t611 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X763 a_n480_n9650.t2 a_n1561_n10022.t5 a_n827_n10054.t1 VDDD.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X764 VSSD.t1077 CLKS.t68 a_4833_n1029.t1 VSSD.t1076 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X765 VSSD.t1075 CLKS.t69 a_n6579_n9484.t1 VSSD.t1041 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X766 VDDD.t1370 a_9355_n9510.t6 SWP[9].t3 VDDD.t1369 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X767 auto_sampling_0.x3.D.t0 a_3411_3531.t5 VSSD.t782 VSSD.t781 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X768 VDDD.t3 CF[4].t7 a_n1561_n9484.t1 VDDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X769 VDDD.t242 CF[7].t7 a_4235_n10022.t1 VDDD.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X770 a_8435_n1029.t3 a_7919_n1029.t3 a_8340_n1029.t3 VSSD.t508 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X771 VDDD.t184 a_n305_n9724.t7 SWN[4].t2 VDDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X772 a_2670_2717.t0 a_2320_2717.t4 a_2575_2717.t0 VDDD.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X773 SWN[3].t1 a_n2237_n9724.t4 VSSD.t129 VSSD.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X774 a_6535_3557.t2 a_6019_3557.t4 a_6440_3557.t0 VSSD.t318 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X775 a_8554_n5624.t0 EN.t45 VSSD.t271 VSSD.t270 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X776 VDDD.t106 a_7275_3531.t5 a_7262_3923.t0 VDDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X777 VDDD.t832 SWP[6].t4 a_6947_n5258.t2 VDDD.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X778 a_8116_2717.t0 a_7950_2717.t4 VSSD.t236 VSSD.t235 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X779 a_n9123_n9484.t0 a_n9289_n9484.t5 VSSD.t632 VSSD.t631 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X780 VSSD.t533 a_6820_n4776.t6 a_6754_n4702.t1 VSSD.t532 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X781 VDDD.t116 CLKS.t70 a_2183_n1599.t2 VDDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X782 a_7248_n9484.t2 a_6333_n9484.t4 a_6901_n9242.t1 VSSD.t744 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X783 a_5245_n1029.t1 a_4055_n1029.t2 a_5136_n1029.t3 VSSD.t478 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X784 VDDD.t714 a_5491_n9724.t4 SWN[7].t3 VDDD.t713 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X785 a_2324_n5080.t0 EN.t46 VDDD.t297 VDDD.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X786 a_1479_3531.t0 EN.t47 VDDD.t1319 VDDD.t1318 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X787 SWN[1].t3 a_n6101_n9724.t5 VDDD.t318 VDDD.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X788 VDDD.t577 a_8752_n4776.t7 DOUT[9].t3 VDDD.t576 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X789 VDDD.t1458 a_n6276_n9484.t5 a_n6101_n9510.t2 VDDD.t1457 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X790 a_8711_n9484.t0 a_8265_n9484.t3 a_8615_n9484.t0 VSSD.t69 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X791 a_2778_3083.t2 a_2154_2717.t4 a_2670_2717.t3 VDDD.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X792 SWN[9].t0 a_9355_n9724.t6 VSSD.t799 VSSD.t798 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X793 a_8520_n9484.t3 cdac_ctrl_0.x1.X.t26 VDDD.t1451 VDDD.t1450 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X794 a_519_n5258.t1 a_393_n5356.t4 a_115_n5372.t1 VSSD.t745 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X795 VSSD.t915 a_251_n1599.t6 CF[0].t0 VSSD.t914 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X796 a_6765_n1029.t0 a_6721_n787.t5 a_6599_n1029.t0 VSSD.t1154 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X797 VDDD.t258 a_4789_n787.t4 a_4679_n663.t1 VDDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X798 a_5276_2717.t0 a_4086_2717.t5 a_5167_2717.t1 VSSD.t416 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X799 a_6176_n4702.t1 a_5730_n5074.t4 a_6080_n4702.t3 VSSD.t1166 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X800 a_8116_2717.t1 a_7950_2717.t5 VDDD.t250 VDDD.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X801 auto_sampling_0.x22.A.t3 a_n454_2691.t6 VDDD.t196 VDDD.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X802 VSSD.t527 CF[8].t8 a_6167_n10022.t0 VSSD.t523 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X803 VSSD.t1074 CLKS.t71 a_8877_n9484.t1 VSSD.t1037 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X804 a_n66_n5074.t0 a_n232_n5074.t2 VSSD.t65 VSSD.t64 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X805 VSSD.t825 CLK.t15 a_6018_2717.t0 VSSD.t824 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X806 a_5330_3923.t0 a_4253_3557.t3 a_5168_3557.t2 VDDD.t607 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X807 a_887_n9484.t1 a_371_n9484.t3 a_792_n9484.t0 VSSD.t112 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X808 a_n4691_n9242.t1 a_n4909_n9484.t4 VDDD.t1074 VDDD.t1073 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X809 VDDD.t1321 EN.t48 a_6529_n5258.t0 VDDD.t1320 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X810 VSSD.t854 a_n784_n1599.t10 out_latch_0.FINAL.t4 VSSD.t853 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X811 VSSD.t846 a_7243_n1055.t5 CF[6].t0 VSSD.t845 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X812 VDDD.t954 a_849_n4702.t4 a_1024_n4776.t1 VDDD.t953 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X813 a_4698_2717.t0 a_4252_2717.t3 a_4602_2717.t3 VSSD.t771 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X814 VSSD.t987 CF[3].t6 a_n3493_n10022.t0 VSSD.t654 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X815 VDDD.t468 a_2943_n1599.t5 a_2874_n1573.t1 VDDD.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X816 out_latch_0.FINAL.t3 a_n784_n1599.t11 VSSD.t856 VSSD.t855 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X817 VDDD.t67 CKO.t16 a_1700_n5074.t1 VDDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X818 a_8739_n5080.t1 a_7662_n5074.t3 a_8577_n4702.t2 VDDD.t951 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X819 VSSD.t233 a_4719_n1331.t4 a_4680_n1457.t0 VSSD.t232 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X820 a_n2058_n9484.t1 CLKS.t72 VSSD.t1073 VSSD.t1035 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X821 a_n8046_n9118.t0 a_n9123_n9484.t3 a_n8208_n9484.t2 VDDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X822 a_925_n787.t1 a_707_n1029.t4 VSSD.t403 VSSD.t402 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X823 a_3979_n5372.t1 a_4257_n5356.t4 a_4213_n5258.t1 VDDD.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X824 a_n2881_n9484.t0 a_n3327_n9484.t3 a_n2977_n9484.t1 VSSD.t335 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X825 a_1105_n9242.t2 a_887_n9484.t4 VDDD.t1067 VDDD.t1066 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X826 VSSD.t999 EN.t49 a_4014_n5624.t0 VSSD.t998 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X827 VSSD.t1072 CLKS.t73 a_n8511_n9662.t1 VSSD.t1071 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X828 VDDD.t1113 CLK.t16 a_6018_2717.t1 VDDD.t1112 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X829 VSSD.t877 CLK.t17 a_7919_n1029.t0 VSSD.t876 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X830 VSSD.t879 CLK.t18 a_191_n1029.t0 VSSD.t878 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X831 a_4656_n9484.t2 cdac_ctrl_0.x1.X.t27 VSSD.t1192 VSSD.t570 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X832 a_n6579_n9484.t0 a_n6623_n9242.t5 a_n6745_n9484.t0 VSSD.t151 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X833 VDDD.t1160 a_1452_n9484.t5 a_1627_n9510.t1 VDDD.t1159 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X834 a_2927_n10028.t1 CLKS.t74 VDDD.t1313 VDDD.t1312 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X835 a_5136_n1029.t1 a_4221_n1029.t5 a_4789_n787.t0 VSSD.t758 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X836 VDDD.t538 CF[5].t7 a_371_n9484.t0 VDDD.t537 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X837 VDDD.t871 a_4821_3799.t4 a_4711_3923.t2 VDDD.t870 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X838 a_n1395_n9484.t0 a_n1561_n9484.t4 VSSD.t1159 VSSD.t870 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X839 a_7602_n9484.t1 CLKS.t75 VSSD.t1013 VSSD.t1012 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X840 a_n7191_n9484.t1 a_n7357_n9484.t6 VDDD.t807 VDDD.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X841 a_n2237_n9724.t2 CLKS.t76 VDDD.t1315 VDDD.t1314 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X842 a_6568_n1573.t1 a_6047_n1599.t4 VDDD.t1044 VDDD.t1043 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X843 a_4410_n4714.t1 a_4366_n5106.t5 a_4244_n4702.t1 VSSD.t93 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X844 VSSD.t921 a_2364_n5482.t6 a_2325_n5356.t0 VSSD.t920 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X845 a_1452_n9650.t2 a_371_n10022.t5 a_1105_n10054.t3 VDDD.t751 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X846 VDDD.t349 a_1024_n4776.t7 DOUT[1].t2 VDDD.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X847 VSSD.t732 a_7423_n9510.t3 a_7357_n9484.t0 VSSD.t303 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X848 a_115_n5372.t3 a_432_n5482.t6 a_390_n5624.t1 VSSD.t993 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X849 a_n2869_n9118.t0 a_n3493_n9484.t3 a_n2977_n9484.t3 VDDD.t1277 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X850 VSSD.t543 COMP_P.t2 a_n10393_n9484.t2 VSSD.t260 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X851 VDDD.t1091 a_n784_n1599.t12 out_latch_0.FINAL.t14 VDDD.t1090 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X852 SWN[7].t2 a_5491_n9724.t5 VDDD.t716 VDDD.t715 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X853 a_5985_n4714.t3 SWP[7].t5 VDDD.t1279 VDDD.t1278 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X854 VSSD.t541 a_6807_n1599.t5 a_6738_n1573.t1 VSSD.t540 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X855 a_4875_n1599.t2 a_4680_n1457.t5 a_5185_n1207.t0 VSSD.t778 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X856 VSSD.t1070 CLKS.t77 a_6765_n1029.t1 VSSD.t1069 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X857 a_5015_n5258.t3 a_4296_n5482.t3 a_4452_n5387.t2 VSSD.t1142 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X858 VSSD.t414 auto_sampling_0.x24.A.t16 CLKS.t8 VSSD.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X859 a_956_2959.t1 a_738_2717.t4 VDDD.t443 VDDD.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X860 a_8931_n4714.t0 EN.t50 VSSD.t1001 VSSD.t1000 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X861 a_n2869_n9118.t2 CLKS.t78 VDDD.t1317 VDDD.t1316 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X862 a_n1543_3557.t1 a_n1709_3557.t5 VDDD.t1162 VDDD.t1161 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X863 a_n8868_n9484.t3 cdac_ctrl_0.x1.X.t28 VDDD.t1453 VDDD.t1452 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X864 VDDD.t990 a_3411_3531.t6 auto_sampling_0.x3.D.t3 VDDD.t989 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X865 a_1413_3557.t1 a_223_3557.t5 a_1304_3557.t3 VSSD.t1194 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X866 a_8670_n1573.t0 a_8583_n1331.t6 a_8266_n1441.t0 VDDD.t1329 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X867 a_8574_3083.t0 EN.t51 VDDD.t1323 VDDD.t1322 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X868 SWN[8].t3 a_7423_n9724.t4 VDDD.t1387 VDDD.t1386 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X869 VDDD.t925 COMP_P.t3 a_n10393_n9484.t3 VDDD.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X870 a_6901_n10054.t3 a_6683_n9650.t5 VDDD.t1196 VDDD.t1195 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X871 a_8117_3557.t1 a_7951_3557.t4 VDDD.t1206 VDDD.t1205 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X872 CF[4].t1 a_7979_n1599.t4 VSSD.t385 VSSD.t384 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X873 a_2671_3557.t2 a_2321_3557.t3 a_2576_3557.t3 VDDD.t1223 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X874 SWP[8].t0 a_7423_n9510.t4 VSSD.t734 VSSD.t733 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X875 SWP[4].t1 a_n305_n9510.t5 VSSD.t736 VSSD.t139 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X876 a_7878_n5624.t1 a_7843_n5372.t4 a_7556_n5650.t1 VSSD.t155 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X877 a_4719_n1331.t1 CLK.t19 VDDD.t1115 VDDD.t1114 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X878 VDDD.t898 a_7423_n9510.t5 a_7410_n9118.t0 VDDD.t897 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X879 a_2544_n1029.t0 CF[9].t6 VSSD.t255 VSSD.t254 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X880 a_6588_n9662.t2 cdac_ctrl_0.x2.X.t25 VSSD.t884 VSSD.t227 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X881 a_8684_2959.t2 a_8466_2717.t4 VDDD.t1170 VDDD.t1169 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X882 out_latch_0.FINAL.t2 a_n784_n1599.t13 VSSD.t858 VSSD.t857 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X883 VDDD.t732 a_7248_n9650.t4 a_7423_n9724.t0 VDDD.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X884 a_8012_n4702.t3 a_7662_n5074.t4 a_7917_n4714.t3 VDDD.t952 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X885 a_284_n4702.t1 a_n66_n5074.t4 a_189_n4714.t0 VDDD.t1276 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X886 a_9302_n1573.t1 a_8544_n1457.t3 a_8739_n1599.t3 VDDD.t841 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X887 a_5490_n1029.t1 CLKS.t79 VSSD.t1068 VSSD.t1067 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X888 VDDD.t1028 a_925_n787.t5 a_815_n663.t1 VDDD.t1027 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X889 a_n3327_n10022.t0 a_n3493_n10022.t5 VSSD.t60 VSSD.t59 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X890 a_537_n10022.t1 a_371_n10022.t6 VDDD.t753 VDDD.t752 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X891 a_n6623_n9242.t2 a_n6841_n9484.t4 VDDD.t459 VDDD.t458 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X892 VDDD.t1325 EN.t52 a_8461_n5258.t0 VDDD.t1324 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X893 a_6529_n5258.t1 a_6315_n5258.t5 VDDD.t957 VDDD.t956 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X894 VSSD.t860 a_n784_n1599.t14 out_latch_0.FINAL.t1 VSSD.t859 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X895 VSSD.t293 a_9175_n1055.t7 CF[5].t0 VSSD.t292 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X896 VSSD.t1129 a_n4169_n9510.t8 a_n4235_n9484.t0 VSSD.t77 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X897 a_1866_n5074.t0 a_1700_n5074.t4 VSSD.t439 VSSD.t438 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X898 a_4751_n9650.t2 a_4401_n10022.t3 a_4656_n9662.t1 VDDD.t1189 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X899 a_2434_n5106.t0 a_2216_n4702.t5 VSSD.t177 VSSD.t176 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X900 VDDD.t69 CKO.t17 a_n232_n5074.t1 VDDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X901 a_573_n1207.t0 a_538_n1441.t4 a_251_n1599.t0 VSSD.t415 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X902 a_n827_n9242.t0 a_n1045_n9484.t4 VSSD.t389 VSSD.t388 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X903 SWP[8].t1 a_7423_n9510.t6 VDDD.t1145 VDDD.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X904 SWP[4].t3 a_n305_n9510.t6 VDDD.t218 VDDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X905 VDDD.t1117 CLK.t20 a_6019_3557.t1 VDDD.t1116 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X906 VSSD.t241 a_8316_n5387.t4 a_8247_n5258.t1 VSSD.t240 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X907 a_6796_2717.t1 a_6752_2959.t5 a_6630_2717.t0 VSSD.t156 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X908 a_6333_n10022.t1 a_6167_n10022.t6 VDDD.t1175 VDDD.t1174 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X909 a_6186_n5624.t1 a_5624_n5650.t5 VSSD.t905 VSSD.t904 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X910 VSSD.t552 a_5311_n1055.t5 a_5245_n1029.t0 VSSD.t551 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X911 a_5342_2691.t1 a_5167_2717.t4 a_5521_2717.t1 VSSD.t296 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X912 VSSD.t800 a_9355_n9724.t7 a_9289_n9650.t1 VSSD.t498 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X913 a_n3990_n9484.t1 CLKS.t80 VSSD.t1066 VSSD.t1024 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X914 VDDD.t978 CF[0].t7 a_n9289_n10022.t0 VDDD.t977 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X915 a_3384_n9484.t3 a_2303_n9484.t4 a_3037_n9242.t3 VDDD.t1079 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X916 VSSD.t10 EN.t53 a_4410_n4714.t0 VSSD.t9 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X917 a_834_2717.t1 a_388_2717.t4 a_738_2717.t2 VSSD.t707 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X918 cdac_ctrl_0.x2.X.t8 a_n10393_n10028.t14 VDDD.t400 VDDD.t399 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X919 a_1614_n10028.t1 a_537_n10022.t4 a_1452_n9650.t0 VDDD.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X920 a_612_n1029.t0 EN.t54 VSSD.t12 VSSD.t11 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X921 VSSD.t14 EN.t55 a_5946_n5624.t0 VSSD.t13 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X922 a_1627_n9510.t0 CLKS.t81 VDDD.t1188 VDDD.t1187 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X923 a_n1543_3557.t0 a_n1709_3557.t6 VSSD.t831 VSSD.t830 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X924 a_n1140_n9662.t3 cdac_ctrl_0.x2.X.t26 VDDD.t1119 VDDD.t1118 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X925 CLKS.t9 auto_sampling_0.x24.A.t17 VDDD.t472 VDDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X926 a_n1288_3557.t2 auto_sampling_0.x21.Q.t4 VSSD.t1187 VSSD.t1186 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X927 a_n1288_3557.t3 auto_sampling_0.x21.Q.t5 VDDD.t1433 VDDD.t1432 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X928 a_n6623_n10054.t1 a_n6841_n9650.t5 VDDD.t1283 VDDD.t1282 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X929 VDDD.t710 a_957_3799.t5 a_847_3923.t1 VDDD.t709 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X930 VDDD.t327 a_5167_2717.t5 a_5342_2691.t2 VDDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X931 a_6315_n5258.t1 a_6228_n5482.t2 a_5911_n5372.t1 VDDD.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X932 VDDD.t1377 a_588_n5387.t4 a_519_n5258.t3 VDDD.t1376 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X933 VDDD.t254 a_8577_n4702.t5 a_8752_n4776.t1 VDDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X934 a_2778_3083.t0 EN.t56 VDDD.t11 VDDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X935 VSSD.t173 a_n10393_n9484.t12 cdac_ctrl_0.x1.X.t4 VSSD.t172 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X936 a_9534_n9484.t1 CLKS.t82 VSSD.t1065 VSSD.t1018 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X937 a_n6733_n10028.t1 a_n7357_n10022.t5 a_n6841_n9650.t3 VDDD.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X938 VSSD.t1064 CLKS.t83 a_6369_n1207.t1 VSSD.t1063 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X939 a_8117_3557.t0 a_7951_3557.t5 VSSD.t947 VSSD.t946 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X940 a_8653_n787.t0 a_8435_n1029.t4 VSSD.t401 VSSD.t400 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X941 a_n10393_n9484.t4 COMP_P.t4 VSSD.t743 VSSD.t418 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X942 a_6342_n4714.t1 a_6298_n5106.t5 a_6176_n4702.t0 VSSD.t330 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X943 a_n8555_n10054.t2 a_n8773_n9650.t4 VDDD.t846 VDDD.t845 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X944 a_8531_n1029.t1 a_8085_n1029.t3 a_8435_n1029.t0 VSSD.t949 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X945 a_n2412_n9650.t3 a_n3327_n10022.t5 a_n2759_n10054.t3 VSSD.t157 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X946 a_4507_2717.t3 auto_sampling_0.x15.D.t4 VDDD.t866 VDDD.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X947 a_n4909_n9484.t2 a_n5425_n9484.t4 a_n5004_n9484.t3 VSSD.t711 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X948 a_4820_2959.t3 a_4602_2717.t4 VDDD.t860 VDDD.t859 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X949 VSSD.t881 CLK.t21 a_4086_2717.t0 VSSD.t880 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X950 VSSD.t92 a_8739_n1599.t4 a_8670_n1573.t2 VSSD.t91 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X951 a_2281_n5258.t0 a_1760_n5650.t4 VDDD.t722 VDDD.t721 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X952 VDDD.t886 a_n10393_n9484.t13 cdac_ctrl_0.x1.X.t12 VDDD.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X953 a_1574_n1573.t0 a_816_n1457.t3 a_1011_n1599.t0 VDDD.t1164 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X954 VDDD.t108 a_7275_3531.t6 auto_sampling_0.x11.D.t2 VDDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X955 a_6947_n5258.t1 a_6228_n5482.t3 a_6384_n5387.t2 VSSD.t608 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X956 a_5277_3557.t0 a_4087_3557.t7 a_5168_3557.t1 VSSD.t1128 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X957 SWP[3].t1 a_n2237_n9510.t4 VSSD.t88 VSSD.t87 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X958 VDDD.t530 a_n2759_n9242.t4 a_n2869_n9118.t1 VDDD.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X959 VDDD.t302 a_n480_n9650.t5 a_n305_n9724.t1 VDDD.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X960 a_1806_n9662.t1 CLKS.t84 VSSD.t1062 VSSD.t1061 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X961 VSSD.t811 a_3410_2691.t5 a_3344_2717.t0 VSSD.t810 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X962 VDDD.t1352 a_n453_3531.t6 auto_sampling_0.x7.Q.t2 VDDD.t1351 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X963 a_n6745_n9650.t0 a_n7191_n10022.t3 a_n6841_n9650.t1 VSSD.t890 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X964 a_4751_n9650.t1 a_4235_n10022.t6 a_4656_n9662.t0 VSSD.t150 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X965 a_n10393_n9484.t5 COMP_P.t5 VDDD.t927 VDDD.t926 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X966 VSSD.t883 CLK.t22 a_6019_3557.t0 VSSD.t882 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X967 VSSD.t664 a_3692_n5650.t5 DOUT[4].t0 VSSD.t663 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X968 a_6535_3557.t1 a_6185_3557.t4 a_6440_3557.t1 VDDD.t532 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X969 a_8085_n1029.t0 a_7919_n1029.t4 VSSD.t510 VSSD.t509 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X970 a_9180_n9650.t2 a_8265_n10022.t4 a_8833_n10054.t1 VSSD.t70 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X971 a_4699_3557.t0 a_4253_3557.t4 a_4603_3557.t3 VSSD.t500 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X972 VSSD.t961 a_1627_n9724.t5 a_1561_n9650.t0 VSSD.t801 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X973 VDDD.t246 a_4719_n1331.t5 a_4680_n1457.t1 VDDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X974 VDDD.t1018 CLK.t23 a_4086_2717.t1 VDDD.t1017 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X975 a_1561_n9650.t1 a_371_n10022.t7 a_1452_n9650.t3 VSSD.t601 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X976 a_2469_n9484.t0 a_2303_n9484.t5 VSSD.t838 VSSD.t790 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X977 VSSD.t875 a_9487_n4848.t3 CKO.t1 VSSD.t874 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X978 a_8265_n9484.t1 a_8099_n9484.t5 VDDD.t20 VDDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X979 a_983_n9484.t0 a_537_n9484.t3 a_887_n9484.t3 VSSD.t591 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X980 SWP[9].t0 a_9355_n9510.t7 VSSD.t1141 VSSD.t798 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X981 SWP[3].t3 a_n2237_n9510.t5 VDDD.t91 VDDD.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X982 a_7370_n1573.t0 a_6651_n1331.t5 a_6807_n1599.t3 VSSD.t1180 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X983 VSSD.t1060 CLKS.t85 a_5013_n9484.t0 VSSD.t1008 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X984 a_n6101_n9724.t0 a_n6276_n9650.t5 a_n5922_n9662.t0 VSSD.t756 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X985 a_n2412_n9484.t3 a_n3493_n9484.t4 a_n2759_n9242.t1 VDDD.t436 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X986 a_5167_2717.t0 a_4086_2717.t6 a_4820_2959.t0 VDDD.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X987 a_6643_3923.t2 a_6019_3557.t5 a_6535_3557.t3 VDDD.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X988 VSSD.t976 SWP[0].t4 a_1151_n5258.t2 VSSD.t975 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X989 a_7117_n1207.t1 a_6738_n1573.t4 a_7045_n1207.t0 VSSD.t530 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X990 a_2216_n4702.t1 a_1700_n5074.t5 a_2121_n4714.t2 VSSD.t440 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X991 a_n8555_n9242.t2 a_n8773_n9484.t5 VSSD.t336 VSSD.t85 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X992 a_n949_n9484.t1 a_n1395_n9484.t4 a_n1045_n9484.t2 VSSD.t590 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X993 VSSD.t16 EN.t57 a_8728_2717.t0 VSSD.t15 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X994 a_9206_2691.t1 a_9031_2717.t4 a_9385_2717.t1 VSSD.t555 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X995 CF[0].t3 a_251_n1599.t7 VDDD.t87 VDDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X996 SWP[9].t2 a_9355_n9510.t8 VDDD.t1372 VDDD.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X997 a_n2303_n9650.t1 a_n3493_n10022.t6 a_n2412_n9650.t0 VSSD.t61 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X998 VSSD.t130 a_n2237_n9724.t5 SWN[3].t0 VSSD.t89 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X999 VDDD.t1358 a_n2237_n9724.t6 SWN[3].t3 VDDD.t1357 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1000 VDDD.t1356 a_8833_n10054.t4 a_8723_n10028.t1 VDDD.t1355 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1001 VDDD.t277 a_3410_2691.t6 a_3397_3083.t1 VDDD.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1002 VSSD.t407 a_5342_2691.t7 auto_sampling_0.x16.D.t0 VSSD.t406 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1003 a_942_n1573.t0 a_816_n1457.t4 a_538_n1441.t1 VSSD.t927 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1004 a_6807_n1599.t2 a_6651_n1331.t6 a_6952_n1573.t0 VDDD.t1427 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1005 a_3559_n9510.t2 CLKS.t86 VDDD.t820 VDDD.t819 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1006 VDDD.t685 a_9031_2717.t5 a_9206_2691.t2 VDDD.t684 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1007 a_8160_n5482.t0 CKO.t18 VSSD.t74 VSSD.t73 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1008 a_6642_3083.t0 EN.t58 VDDD.t13 VDDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1009 DOUT[9].t2 a_8752_n4776.t8 VDDD.t579 VDDD.t578 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1010 a_8541_n1207.t1 a_7979_n1599.t5 VSSD.t387 VSSD.t386 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1011 VSSD.t1151 a_7423_n9724.t5 SWN[8].t0 VSSD.t917 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1012 VSSD.t169 a_n305_n9724.t8 SWN[4].t0 VSSD.t168 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1013 a_8247_n5258.t3 a_8160_n5482.t6 a_7843_n5372.t2 VDDD.t485 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1014 CF[6].t3 a_7243_n1055.t6 VDDD.t1089 VDDD.t1088 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1015 VDDD.t356 a_n8555_n10054.t5 a_n8665_n10028.t1 VDDD.t355 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1016 a_1452_n9650.t1 a_537_n10022.t5 a_1105_n10054.t2 VSSD.t95 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1017 a_4656_n9662.t3 cdac_ctrl_0.x2.X.t27 VDDD.t1121 VDDD.t1120 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1018 VDDD.t822 CLKS.t87 a_1156_n1573.t2 VDDD.t821 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1019 a_6298_n5106.t3 a_6080_n4702.t5 VDDD.t1334 VDDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1020 a_792_n9662.t3 cdac_ctrl_0.x2.X.t28 VDDD.t1123 VDDD.t1122 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1021 a_2927_n9118.t1 CLKS.t88 VDDD.t824 VDDD.t823 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1022 a_n1140_n9662.t2 cdac_ctrl_0.x2.X.t29 VSSD.t885 VSSD.t363 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1023 a_n66_n5074.t1 a_n232_n5074.t3 VDDD.t71 VDDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1024 a_251_n1599.t1 a_538_n1441.t5 VDDD.t476 VDDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1025 a_7274_2691.t2 EN.t59 VDDD.t1198 VDDD.t1197 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1026 CLKS.t10 auto_sampling_0.x24.A.t18 VDDD.t474 VDDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1027 a_6588_n9662.t3 cdac_ctrl_0.x2.X.t30 VDDD.t706 VDDD.t705 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1028 VSSD.t257 CF[9].t7 a_8099_n9484.t0 VSSD.t256 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1029 a_8120_n5080.t1 a_7496_n5074.t2 a_8012_n4702.t0 VDDD.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1030 a_643_2717.t1 auto_sampling_0.x22.A.t6 VDDD.t622 VDDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1031 VDDD.t1020 CLK.t24 a_4087_3557.t1 VDDD.t1019 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1032 a_2857_n787.t2 a_2639_n1029.t5 VDDD.t882 VDDD.t881 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1033 VDDD.t509 a_n975_3799.t4 a_n1085_3923.t1 VDDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1034 VDDD.t726 a_3559_n9724.t6 a_3546_n10028.t0 VDDD.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1035 a_5136_n1029.t2 a_4055_n1029.t3 a_4789_n787.t1 VDDD.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1036 a_3738_n9662.t1 CLKS.t89 VSSD.t1059 VSSD.t1058 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1037 VSSD.t943 EN.t60 a_2932_2717.t0 VSSD.t942 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1038 a_n6114_n10028.t0 a_n7191_n10022.t4 a_n6276_n9650.t1 VDDD.t1168 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1039 DOUT[4].t3 a_3692_n5650.t6 VDDD.t138 VDDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1040 a_942_n1573.t1 a_855_n1331.t6 a_538_n1441.t3 VDDD.t1156 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1041 a_4508_3557.t2 auto_sampling_0.x3.D.t4 VDDD.t734 VDDD.t733 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1042 a_n8677_n9650.t0 a_n9123_n10022.t5 a_n8773_n9650.t2 VSSD.t135 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1043 VDDD.t64 a_1452_n9650.t5 a_1627_n9724.t1 VDDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1044 a_5491_n9510.t1 a_5316_n9484.t5 a_5670_n9484.t0 VSSD.t243 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1045 a_9487_n4848.t0 out_latch_0.FINAL.t18 a_9661_n4742.t0 VSSD.t760 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1046 VSSD.t907 a_5624_n5650.t6 DOUT[6].t0 VSSD.t906 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1047 a_n4344_n9484.t0 a_n5259_n9484.t4 a_n4691_n9242.t0 VSSD.t615 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1048 VDDD.t5 CF[4].t8 a_n1561_n10022.t1 VDDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1049 VSSD.t49 a_1478_2691.t5 auto_sampling_0.x14.D.t0 VSSD.t48 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1050 a_538_n1441.t2 a_855_n1331.t7 a_813_n1207.t0 VSSD.t924 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1051 a_n275_2717.t0 EN.t61 VSSD.t945 VSSD.t944 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1052 a_6797_3557.t1 a_6753_3799.t5 a_6631_3557.t1 VSSD.t528 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1053 a_6315_n5258.t0 a_6189_n5356.t5 a_5911_n5372.t3 VSSD.t939 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1054 a_2781_n4702.t0 a_1700_n5074.t6 a_2434_n5106.t2 VDDD.t938 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1055 VSSD.t815 a_6047_n1599.t5 CF[3].t1 VSSD.t814 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1056 a_5343_3531.t2 a_5168_3557.t5 a_5522_3557.t1 VSSD.t770 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1057 VDDD.t378 a_3379_n1055.t7 CF[8].t0 VDDD.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1058 a_2819_n9650.t3 a_2469_n10022.t4 a_2724_n9662.t0 VDDD.t524 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1059 VDDD.t1010 a_9355_n9724.t8 a_9342_n10028.t0 VDDD.t1009 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1060 a_835_3557.t1 a_389_3557.t3 a_739_3557.t3 VSSD.t20 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1061 VDDD.t668 CF[2].t7 a_n5425_n9484.t1 VDDD.t667 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1062 a_n6101_n9724.t2 CLKS.t90 VDDD.t848 VDDD.t847 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1063 VDDD.t1288 CF[3].t7 a_n3493_n10022.t1 VDDD.t1287 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1064 VDDD.t1299 a_4969_n9242.t4 a_4859_n9118.t2 VDDD.t1298 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1065 a_432_n5482.t0 CKO.t19 VSSD.t205 VSSD.t204 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1066 a_6683_n9484.t2 a_6167_n9484.t5 a_6588_n9484.t2 VSSD.t201 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1067 a_1249_n1207.t1 CLKS.t91 VSSD.t1057 VSSD.t1056 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1068 VSSD.t122 auto_sampling_0.x23.A.t8 auto_sampling_0.x24.A.t2 VSSD.t121 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1069 a_n784_n1599.t4 CF[0].t8 VDDD.t980 VDDD.t979 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1070 a_6228_n5482.t1 CKO.t20 VDDD.t224 VDDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1071 a_9049_n1207.t1 a_8670_n1573.t5 a_8977_n1207.t0 VSSD.t297 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1072 CF[9].t3 a_1447_n1055.t6 VDDD.t230 VDDD.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1073 VDDD.t1290 CF[3].t8 a_5438_n1573.t3 VDDD.t1289 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1074 a_4148_n4702.t1 a_3632_n5074.t6 a_4053_n4714.t0 VSSD.t374 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1075 a_6779_n9650.t1 a_6333_n10022.t4 a_6683_n9650.t3 VSSD.t443 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1076 a_n784_n1599.t0 CF[0].t9 VDDD.t423 VDDD.t422 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1077 a_2927_n9118.t2 a_2303_n9484.t6 a_2819_n9484.t3 VDDD.t1080 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1078 VDDD.t1327 a_1011_n1599.t5 a_942_n1573.t3 VDDD.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1079 a_3493_n9484.t0 a_2303_n9484.t7 a_3384_n9484.t2 VSSD.t839 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1080 VSSD.t611 a_588_n5387.t5 a_519_n5258.t0 VSSD.t610 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1081 VDDD.t55 a_7274_2691.t5 a_7261_3083.t1 VDDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1082 VSSD.t723 a_9206_2691.t8 auto_sampling_0.x21.Q.t0 VSSD.t722 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1083 a_6440_3557.t2 auto_sampling_0.x5.D.t5 VSSD.t642 VSSD.t641 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1084 VDDD.t1093 a_n784_n1599.t15 out_latch_0.FINAL.t13 VDDD.t1092 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1085 VSSD.t431 a_4888_n4776.t5 a_4822_n4702.t1 VSSD.t430 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1086 cdac_ctrl_0.x2.X.t9 a_n10393_n10028.t15 VSSD.t350 VSSD.t349 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1087 a_3037_n10054.t1 a_2819_n9650.t5 VSSD.t179 VSSD.t178 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1088 VDDD.t216 a_2434_n5106.t5 a_2324_n5080.t2 VDDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1089 a_849_n4702.t2 a_n232_n5074.t4 a_502_n5106.t1 VDDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1090 a_1478_2691.t0 EN.t62 VDDD.t1200 VDDD.t1199 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1091 VSSD.t433 a_4888_n4776.t6 DOUT[5].t1 VSSD.t432 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1092 VDDD.t279 a_3410_2691.t7 auto_sampling_0.x15.D.t2 VDDD.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1093 DOUT[2].t1 a_1760_n5650.t5 VSSD.t714 VSSD.t713 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1094 VSSD.t287 a_n6101_n9724.t6 a_n6167_n9650.t0 VSSD.t286 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1095 VSSD.t371 CF[0].t10 a_n9289_n9484.t0 VSSD.t370 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1096 VDDD.t1022 CLK.t25 a_2123_n1029.t1 VDDD.t1021 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1097 a_5013_n9484.t1 a_4969_n9242.t5 a_4847_n9484.t1 VSSD.t926 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1098 a_5329_3083.t0 a_4252_2717.t4 a_5167_2717.t3 VDDD.t972 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1099 a_n6936_n9484.t3 cdac_ctrl_0.x1.X.t29 VSSD.t896 VSSD.t625 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1100 VDDD.t1202 EN.t63 a_n172_n5650.t2 VDDD.t1201 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1101 VSSD.t373 CF[0].t11 a_n784_n1599.t1 VSSD.t372 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1102 a_7243_n1055.t0 CLKS.t92 VDDD.t850 VDDD.t849 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1103 a_3559_n9724.t2 CLKS.t93 VDDD.t852 VDDD.t851 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1104 VSSD.t804 CLK.t26 a_4087_3557.t0 VSSD.t803 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1105 a_956_2959.t0 a_738_2717.t5 VSSD.t909 VSSD.t908 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1106 VSSD.t983 SWP[8].t5 a_8879_n5258.t0 VSSD.t982 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1107 a_8340_n1029.t2 CF[6].t6 VDDD.t134 VDDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1108 a_6952_n1573.t1 a_6738_n1573.t5 VDDD.t651 VDDD.t650 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1109 a_612_n1029.t1 EN.t64 VDDD.t1204 VDDD.t1203 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1110 a_7423_n9724.t1 a_7248_n9650.t5 a_7602_n9662.t0 VSSD.t584 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1111 a_n4235_n9484.t1 a_n5425_n9484.t5 a_n4344_n9484.t2 VSSD.t426 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1112 auto_sampling_0.x21.D.t0 a_7274_2691.t6 VSSD.t56 VSSD.t55 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1113 a_n467_3083.t1 a_n1544_2717.t4 a_n629_2717.t0 VDDD.t430 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1114 a_2956_n4776.t2 a_2781_n4702.t5 a_3135_n4714.t1 VSSD.t988 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1115 VSSD.t952 a_3411_3531.t7 a_3345_3557.t1 VSSD.t951 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1116 a_n827_n10054.t2 a_n1045_n9650.t4 VDDD.t588 VDDD.t587 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1117 VDDD.t479 COMP_N.t4 a_n10393_n10028.t4 VDDD.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1118 a_5491_n9724.t2 CLKS.t94 VDDD.t262 VDDD.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1119 VDDD.t439 a_9032_3557.t4 a_9207_3531.t1 VDDD.t438 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1120 a_6643_3923.t0 EN.t65 VDDD.t625 VDDD.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1121 a_5911_n5372.t0 a_6228_n5482.t4 a_6186_n5624.t0 VSSD.t609 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1122 a_n1086_3083.t1 a_n1710_2717.t3 a_n1194_2717.t2 VDDD.t1171 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1123 a_n126_n9484.t1 CLKS.t95 VSSD.t1055 VSSD.t1006 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1124 a_n1045_n9484.t1 a_n1561_n9484.t5 a_n1140_n9484.t0 VSSD.t284 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1125 a_8230_n5106.t3 a_8012_n4702.t5 VDDD.t570 VDDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1126 out_latch_0.FINAL.t0 a_n784_n1599.t16 VSSD.t1191 VSSD.t1190 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1127 a_4053_n4714.t2 SWP[5].t5 VDDD.t796 VDDD.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1128 VSSD.t1054 CLKS.t96 a_n2715_n9484.t1 VSSD.t1053 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1129 a_1149_n9662.t0 a_1105_n10054.t5 a_983_n9650.t0 VSSD.t133 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1130 a_n4801_n10028.t1 CLKS.t97 VDDD.t264 VDDD.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1131 a_8520_n9484.t2 cdac_ctrl_0.x1.X.t30 VSSD.t898 VSSD.t897 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1132 a_n6841_n9650.t2 a_n7357_n10022.t6 a_n6936_n9662.t3 VSSD.t4 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1133 VDDD.t963 a_7979_n1599.t6 CF[4].t2 VDDD.t962 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1134 a_4571_n1029.t2 a_4055_n1029.t4 a_4476_n1029.t3 VSSD.t109 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1135 a_3083_n5258.t1 a_2364_n5482.t7 a_2520_n5387.t0 VSSD.t922 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1136 a_1866_n5074.t1 a_1700_n5074.t7 VDDD.t940 VDDD.t939 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1137 a_6721_n787.t1 a_6503_n1029.t5 VDDD.t518 VDDD.t517 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1138 a_9000_n1029.t0 a_7919_n1029.t5 a_8653_n787.t2 VDDD.t623 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1139 a_4690_n5624.t0 EN.t66 VSSD.t512 VSSD.t511 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1140 VSSD.t514 EN.t67 a_6796_2717.t0 VSSD.t513 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1141 VDDD.t1389 SWP[2].t5 a_3083_n5258.t3 VDDD.t1388 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1142 a_8372_3557.t2 auto_sampling_0.x11.D.t5 VDDD.t376 VDDD.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1143 a_8615_n9484.t1 a_8265_n9484.t4 a_8520_n9484.t0 VDDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1144 a_n7191_n10022.t1 a_n7357_n10022.t7 VDDD.t7 VDDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1145 VDDD.t24 a_n8033_n9724.t5 a_n8046_n10028.t0 VDDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1146 a_3384_n9484.t1 a_2469_n9484.t5 a_3037_n9242.t2 VSSD.t589 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1147 a_1381_n1029.t1 a_191_n1029.t5 a_1272_n1029.t1 VSSD.t325 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1148 a_2520_n5387.t2 a_2325_n5356.t4 a_2830_n5624.t1 VSSD.t842 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1149 a_n1194_2717.t0 a_n1544_2717.t5 a_n1289_2717.t0 VDDD.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1150 DOUT[6].t3 a_5624_n5650.t7 VDDD.t1139 VDDD.t1138 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1151 VDDD.t45 a_1478_2691.t6 a_1465_3083.t0 VDDD.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1152 a_8684_2959.t1 a_8466_2717.t5 VSSD.t862 VSSD.t861 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1153 VDDD.t920 a_4820_2959.t4 a_4710_3083.t2 VDDD.t919 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1154 a_357_n1029.t0 a_191_n1029.t6 VSSD.t327 VSSD.t326 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1155 VDDD.t1135 a_3204_n1029.t4 a_3379_n1055.t0 VDDD.t1134 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1156 a_n6276_n9484.t3 a_n7191_n9484.t3 a_n6623_n9242.t3 VSSD.t889 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1157 CF[3].t0 a_6047_n1599.t6 VSSD.t817 VSSD.t816 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1158 VSSD.t516 EN.t68 a_8729_3557.t0 VSSD.t515 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1159 VDDD.t266 CLKS.t98 a_8884_n1573.t2 VDDD.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1160 a_9207_3531.t2 a_9032_3557.t5 a_9386_3557.t1 VSSD.t390 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1161 VDDD.t1087 a_7243_n1055.t7 a_7230_n663.t0 VDDD.t1086 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1162 a_8833_n9242.t2 a_8615_n9484.t4 VSSD.t962 VSSD.t344 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1163 a_n5259_n9484.t0 a_n5425_n9484.t6 VDDD.t834 VDDD.t833 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1164 a_8752_n4776.t0 EN.t69 VDDD.t627 VDDD.t626 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1165 a_2901_n1029.t0 a_2857_n787.t4 a_2735_n1029.t1 VSSD.t134 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1166 a_537_n9484.t1 a_371_n9484.t4 VDDD.t1404 VDDD.t1403 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1167 a_2312_n4702.t1 a_1866_n5074.t4 a_2216_n4702.t2 VSSD.t451 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1168 a_n8868_n9662.t2 cdac_ctrl_0.x2.X.t31 VSSD.t568 VSSD.t365 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1169 VSSD.t3 CF[4].t9 a_n1561_n9484.t0 VSSD.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1170 VSSD.t484 a_5343_3531.t7 auto_sampling_0.x5.D.t0 VSSD.t483 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1171 VSSD.t125 CF[6].t7 a_2303_n10022.t0 VSSD.t123 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1172 a_n937_n9118.t1 a_n1561_n9484.t6 a_n1045_n9484.t0 VDDD.t1394 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1173 a_1447_n1055.t2 CLKS.t99 VDDD.t969 VDDD.t968 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1174 VDDD.t85 CF[1].t6 a_n7357_n9484.t0 VDDD.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1175 VDDD.t766 a_6228_n5482.t5 a_6189_n5356.t0 VDDD.t765 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1176 CF[7].t2 a_5311_n1055.t6 VDDD.t681 VDDD.t680 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1177 a_9032_3557.t0 a_7951_3557.t6 a_8685_3799.t0 VDDD.t1207 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1178 SWN[0].t1 a_n8033_n9724.t6 VSSD.t33 VSSD.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1179 a_2544_n1029.t1 CF[9].t8 VDDD.t1381 VDDD.t1380 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1180 a_n520_2717.t1 a_n1710_2717.t4 a_n629_2717.t2 VSSD.t930 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1181 a_2943_n1599.t2 a_2748_n1457.t4 a_3253_n1207.t1 VSSD.t660 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1182 auto_sampling_0.x14.D.t1 a_1478_2691.t7 VSSD.t51 VSSD.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1183 a_1303_2717.t1 a_388_2717.t5 a_956_2959.t2 VSSD.t708 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1184 VDDD.t335 a_7423_n9724.t6 SWN[8].t2 VDDD.t334 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1185 a_6999_n4714.t0 EN.t70 VSSD.t518 VSSD.t517 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1186 VDDD.t971 CLKS.t100 a_7979_n1599.t2 VDDD.t970 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1187 a_357_n1029.t1 a_191_n1029.t7 VDDD.t365 VDDD.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1188 a_4875_n5080.t1 a_3798_n5074.t3 a_4713_n4702.t2 VDDD.t911 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1189 out_latch_0.FINAL.t12 a_n784_n1599.t17 VDDD.t1441 VDDD.t1440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1190 a_4859_n9118.t0 a_4235_n9484.t5 a_4751_n9484.t0 VDDD.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1191 SWN[5].t3 a_1627_n9724.t6 VDDD.t1032 VDDD.t1031 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1192 VDDD.t451 a_3236_3557.t4 a_3411_3531.t2 VDDD.t450 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1193 VDDD.t1111 a_9180_n9484.t5 a_9355_n9510.t1 VDDD.t1110 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1194 DOUT[5].t0 a_4888_n4776.t7 VSSD.t435 VSSD.t434 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1195 VDDD.t728 a_7274_2691.t7 auto_sampling_0.x21.D.t2 VDDD.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1196 VSSD.t90 a_n2237_n9510.t6 SWP[3].t0 VSSD.t89 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1197 VDDD.t1024 CLK.t27 a_5987_n1029.t1 VDDD.t1023 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1198 a_7556_n5650.t2 a_7843_n5372.t5 VDDD.t163 VDDD.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1199 a_n172_n5650.t1 a_115_n5372.t5 VDDD.t789 VDDD.t788 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1200 VDDD.t198 a_n454_2691.t7 auto_sampling_0.x22.A.t2 VDDD.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1201 a_n2977_n9484.t2 a_n3327_n9484.t4 a_n3072_n9484.t3 VDDD.t1226 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1202 a_n2715_n9484.t0 a_n2759_n9242.t5 a_n2881_n9484.t1 VSSD.t142 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1203 a_925_n787.t2 a_707_n1029.t5 VDDD.t457 VDDD.t456 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1204 a_4820_2959.t2 a_4602_2717.t5 VSSD.t681 VSSD.t680 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1205 a_6945_n9484.t0 a_6901_n9242.t5 a_6779_n9484.t0 VSSD.t505 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1206 a_2576_3557.t2 auto_sampling_0.x2.D.t5 VDDD.t996 VDDD.t995 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1207 a_8977_n1207.t1 CLKS.t101 VSSD.t1052 VSSD.t1051 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1208 a_1272_n1029.t3 a_357_n1029.t5 a_925_n787.t3 VSSD.t866 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1209 VSSD.t80 a_3559_n9724.t7 SWN[6].t0 VSSD.t79 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1210 VDDD.t586 a_6384_n5387.t4 a_6315_n5258.t3 VDDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1211 a_4762_n5624.t1 a_4383_n5258.t4 a_4690_n5624.t1 VSSD.t703 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1212 VDDD.t393 a_6645_n4702.t5 a_6820_n4776.t2 VDDD.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1213 VSSD.t918 a_7423_n9510.t7 SWP[8].t2 VSSD.t917 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1214 VDDD.t299 a_n827_n10054.t5 a_n937_n10028.t1 VDDD.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1215 VSSD.t198 a_n305_n9510.t7 SWP[4].t0 VSSD.t168 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1216 VDDD.t93 a_n2237_n9510.t7 SWP[3].t2 VDDD.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1217 a_2704_n1573.t0 a_2183_n1599.t7 VDDD.t1265 VDDD.t1264 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1218 a_4888_n4776.t2 a_4713_n4702.t5 a_5067_n4714.t1 VSSD.t837 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1219 VSSD.t1121 EN.t71 a_2933_3557.t0 VSSD.t1120 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1220 VDDD.t1309 a_1447_n1055.t7 a_1434_n663.t0 VDDD.t1308 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1221 a_8686_n4702.t1 a_7496_n5074.t3 a_8577_n4702.t0 VSSD.t408 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1222 a_1105_n9242.t1 a_887_n9484.t5 VSSD.t828 VSSD.t493 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1223 VDDD.t402 a_n10393_n10028.t16 cdac_ctrl_0.x2.X.t10 VDDD.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1224 VDDD.t1034 a_1627_n9724.t7 a_1614_n10028.t0 VDDD.t1033 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1225 a_n2977_n9484.t0 a_n3493_n9484.t5 a_n3072_n9484.t0 VSSD.t58 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1226 a_6901_n9242.t3 a_6683_n9484.t5 VDDD.t1082 VDDD.t1081 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1227 VSSD.t461 a_1479_3531.t6 auto_sampling_0.x2.D.t1 VSSD.t460 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1228 a_392_n5080.t0 EN.t72 VDDD.t1345 VDDD.t1344 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1229 VSSD.t334 a_3379_n1055.t8 a_3313_n1029.t0 VSSD.t333 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1230 VSSD.t1050 CLKS.t102 a_2901_n1029.t1 VSSD.t1049 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1231 VSSD.t1048 CLKS.t103 a_n4647_n9484.t1 VSSD.t1047 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1232 VDDD.t1147 a_7423_n9510.t8 SWP[8].t3 VDDD.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1233 VSSD.t1046 CLKS.t104 a_6945_n9662.t1 VSSD.t1045 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1234 VSSD.t456 a_9487_n5472.t3 CKO.t2 VSSD.t455 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1235 a_1452_n9484.t1 a_371_n9484.t5 a_1105_n9242.t0 VDDD.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1236 VDDD.t220 a_n305_n9510.t8 SWP[4].t2 VDDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1237 a_n8773_n9650.t1 a_n9289_n10022.t6 a_n8868_n9662.t0 VSSD.t116 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1238 a_8879_n5258.t2 a_8121_n5356.t4 a_8316_n5387.t1 VDDD.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1239 VSSD.t449 CF[5].t8 a_371_n9484.t1 VSSD.t447 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1240 a_392_n5080.t1 a_n232_n5074.t5 a_284_n4702.t2 VDDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1241 a_5521_2717.t0 EN.t73 VSSD.t1123 VSSD.t1122 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1242 a_7248_n9650.t0 a_6167_n10022.t7 a_6901_n10054.t0 VDDD.t1176 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1243 a_n7191_n9484.t0 a_n7357_n9484.t7 VSSD.t572 VSSD.t521 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1244 a_n2237_n9510.t0 a_n2412_n9484.t4 a_n2058_n9484.t0 VSSD.t380 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1245 VDDD.t559 a_956_2959.t5 a_846_3083.t1 VDDD.t558 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1246 a_n827_n10054.t3 a_n1045_n9650.t5 VSSD.t489 VSSD.t388 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1247 auto_sampling_0.x24.A.t3 auto_sampling_0.x23.A.t9 VDDD.t190 VDDD.t189 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1248 VDDD.t653 a_6820_n4776.t7 DOUT[7].t3 VDDD.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1249 VSSD.t1125 EN.t74 a_n932_2717.t0 VSSD.t1124 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1250 a_n629_2717.t3 a_n1710_2717.t5 a_n976_2959.t3 VDDD.t1172 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1251 a_4014_n5624.t1 a_3979_n5372.t4 a_3692_n5650.t1 VSSD.t593 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1252 VDDD.t1155 a_n4344_n9484.t4 a_n4169_n9510.t1 VDDD.t1154 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1253 a_n976_2959.t2 a_n1194_2717.t5 VDDD.t549 VDDD.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1254 VSSD.t1044 CLKS.t105 a_4437_n1207.t0 VSSD.t1043 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1255 VSSD.t226 a_9207_3531.t7 auto_sampling_0.x11.Q.t0 VSSD.t225 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1256 a_n8665_n9118.t0 a_n9289_n9484.t6 a_n8773_n9484.t3 VDDD.t793 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1257 DOUT[0].t0 a_n172_n5650.t8 VSSD.t640 VSSD.t639 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1258 a_4833_n1029.t0 a_4789_n787.t5 a_4667_n1029.t1 VSSD.t244 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1259 a_2724_n9662.t1 cdac_ctrl_0.x2.X.t32 VSSD.t569 VSSD.t97 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1260 a_4452_n5387.t3 a_4296_n5482.t4 a_4597_n5258.t2 VDDD.t1373 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1261 a_n4647_n9662.t0 a_n4691_n10054.t5 a_n4813_n9650.t1 VSSD.t464 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1262 a_8877_n9662.t0 a_8833_n10054.t5 a_8711_n9650.t0 VSSD.t452 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1263 a_4244_n4702.t0 a_3798_n5074.t4 a_4148_n4702.t3 VSSD.t737 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1264 auto_sampling_0.x23.A.t2 auto_sampling_0.x22.A.t7 VDDD.t769 VDDD.t768 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1265 a_6599_n1029.t1 a_6153_n1029.t4 a_6503_n1029.t0 VSSD.t62 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1266 VDDD.t557 a_1479_3531.t7 a_1466_3923.t0 VDDD.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1267 a_2320_2717.t0 a_2154_2717.t5 VSSD.t397 VSSD.t396 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1268 VDDD.t168 a_8160_n5482.t7 a_8121_n5356.t1 VDDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1269 a_5167_2717.t2 a_4252_2717.t5 a_4820_2959.t1 VSSD.t772 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1270 a_n2759_n9242.t3 a_n2977_n9484.t5 VDDD.t62 VDDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1271 VSSD.t554 a_5311_n1055.t7 CF[7].t1 VSSD.t553 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1272 a_7979_n1599.t1 a_8266_n1441.t5 VDDD.t1397 VDDD.t1396 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1273 a_n931_3557.t1 a_n975_3799.t5 a_n1097_3557.t1 VSSD.t361 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1274 VDDD.t890 a_n827_n9242.t4 a_n937_n9118.t0 VDDD.t889 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1275 a_9162_n663.t1 a_8085_n1029.t4 a_9000_n1029.t1 VDDD.t1208 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1276 VDDD.t102 a_7100_3557.t5 a_7275_3531.t2 VDDD.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1277 a_738_2717.t1 a_222_2717.t7 a_643_2717.t2 VSSD.t670 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1278 a_957_3799.t1 a_739_3557.t5 VSSD.t299 VSSD.t298 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1279 VSSD.t1131 a_n453_3531.t7 a_n519_3557.t1 VSSD.t1130 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1280 a_4711_3923.t0 EN.t75 VDDD.t1347 VDDD.t1346 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1281 a_2322_n5624.t0 a_1760_n5650.t6 VSSD.t716 VSSD.t715 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1282 a_9487_n4848.t2 CLKS.t106 VDDD.t913 VDDD.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1283 auto_sampling_0.x22.A.t0 a_n454_2691.t8 VSSD.t185 VSSD.t184 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1284 VSSD.t753 a_5491_n9724.t6 a_5425_n9650.t1 VSSD.t566 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1285 a_8577_n4702.t3 a_7662_n5074.t5 a_8230_n5106.t1 VSSD.t763 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1286 VSSD.t796 a_2787_n1331.t5 a_2748_n1457.t0 VSSD.t795 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1287 a_n6114_n9118.t1 a_n7191_n9484.t4 a_n6276_n9484.t2 VDDD.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1288 a_2819_n9650.t0 a_2303_n10022.t4 a_2724_n9662.t3 VSSD.t190 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1289 a_2047_n5372.t1 a_2325_n5356.t5 a_2281_n5258.t1 VDDD.t1083 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1290 auto_sampling_0.x11.D.t0 a_7275_3531.t7 VSSD.t103 VSSD.t102 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1291 a_7100_3557.t2 a_6185_3557.t5 a_6753_3799.t1 VSSD.t446 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1292 CLKS.t0 auto_sampling_0.x24.A.t19 VSSD.t159 VSSD.t158 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1293 a_n4909_n9650.t2 a_n5259_n10022.t3 a_n5004_n9662.t1 VDDD.t981 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1294 a_6738_n1573.t2 a_6612_n1457.t4 a_6334_n1441.t2 VSSD.t863 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1295 a_6534_2717.t3 a_6184_2717.t5 a_6439_2717.t3 VDDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1296 a_2320_2717.t1 a_2154_2717.t6 VDDD.t844 VDDD.t843 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1297 cdac_ctrl_0.x1.X.t3 a_n10393_n9484.t14 VSSD.t720 VSSD.t349 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1298 VSSD.t1127 EN.t76 a_2082_n5624.t0 VSSD.t1126 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1299 VSSD.t1042 CLKS.t107 a_n6579_n9662.t0 VSSD.t1041 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1300 a_8340_n1029.t1 CF[6].t8 VSSD.t575 VSSD.t574 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1301 a_5478_n10028.t1 a_4401_n10022.t4 a_5316_n9650.t3 VDDD.t1190 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1302 a_n4909_n9484.t0 a_n5259_n9484.t5 a_n5004_n9484.t0 VDDD.t767 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1303 a_n4344_n9650.t1 a_n5425_n10022.t5 a_n4691_n10054.t0 VDDD.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1304 a_n6841_n9650.t0 a_n7191_n10022.t5 a_n6936_n9662.t0 VDDD.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1305 a_n2237_n9510.t2 CLKS.t108 VDDD.t915 VDDD.t914 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1306 a_n9123_n10022.t1 a_n9289_n10022.t7 VSSD.t742 VSSD.t631 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1307 VSSD.t754 a_5491_n9724.t7 SWN[7].t1 VSSD.t602 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1308 a_n480_n9484.t3 a_n1561_n9484.t7 a_n827_n9242.t2 VDDD.t1395 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1309 a_7662_n5074.t0 a_7496_n5074.t4 VSSD.t410 VSSD.t409 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1310 a_9194_3923.t1 a_8117_3557.t4 a_9032_3557.t3 VDDD.t1364 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1311 a_5670_n9484.t1 CLKS.t109 VSSD.t1040 VSSD.t1039 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1312 VDDD.t41 a_8316_n5387.t5 a_8247_n5258.t0 VDDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1313 VSSD.t690 EN.t77 a_6797_3557.t0 VSSD.t689 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1314 a_6642_3083.t1 a_6018_2717.t5 a_6534_2717.t1 VDDD.t357 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1315 a_7410_n10028.t1 a_6333_n10022.t5 a_7248_n9650.t2 VDDD.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1316 cdac_ctrl_0.x1.X.t11 a_n10393_n9484.t15 VDDD.t888 VDDD.t887 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1317 VDDD.t449 a_8653_n787.t5 a_8543_n663.t1 VDDD.t448 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1318 a_9140_2717.t1 a_7950_2717.t6 a_9031_2717.t0 VSSD.t237 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1319 a_4636_n1573.t1 a_4115_n1599.t6 VDDD.t1254 VDDD.t1253 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1320 a_n1086_3083.t0 EN.t78 VDDD.t869 VDDD.t868 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1321 VDDD.t433 a_n629_2717.t4 a_n454_2691.t1 VDDD.t432 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1322 VDDD.t718 CF[6].t9 a_2303_n10022.t1 VDDD.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1323 VDDD.t75 a_n8208_n9650.t5 a_n8033_n9724.t0 VDDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1324 a_n5259_n10022.t1 a_n5425_n10022.t6 VDDD.t774 VDDD.t773 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1325 a_n371_n9650.t0 a_n1561_n10022.t6 a_n480_n9650.t3 VSSD.t285 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1326 a_8685_3799.t2 a_8467_3557.t5 VSSD.t369 VSSD.t368 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1327 VDDD.t1000 a_3037_n10054.t5 a_2927_n10028.t0 VDDD.t999 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1328 a_8833_n9242.t3 a_8615_n9484.t5 VDDD.t1236 VDDD.t1235 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1329 VSSD.t702 a_4875_n1599.t5 a_4806_n1573.t2 VSSD.t701 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1330 a_7423_n9510.t2 CLKS.t110 VDDD.t312 VDDD.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1331 a_8562_2717.t0 a_8116_2717.t4 a_8466_2717.t3 VSSD.t338 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1332 a_792_n9484.t2 cdac_ctrl_0.x1.X.t31 VSSD.t900 VSSD.t899 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1333 VDDD.t89 a_251_n1599.t8 CF[0].t2 VDDD.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1334 a_9289_n9650.t0 a_8099_n10022.t7 a_9180_n9650.t1 VSSD.t22 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1335 VSSD.t1038 CLKS.t111 a_8877_n9662.t1 VSSD.t1037 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1336 a_9385_2717.t0 EN.t79 VSSD.t692 VSSD.t691 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1337 a_n6936_n9484.t2 cdac_ctrl_0.x1.X.t32 VDDD.t661 VDDD.t660 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1338 SWN[2].t2 a_n4169_n9724.t7 VDDD.t79 VDDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1339 a_9000_n1029.t2 a_8085_n1029.t5 a_8653_n787.t3 VSSD.t950 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1340 a_3366_n663.t1 a_2289_n1029.t5 a_3204_n1029.t0 VDDD.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1341 VSSD.t352 a_n10393_n10028.t17 cdac_ctrl_0.x2.X.t11 VSSD.t351 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1342 a_887_n9484.t2 a_537_n9484.t4 a_792_n9484.t1 VDDD.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1343 a_n8555_n10054.t0 a_n8773_n9650.t5 VSSD.t86 VSSD.t85 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1344 VDDD.t1443 a_n784_n1599.t18 out_latch_0.FINAL.t11 VDDD.t1442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1345 a_4221_n1029.t0 a_4055_n1029.t5 VSSD.t111 VSSD.t110 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1346 a_n2058_n9662.t1 CLKS.t112 VSSD.t1036 VSSD.t1035 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1347 DOUT[7].t2 a_6820_n4776.t8 VDDD.t655 VDDD.t654 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1348 VDDD.t136 a_8685_3799.t5 a_8575_3923.t2 VDDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1349 a_n1193_3557.t3 a_n1709_3557.t7 a_n1288_3557.t1 VSSD.t829 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1350 a_n4169_n9510.t0 a_n4344_n9484.t5 a_n3990_n9484.t0 VSSD.t560 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1351 a_6609_n1207.t1 a_6047_n1599.t7 VSSD.t819 VSSD.t818 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1352 cdac_ctrl_0.x2.X.t12 a_n10393_n10028.t18 VSSD.t353 VSSD.t246 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1353 auto_sampling_0.x2.D.t0 a_1479_3531.t8 VSSD.t463 VSSD.t462 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1354 VDDD.t314 CLKS.t113 a_5020_n1573.t1 VDDD.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1355 a_1304_3557.t1 a_389_3557.t4 a_957_3799.t3 VSSD.t21 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1356 a_6334_n1441.t3 a_6651_n1331.t7 a_6609_n1207.t0 VSSD.t1181 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1357 out_latch_0.FINAL.t10 a_n784_n1599.t19 VDDD.t1445 VDDD.t1444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1358 a_4401_n9484.t1 a_4235_n9484.t6 VDDD.t153 VDDD.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1359 a_5946_n5624.t1 a_5911_n5372.t5 a_5624_n5650.t2 VSSD.t214 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1360 a_6184_2717.t0 a_6018_2717.t6 VSSD.t323 VSSD.t322 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1361 VDDD.t702 a_5491_n9510.t6 a_5478_n9118.t0 VDDD.t701 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1362 a_3506_n1573.t0 a_2787_n1331.t6 a_2943_n1599.t0 VSSD.t797 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1363 a_6503_n1029.t1 a_6153_n1029.t5 a_6408_n1029.t1 VDDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1364 a_4656_n9662.t2 cdac_ctrl_0.x2.X.t33 VSSD.t571 VSSD.t570 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1365 VSSD.t1031 CLKS.t114 a_1149_n9484.t1 VSSD.t1030 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1366 a_6384_n5387.t3 a_6228_n5482.t6 a_6529_n5258.t2 VDDD.t955 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1367 a_n6579_n9662.t1 a_n6623_n10054.t4 a_n6745_n9650.t1 VSSD.t151 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1368 CF[7].t0 a_5311_n1055.t8 VSSD.t181 VSSD.t180 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1369 VDDD.t836 a_3037_n9242.t4 a_2927_n9118.t0 VDDD.t835 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1370 a_7370_n1573.t3 a_6612_n1457.t5 a_6807_n1599.t0 VDDD.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1371 a_n4691_n9242.t2 a_n4909_n9484.t5 VSSD.t836 VSSD.t834 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1372 VSSD.t183 CF[5].t9 a_9302_n1573.t2 VSSD.t182 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1373 SWP[0].t1 a_n8033_n9510.t5 VSSD.t964 VSSD.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1374 VDDD.t1238 a_n8555_n9242.t4 a_n8665_n9118.t1 VDDD.t1237 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1375 a_4821_3799.t2 a_4603_3557.t5 VSSD.t706 VSSD.t705 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1376 a_n1395_n10022.t1 a_n1561_n10022.t7 VSSD.t871 VSSD.t870 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1377 a_4597_n5258.t1 a_4383_n5258.t5 VDDD.t873 VDDD.t872 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1378 a_3398_3923.t1 a_2321_3557.t4 a_3236_3557.t3 VDDD.t1224 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1379 a_7602_n9662.t1 CLKS.t115 VSSD.t1034 VSSD.t1012 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1380 VSSD.t925 a_n2237_n9510.t8 a_n2303_n9484.t0 VSSD.t127 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1381 a_2321_3557.t1 a_2155_3557.t5 VDDD.t659 VDDD.t658 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1382 VDDD.t929 a_n6101_n9510.t8 a_n6114_n9118.t0 VDDD.t928 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1383 VDDD.t170 CLKS.t116 a_251_n1599.t2 VDDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1384 VSSD.t175 auto_sampling_0.x23.A.t10 auto_sampling_0.x24.A.t4 VSSD.t174 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1385 VSSD.t486 a_6384_n5387.t5 a_6315_n5258.t2 VSSD.t485 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1386 VDDD.t453 a_2857_n787.t5 a_2747_n663.t1 VDDD.t452 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1387 a_3344_2717.t1 a_2154_2717.t7 a_3235_2717.t2 VSSD.t671 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1388 a_4254_n5624.t0 a_3692_n5650.t7 VSSD.t132 VSSD.t131 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1389 a_6611_n663.t1 a_5987_n1029.t6 a_6503_n1029.t3 VDDD.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1390 a_6184_2717.t1 a_6018_2717.t7 VDDD.t359 VDDD.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1391 VSSD.t304 a_7423_n9724.t7 a_7357_n9650.t0 VSSD.t303 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1392 a_8265_n9484.t0 a_8099_n9484.t6 VSSD.t25 VSSD.t24 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1393 VSSD.t694 EN.t80 a_2478_n4714.t0 VSSD.t693 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1394 a_995_n10028.t2 CLKS.t117 VDDD.t172 VDDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1395 a_6645_n4702.t0 a_5564_n5074.t7 a_6298_n5106.t0 VDDD.t759 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1396 a_3559_n9510.t1 a_3384_n9484.t5 a_3738_n9484.t0 VSSD.t465 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1397 VSSD.t617 auto_sampling_0.x22.A.t8 auto_sampling_0.x23.A.t0 VSSD.t616 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1398 a_8670_n1573.t1 a_8544_n1457.t4 a_8266_n1441.t2 VSSD.t667 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1399 SWP[0].t3 a_n8033_n9510.t6 VDDD.t1248 VDDD.t1247 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1400 a_3081_n9484.t0 a_3037_n9242.t5 a_2915_n9484.t0 VSSD.t538 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1401 a_2766_2717.t0 a_2320_2717.t5 a_2670_2717.t1 VSSD.t300 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1402 a_n5004_n9484.t1 cdac_ctrl_0.x1.X.t33 VSSD.t537 VSSD.t536 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1403 VDDD.t140 a_3692_n5650.t8 DOUT[4].t2 VDDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1404 a_3589_2717.t1 EN.t81 VSSD.t696 VSSD.t695 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1405 a_5113_n1207.t0 CLKS.t118 VSSD.t1033 VSSD.t1032 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1406 VSSD.t207 CKO.t21 a_7496_n5074.t0 VSSD.t206 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1407 VSSD.t990 a_4115_n1599.t7 CF[2].t1 VSSD.t989 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1408 a_n8208_n9484.t0 a_n9289_n9484.t7 a_n8555_n9242.t0 VDDD.t794 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1409 auto_sampling_0.x24.A.t5 auto_sampling_0.x23.A.t11 VDDD.t192 VDDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1410 VSSD.t1148 a_3559_n9510.t6 SWP[6].t0 VSSD.t79 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1411 VSSD.t653 SWP[6].t5 a_6947_n5258.t3 VSSD.t652 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1412 a_4383_n5258.t3 a_4296_n5482.t5 a_3979_n5372.t3 VDDD.t1374 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1413 a_n4169_n9510.t2 CLKS.t119 VDDD.t487 VDDD.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1414 auto_sampling_0.x12.D.t0 auto_sampling_0.x11.Q.t5 VSSD.t295 VSSD.t294 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1415 auto_sampling_0.x5.D.t2 a_5343_3531.t8 VDDD.t584 VDDD.t583 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1416 a_n454_2691.t2 a_n629_2717.t5 a_n275_2717.t1 VSSD.t381 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1417 VDDD.t22 a_n8033_n9724.t7 SWN[0].t2 VDDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1418 VDDD.t114 a_2889_3799.t5 a_2779_3923.t2 VDDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1419 a_5522_3557.t0 EN.t82 VSSD.t698 VSSD.t697 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1420 a_9661_n5596.t1 CLKS.t120 VSSD.t1029 VSSD.t1028 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1421 a_n7854_n9484.t1 CLKS.t121 VSSD.t1027 VSSD.t1026 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1422 VDDD.t670 CF[2].t8 a_3506_n1573.t2 VDDD.t669 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1423 VSSD.t27 a_n8033_n9724.t8 SWN[0].t0 VSSD.t26 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1424 a_958_n4702.t1 a_n232_n5074.t6 a_849_n4702.t3 VSSD.t954 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1425 auto_sampling_0.x7.Q.t3 a_n453_3531.t8 VDDD.t1354 VDDD.t1353 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1426 VDDD.t1383 a_n628_3557.t5 a_n453_3531.t2 VDDD.t1382 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1427 VDDD.t1026 CLK.t28 a_n1709_3557.t1 VDDD.t1025 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1428 CF[4].t3 a_7979_n1599.t7 VDDD.t965 VDDD.t964 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1429 VDDD.t1385 a_3559_n9510.t7 SWP[6].t2 VDDD.t1384 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1430 VDDD.t415 a_2956_n4776.t5 a_2943_n5080.t0 VDDD.t414 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1431 a_9355_n9510.t2 CLKS.t122 VDDD.t489 VDDD.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1432 a_n305_n9724.t2 CLKS.t123 VDDD.t491 VDDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1433 a_4969_n10054.t1 a_4751_n9650.t5 VDDD.t333 VDDD.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1434 VSSD.t595 a_2956_n4776.t6 DOUT[3].t1 VSSD.t594 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1435 VSSD.t84 CF[1].t7 a_1574_n1573.t2 VSSD.t83 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1436 out_latch_0.FINAL.t9 a_n784_n1599.t20 VDDD.t1447 VDDD.t1446 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1437 VSSD.t78 a_n4169_n9724.t8 a_n4235_n9650.t0 VSSD.t77 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1438 a_2321_3557.t0 a_2155_3557.t6 VSSD.t428 VSSD.t427 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1439 a_n4813_n9650.t0 a_n5259_n10022.t4 a_n4909_n9650.t3 VSSD.t614 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1440 VSSD.t354 a_n10393_n10028.t19 cdac_ctrl_0.x2.X.t13 VSSD.t248 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1441 a_5168_3557.t3 a_4253_3557.t5 a_4821_3799.t1 VSSD.t501 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1442 a_588_n5387.t2 a_393_n5356.t5 a_898_n5624.t0 VSSD.t746 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1443 VDDD.t1449 a_n784_n1599.t21 out_latch_0.FINAL.t8 VDDD.t1448 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1444 VSSD.t253 a_1760_n5650.t7 DOUT[2].t0 VSSD.t252 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X1445 a_6153_n1029.t0 a_5987_n1029.t7 VSSD.t683 VSSD.t682 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1446 VDDD.t984 CF[7].t8 a_4235_n9484.t1 VDDD.t983 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1447 a_n3990_n9662.t1 CLKS.t124 VSSD.t1025 VSSD.t1024 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1448 VDDD.t581 a_5316_n9650.t4 a_5491_n9724.t0 VDDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1449 VDDD.t1006 a_2787_n1331.t7 a_2748_n1457.t1 VDDD.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1450 a_739_3557.t1 a_223_3557.t6 a_644_3557.t1 VSSD.t643 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1451 a_2927_n10028.t2 a_2303_n10022.t5 a_2819_n9650.t1 VDDD.t1151 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1452 VDDD.t483 CLKS.t125 a_6952_n1573.t2 VDDD.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1453 a_5020_n1573.t2 a_4806_n1573.t4 VDDD.t1098 VDDD.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1454 a_5478_n9118.t1 a_4401_n9484.t5 a_5316_n9484.t2 VDDD.t1182 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1455 a_8266_n1441.t1 a_8583_n1331.t7 a_8541_n1207.t0 VSSD.t1004 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1456 a_1447_n1055.t1 a_1272_n1029.t5 a_1626_n1029.t0 VSSD.t953 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1457 a_6333_n9484.t0 a_6167_n9484.t6 VDDD.t1103 VDDD.t1102 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1458 a_5438_n1573.t0 a_4719_n1331.t6 a_4875_n1599.t1 VSSD.t234 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1459 VSSD.t1023 CLKS.t126 a_3081_n9484.t1 VSSD.t1022 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1460 VSSD.t1021 CLKS.t127 a_n783_n9484.t1 VSSD.t1020 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1461 a_6185_3557.t1 a_6019_3557.t6 VDDD.t354 VDDD.t353 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1462 a_5185_n1207.t1 a_4806_n1573.t5 a_5113_n1207.t1 VSSD.t864 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1463 VSSD.t161 auto_sampling_0.x24.A.t20 CLKS.t1 VSSD.t160 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1464 VDDD.t1132 CF[1].t8 a_n7357_n10022.t1 VDDD.t1131 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1465 a_2915_n9650.t1 a_2469_n10022.t5 a_2819_n9650.t2 VSSD.t444 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1466 a_n6623_n9242.t1 a_n6841_n9484.t5 VSSD.t405 VSSD.t404 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1467 a_9534_n9662.t1 CLKS.t128 VSSD.t1019 VSSD.t1018 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1468 a_5067_n4714.t0 EN.t83 VSSD.t1168 VSSD.t1167 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1469 VDDD.t1360 a_n2237_n9724.t7 a_n2250_n10028.t0 VDDD.t1359 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1470 VSSD.t581 a_7274_2691.t8 a_7208_2717.t1 VSSD.t580 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1471 a_8371_2717.t3 auto_sampling_0.x21.D.t5 VDDD.t128 VDDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1472 VSSD.t806 CLK.t29 a_7950_2717.t0 VSSD.t805 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1473 a_8615_n9650.t3 a_8265_n10022.t5 a_8520_n9662.t1 VDDD.t374 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1474 a_849_n4702.t1 a_n66_n5074.t5 a_502_n5106.t0 VSSD.t977 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1475 VDDD.t174 auto_sampling_0.x24.A.t21 CLKS.t2 VDDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1476 VSSD.t467 CLK.t30 a_222_2717.t0 VSSD.t466 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1477 VSSD.t469 CLK.t31 a_n1709_3557.t0 VSSD.t468 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1478 a_9141_3557.t0 a_7951_3557.t7 a_9032_3557.t1 VSSD.t948 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1479 VSSD.t963 CF[2].t9 a_n5425_n9484.t0 VSSD.t673 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1480 a_8577_n4702.t1 a_7496_n5074.t5 a_8230_n5106.t0 VDDD.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1481 a_n1045_n9484.t3 a_n1395_n9484.t5 a_n1140_n9484.t3 VDDD.t739 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1482 a_n4801_n10028.t2 a_n5425_n10022.t7 a_n4909_n9650.t0 VDDD.t775 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1483 VDDD.t1141 a_5624_n5650.t8 DOUT[6].t2 VDDD.t1140 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1484 a_7917_n4714.t0 SWP[9].t5 VSSD.t769 VSSD.t768 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1485 a_189_n4714.t2 SWP[1].t4 VSSD.t887 VSSD.t886 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1486 a_4864_2717.t1 a_4820_2959.t5 a_4698_2717.t1 VSSD.t741 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1487 a_6228_n5482.t0 CKO.t22 VSSD.t209 VSSD.t208 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1488 a_6820_n4776.t0 EN.t84 VDDD.t1407 VDDD.t1406 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1489 auto_sampling_0.x11.Q.t2 a_9207_3531.t8 VDDD.t232 VDDD.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1490 a_7045_n1207.t1 CLKS.t129 VSSD.t1017 VSSD.t1016 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1491 a_3410_2691.t1 a_3235_2717.t4 a_3589_2717.t0 VSSD.t529 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1492 a_8563_3557.t0 a_8117_3557.t5 a_8467_3557.t3 VSSD.t1135 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1493 VDDD.t566 CLK.t32 a_7950_2717.t1 VDDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1494 VSSD.t603 a_5491_n9510.t7 SWP[7].t0 VSSD.t602 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1495 CLKSB.t0 CLKS.t130 VSSD.t1015 VSSD.t1014 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1496 a_9031_2717.t1 a_7950_2717.t7 a_8684_2959.t0 VDDD.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1497 a_9386_3557.t0 EN.t85 VSSD.t1170 VSSD.t1169 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1498 VDDD.t568 CLK.t33 a_222_2717.t1 VDDD.t567 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1499 a_8723_n9118.t0 a_8099_n9484.t7 a_8615_n9484.t3 VDDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1500 a_502_n5106.t3 a_284_n4702.t5 VSSD.t710 VSSD.t709 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1501 a_4507_2717.t2 auto_sampling_0.x15.D.t5 VSSD.t688 VSSD.t687 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1502 VDDD.t1036 a_1627_n9724.t8 SWN[5].t2 VDDD.t1035 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1503 a_2469_n10022.t0 a_2303_n10022.t6 VSSD.t791 VSSD.t790 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1504 a_4366_n5106.t2 a_4148_n4702.t5 VDDD.t429 VDDD.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1505 SWN[3].t2 a_n2237_n9724.t8 VDDD.t1362 VDDD.t1361 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1506 a_9109_n1029.t0 a_7919_n1029.t6 a_9000_n1029.t3 VSSD.t969 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1507 a_9355_n9724.t2 CLKS.t131 VDDD.t464 VDDD.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1508 a_995_n9118.t1 CLKS.t132 VDDD.t466 VDDD.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1509 VDDD.t649 a_3235_2717.t5 a_3410_2691.t0 VDDD.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1510 a_8833_n10054.t2 a_8615_n9650.t5 VSSD.t345 VSSD.t344 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1511 VDDD.t120 a_8230_n5106.t5 a_8120_n5080.t2 VDDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1512 a_6188_n5080.t0 EN.t86 VDDD.t1409 VDDD.t1408 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1513 a_4221_n1029.t1 a_4055_n1029.t6 VDDD.t122 VDDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1514 VSSD.t1011 CLKS.t133 a_969_n1029.t1 VSSD.t1010 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1515 VSSD.t1009 CLKS.t134 a_5013_n9662.t1 VSSD.t1008 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1516 VDDD.t755 a_5491_n9510.t8 SWP[7].t2 VDDD.t754 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1517 VDDD.t496 a_4888_n4776.t8 a_4875_n5080.t0 VDDD.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1518 VDDD.t81 a_3559_n9724.t8 SWN[6].t2 VDDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1519 a_855_n1331.t0 CLK.t34 VSSD.t471 VSSD.t470 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1520 a_6185_3557.t0 a_6019_3557.t7 VSSD.t67 VSSD.t66 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1521 a_n8665_n10028.t2 CLKS.t135 VDDD.t1214 VDDD.t1213 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1522 a_n783_n9484.t0 a_n827_n9242.t5 a_n949_n9484.t0 VSSD.t272 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1523 VSSD.t721 a_n10393_n9484.t16 cdac_ctrl_0.x1.X.t2 VSSD.t351 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1524 VSSD.t473 CLK.t35 a_5987_n1029.t0 VSSD.t472 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1525 a_4679_n663.t0 a_4055_n1029.t7 a_4571_n1029.t3 VDDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1526 VDDD.t1411 EN.t87 a_7556_n5650.t0 VDDD.t1410 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1527 DOUT[2].t2 a_1760_n5650.t8 VDDD.t281 VDDD.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1528 VSSD.t47 a_1478_2691.t8 a_1412_2717.t0 VSSD.t46 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1529 a_2575_2717.t2 auto_sampling_0.x14.D.t5 VDDD.t1256 VDDD.t1255 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1530 VSSD.t475 CLK.t36 a_2154_2717.t0 VSSD.t474 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1531 a_n2412_n9484.t1 a_n3327_n9484.t5 a_n2759_n9242.t0 VSSD.t157 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1532 cdac_ctrl_0.x1.X.t1 a_n10393_n9484.t17 VSSD.t247 VSSD.t246 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1533 CF[1].t0 a_2183_n1599.t8 VSSD.t974 VSSD.t973 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1534 VDDD.t645 CF[8].t9 a_6167_n9484.t1 VDDD.t644 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1535 a_3345_3557.t0 a_2155_3557.t7 a_3236_3557.t1 VSSD.t429 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1536 a_2082_n5624.t1 a_2047_n5372.t5 a_1760_n5650.t2 VSSD.t940 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1537 VDDD.t992 a_n2412_n9484.t5 a_n2237_n9510.t1 VDDD.t991 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1538 a_3379_n1055.t1 a_3204_n1029.t5 a_3558_n1029.t0 VSSD.t901 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1539 VDDD.t1292 CF[3].t9 a_n3493_n9484.t1 VDDD.t1291 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1540 VDDD.t270 a_n10393_n9484.t18 cdac_ctrl_0.x1.X.t10 VDDD.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1541 a_7662_n5074.t1 a_7496_n5074.t6 VDDD.t884 VDDD.t883 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1542 a_2470_n1441.t3 a_2748_n1457.t5 a_2704_n1573.t1 VDDD.t837 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1543 auto_sampling_0.x3.D.t2 a_3411_3531.t8 VDDD.t1210 VDDD.t1209 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1544 a_4751_n9484.t1 a_4235_n9484.t7 a_4656_n9484.t0 VSSD.t150 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1545 a_n6745_n9484.t1 a_n7191_n9484.t5 a_n6841_n9484.t3 VSSD.t890 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1546 a_2767_3557.t1 a_2321_3557.t5 a_2671_3557.t3 VSSD.t956 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1547 VDDD.t339 CLK.t37 a_2154_2717.t1 VDDD.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1548 cdac_ctrl_0.x1.X.t9 a_n10393_n9484.t19 VDDD.t272 VDDD.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1549 VDDD.t606 a_6901_n10054.t5 a_6791_n10028.t1 VDDD.t605 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1550 CLKS.t3 auto_sampling_0.x24.A.t22 VSSD.t163 VSSD.t162 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1551 a_9180_n9484.t0 a_8265_n9484.t5 a_8833_n9242.t0 VSSD.t70 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1552 a_4847_n9650.t0 a_4401_n10022.t5 a_4751_n9650.t3 VSSD.t935 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1553 a_8316_n5387.t0 a_8121_n5356.t5 a_8626_n5624.t1 VSSD.t699 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1554 a_1561_n9484.t0 a_371_n9484.t6 a_1452_n9484.t0 VSSD.t601 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1555 DOUT[1].t0 a_1024_n4776.t8 VSSD.t314 VSSD.t313 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1556 a_n5259_n9484.t1 a_n5425_n9484.t7 VSSD.t658 VSSD.t424 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1557 VSSD.t597 a_2956_n4776.t7 a_2890_n4702.t1 VSSD.t596 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1558 a_537_n9484.t0 a_371_n9484.t7 VSSD.t29 VSSD.t28 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1559 a_3692_n5650.t2 a_3979_n5372.t5 VDDD.t744 VDDD.t743 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1560 a_1105_n10054.t1 a_887_n9650.t5 VSSD.t494 VSSD.t493 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1561 a_n1544_2717.t0 a_n1710_2717.t6 VSSD.t986 VSSD.t985 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1562 VDDD.t341 CLK.t38 a_7951_3557.t1 VDDD.t340 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1563 VDDD.t320 a_n6101_n9724.t7 SWN[1].t2 VDDD.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1564 VDDD.t343 CLK.t39 a_223_3557.t1 VDDD.t342 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1565 VSSD.t895 CF[1].t9 a_n7357_n9484.t1 VSSD.t81 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1566 VSSD.t766 a_6228_n5482.t7 a_6189_n5356.t1 VSSD.t765 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1567 a_n1289_2717.t2 auto_sampling_0.x12.D.t3 VSSD.t613 VSSD.t612 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1568 a_7274_2691.t0 a_7099_2717.t4 a_7453_2717.t1 VSSD.t627 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1569 VDDD.t155 a_n6623_n10054.t5 a_n6733_n10028.t2 VDDD.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1570 VSSD.t1146 CF[9].t9 a_8099_n10022.t1 VSSD.t256 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1571 VDDD.t1085 a_7243_n1055.t8 CF[6].t2 VDDD.t1084 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1572 a_2724_n9662.t2 cdac_ctrl_0.x2.X.t34 VDDD.t708 VDDD.t707 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1573 SWN[7].t0 a_5491_n9724.t8 VSSD.t755 VSSD.t564 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1574 a_4656_n9484.t3 cdac_ctrl_0.x1.X.t34 VDDD.t663 VDDD.t662 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1575 a_8012_n4702.t2 a_7496_n5074.t7 a_7917_n4714.t2 VSSD.t719 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1576 cdac_ctrl_0.x2.X.t14 a_n10393_n10028.t20 VSSD.t1193 VSSD.t191 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1577 a_284_n4702.t3 a_n232_n5074.t7 a_189_n4714.t1 VSSD.t955 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1578 a_8739_n1599.t2 a_8544_n1457.t5 a_9049_n1207.t0 VSSD.t668 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1579 VSSD.t251 a_3410_2691.t8 auto_sampling_0.x15.D.t0 VSSD.t250 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1580 a_n827_n9242.t1 a_n1045_n9484.t5 VDDD.t435 VDDD.t434 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1581 a_6080_n4702.t2 a_5730_n5074.t5 a_5985_n4714.t1 VDDD.t1401 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1582 a_5491_n9724.t1 a_5316_n9650.t5 a_5670_n9662.t0 VSSD.t243 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1583 a_n2303_n9484.t1 a_n3493_n9484.t6 a_n2412_n9484.t2 VSSD.t61 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1584 a_1024_n4776.t0 a_849_n4702.t5 a_1203_n4714.t0 VSSD.t764 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1585 VDDD.t656 a_9487_n4848.t4 CKO.t0 VDDD.t542 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1586 a_4822_n4702.t0 a_3632_n5074.t7 a_4713_n4702.t0 VSSD.t94 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1587 VDDD.t787 a_7099_2717.t5 a_7274_2691.t1 VDDD.t786 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1588 a_n1544_2717.t1 a_n1710_2717.t7 VDDD.t1286 VDDD.t1285 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1589 a_n937_n9118.t2 CLKS.t136 VDDD.t1216 VDDD.t1215 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1590 a_8085_n1029.t1 a_7919_n1029.t7 VDDD.t1260 VDDD.t1259 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1591 VDDD.t573 auto_sampling_0.x24.A.t23 CLKS.t11 VDDD.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1592 a_4710_3083.t0 EN.t88 VDDD.t1413 VDDD.t1412 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1593 a_3979_n5372.t0 a_4296_n5482.t6 a_4254_n5624.t1 VSSD.t394 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1594 VSSD.t154 a_n8033_n9510.t7 SWP[0].t0 VSSD.t26 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1595 a_6369_n1207.t0 a_6334_n1441.t5 a_6047_n1599.t0 VSSD.t96 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1596 VDDD.t481 COMP_N.t5 a_n10393_n10028.t5 VDDD.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1597 a_643_2717.t0 auto_sampling_0.x22.A.t9 VSSD.t619 VSSD.t618 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1598 a_2121_n4714.t1 SWP[3].t5 VDDD.t43 VDDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1599 a_n4182_n10028.t0 a_n5259_n10022.t5 a_n4344_n9650.t2 VDDD.t982 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1600 a_8120_n5080.t0 EN.t89 VDDD.t373 VDDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1601 a_4602_2717.t0 a_4086_2717.t7 a_4507_2717.t0 VSSD.t417 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1602 a_n8773_n9484.t1 a_n9123_n9484.t4 a_n8868_n9484.t1 VDDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1603 VDDD.t1046 a_6047_n1599.t8 CF[3].t2 VDDD.t1045 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1604 a_n8511_n9484.t0 a_n8555_n9242.t5 a_n8677_n9484.t1 VSSD.t320 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1605 a_5015_n5258.t2 a_4257_n5356.t5 a_4452_n5387.t1 VDDD.t875 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1606 a_1151_n5258.t0 a_432_n5482.t7 a_588_n5387.t0 VSSD.t994 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1607 VDDD.t1055 out_latch_0.FINAL.t19 a_9487_n4848.t1 VDDD.t945 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1608 a_n5004_n9484.t2 cdac_ctrl_0.x1.X.t35 VDDD.t37 VDDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1609 a_2787_n1331.t0 CLK.t40 VSSD.t306 VSSD.t305 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1610 VDDD.t1267 SWP[0].t5 a_1151_n5258.t3 VDDD.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1611 a_6408_n1029.t2 CF[7].t9 VSSD.t777 VSSD.t776 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1612 a_6683_n9484.t0 a_6333_n9484.t5 a_6588_n9484.t3 VDDD.t935 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1613 a_1452_n9484.t3 a_537_n9484.t5 a_1105_n9242.t3 VSSD.t95 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1614 a_n1045_n9650.t1 a_n1395_n10022.t5 a_n1140_n9662.t0 VDDD.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1615 a_n305_n9510.t2 CLKS.t137 VDDD.t1218 VDDD.t1217 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1616 VSSD.t249 a_n10393_n9484.t20 cdac_ctrl_0.x1.X.t0 VSSD.t248 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1617 VDDD.t161 a_n8033_n9510.t8 SWP[0].t2 VDDD.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1618 VDDD.t337 a_7423_n9724.t8 a_7410_n10028.t0 VDDD.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1619 a_8500_n1573.t1 a_7979_n1599.t8 VDDD.t967 VDDD.t966 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1620 a_9193_3083.t1 a_8116_2717.t5 a_9031_2717.t2 VDDD.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1621 cdac_ctrl_0.x2.X.t15 a_n10393_n10028.t21 VDDD.t1455 VDDD.t1454 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1622 a_2469_n10022.t1 a_2303_n10022.t7 VDDD.t1002 VDDD.t1001 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1623 CF[2].t0 a_4115_n1599.t8 VSSD.t992 VSSD.t991 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1624 VSSD.t1134 a_7275_3531.t8 a_7209_3557.t0 VSSD.t1133 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1625 VDDD.t345 CLK.t41 a_2155_3557.t0 VDDD.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1626 VSSD.t308 CLK.t42 a_7951_3557.t0 VSSD.t307 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1627 a_8723_n9118.t2 CLKS.t138 VDDD.t1220 VDDD.t1219 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1628 a_n3327_n9484.t1 a_n3493_n9484.t7 VDDD.t59 VDDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1629 VSSD.t310 CLK.t43 a_223_3557.t0 VSSD.t309 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1630 VSSD.t1177 CF[0].t12 a_n9289_n10022.t1 VSSD.t370 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1631 a_189_n4714.t3 SWP[1].t5 VDDD.t1125 VDDD.t1124 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1632 VDDD.t95 a_8739_n1599.t5 a_8670_n1573.t3 VDDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1633 a_5013_n9662.t0 a_4969_n10054.t5 a_4847_n9650.t1 VSSD.t926 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1634 VDDD.t1153 CKO.t23 a_7496_n5074.t1 VDDD.t1152 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1635 a_3204_n1029.t3 a_2123_n1029.t6 a_2857_n787.t3 VDDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1636 a_n6936_n9662.t1 cdac_ctrl_0.x2.X.t35 VSSD.t626 VSSD.t625 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1637 VSSD.t666 a_9175_n1055.t8 a_9109_n1029.t1 VSSD.t665 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1638 auto_sampling_0.x16.D.t2 a_5342_2691.t8 VDDD.t461 VDDD.t460 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1639 a_1478_2691.t1 a_1303_2717.t5 a_1657_2717.t1 VSSD.t1132 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1640 a_739_3557.t2 a_389_3557.t5 a_644_3557.t0 VDDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1641 VDDD.t1311 a_1447_n1055.t8 CF[9].t2 VDDD.t1310 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1642 VSSD.t1149 a_3559_n9510.t8 a_3493_n9484.t1 VSSD.t578 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1643 a_7248_n9484.t1 a_6167_n9484.t7 a_6901_n9242.t0 VDDD.t1104 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1644 VDDD.t411 a_n10393_n9484.t21 cdac_ctrl_0.x1.X.t8 VDDD.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1645 VDDD.t446 a_4296_n5482.t7 a_4257_n5356.t0 VDDD.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1646 a_4401_n10022.t1 a_4235_n10022.t7 VDDD.t275 VDDD.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1647 SWN[1].t0 a_n6101_n9724.t8 VSSD.t289 VSSD.t288 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1648 VDDD.t1421 CF[0].t13 a_n784_n1599.t5 VDDD.t1420 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1649 a_n8677_n9484.t0 a_n9123_n9484.t5 a_n8773_n9484.t2 VSSD.t135 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1650 a_9487_n5472.t2 CLKS.t139 VDDD.t1070 VDDD.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1651 a_1011_n1599.t1 a_816_n1457.t5 a_1321_n1207.t0 VSSD.t867 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1652 a_4865_3557.t1 a_4821_3799.t5 a_4699_3557.t1 VSSD.t700 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1653 VDDD.t1072 CLKS.t140 a_6047_n1599.t2 VDDD.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1654 a_3411_3531.t1 a_3236_3557.t5 a_3590_3557.t1 VSSD.t457 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1655 a_2943_n5080.t1 a_1866_n5074.t5 a_2781_n4702.t3 VDDD.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1656 a_n8033_n9510.t1 a_n8208_n9484.t5 a_n7854_n9484.t0 VSSD.t531 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1657 VDDD.t543 a_9487_n5472.t4 CKO.t3 VDDD.t542 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1658 a_4713_n4702.t3 a_3798_n5074.t5 a_4366_n5106.t3 VSSD.t738 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1659 a_n466_3923.t0 a_n1543_3557.t5 a_n628_3557.t0 VDDD.t582 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1660 a_n2869_n10028.t0 a_n3493_n10022.t7 a_n2977_n9650.t2 VDDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1661 VDDD.t932 a_7248_n9484.t5 a_7423_n9510.t0 VDDD.t931 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1662 a_2289_n1029.t1 a_2123_n1029.t7 VDDD.t31 VDDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1663 a_847_3923.t2 a_223_3557.t7 a_739_3557.t0 VDDD.t818 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1664 DOUT[3].t0 a_2956_n4776.t8 VSSD.t599 VSSD.t598 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X1665 a_4806_n1573.t0 a_4719_n1331.t7 a_4402_n1441.t0 VDDD.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1666 a_n126_n9662.t1 CLKS.t141 VSSD.t1007 VSSD.t1006 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1667 a_4508_3557.t1 auto_sampling_0.x3.D.t5 VSSD.t588 VSSD.t587 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1668 a_8653_n787.t1 a_8435_n1029.t5 VDDD.t455 VDDD.t454 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1669 VDDD.t1281 a_8684_2959.t5 a_8574_3083.t2 VDDD.t1280 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
R0 a_7068_n1029.n3 a_7068_n1029.n2 636.953
R1 a_7068_n1029.n1 a_7068_n1029.t5 366.856
R2 a_7068_n1029.n2 a_7068_n1029.n0 300.2
R3 a_7068_n1029.n2 a_7068_n1029.n1 225.036
R4 a_7068_n1029.n1 a_7068_n1029.t4 174.056
R5 a_7068_n1029.n0 a_7068_n1029.t3 70.0005
R6 a_7068_n1029.t0 a_7068_n1029.n3 68.0124
R7 a_7068_n1029.n3 a_7068_n1029.t2 63.3219
R8 a_7068_n1029.n0 a_7068_n1029.t1 61.6672
R9 a_7243_n1055.n5 a_7243_n1055.n4 807.871
R10 a_7243_n1055.n2 a_7243_n1055.t7 389.183
R11 a_7243_n1055.n3 a_7243_n1055.n2 251.167
R12 a_7243_n1055.n3 a_7243_n1055.t1 223.571
R13 a_7243_n1055.n0 a_7243_n1055.t8 212.081
R14 a_7243_n1055.n1 a_7243_n1055.t6 212.081
R15 a_7243_n1055.n4 a_7243_n1055.n1 176.576
R16 a_7243_n1055.n2 a_7243_n1055.t3 174.891
R17 a_7243_n1055.n0 a_7243_n1055.t5 139.78
R18 a_7243_n1055.n1 a_7243_n1055.t4 139.78
R19 a_7243_n1055.n5 a_7243_n1055.t2 63.3219
R20 a_7243_n1055.t0 a_7243_n1055.n5 63.3219
R21 a_7243_n1055.n1 a_7243_n1055.n0 61.346
R22 a_7243_n1055.n4 a_7243_n1055.n3 37.7195
R23 VDDD.n1874 VDDD.t130 877.144
R24 VDDD.n254 VDDD.t382 806.511
R25 VDDD.n345 VDDD.t459 806.511
R26 VDDD.n229 VDDD.t1074 806.511
R27 VDDD.n414 VDDD.t62 806.511
R28 VDDD.n204 VDDD.t435 806.511
R29 VDDD.n483 VDDD.t1067 806.511
R30 VDDD.n179 VDDD.t260 806.511
R31 VDDD.n552 VDDD.t1228 806.511
R32 VDDD.n154 VDDD.t1082 806.511
R33 VDDD.n621 VDDD.t1236 806.511
R34 VDDD.n129 VDDD.t1108 806.511
R35 VDDD.n688 VDDD.t1196 806.511
R36 VDDD.n104 VDDD.t333 806.511
R37 VDDD.n757 VDDD.t194 806.511
R38 VDDD.n79 VDDD.t595 806.511
R39 VDDD.n826 VDDD.t588 806.511
R40 VDDD.n54 VDDD.t28 806.511
R41 VDDD.n895 VDDD.t724 806.511
R42 VDDD.n29 VDDD.t1283 806.511
R43 VDDD.n964 VDDD.t846 806.511
R44 VDDD.n2455 VDDD.t689 806.511
R45 VDDD.n2198 VDDD.t331 806.511
R46 VDDD.n2212 VDDD.t351 806.511
R47 VDDD.n2226 VDDD.t704 806.511
R48 VDDD.n2240 VDDD.t683 806.511
R49 VDDD.n2254 VDDD.t421 806.511
R50 VDDD.n2159 VDDD.t549 806.511
R51 VDDD.n1906 VDDD.t443 806.511
R52 VDDD.n1920 VDDD.t1167 806.511
R53 VDDD.n1934 VDDD.t860 806.511
R54 VDDD.n1948 VDDD.t16 806.511
R55 VDDD.n1962 VDDD.t1170 806.511
R56 VDDD.n1383 VDDD.t95 806.511
R57 VDDD.n1397 VDDD.t1234 806.511
R58 VDDD.n1411 VDDD.t361 806.511
R59 VDDD.n1425 VDDD.t468 806.511
R60 VDDD.n1439 VDDD.t1327 806.511
R61 VDDD.n1813 VDDD.t457 806.511
R62 VDDD.n1327 VDDD.t882 806.511
R63 VDDD.n1341 VDDD.t214 806.511
R64 VDDD.n1355 VDDD.t518 806.511
R65 VDDD.n1369 VDDD.t455 806.511
R66 VDDD.n1132 VDDD.t570 806.511
R67 VDDD.n1134 VDDD.t41 806.511
R68 VDDD.n1169 VDDD.t1334 806.511
R69 VDDD.n1171 VDDD.t586 806.511
R70 VDDD.n1206 VDDD.t429 806.511
R71 VDDD.n1208 VDDD.t763 806.511
R72 VDDD.n1243 VDDD.t1016 806.511
R73 VDDD.n1245 VDDD.t165 806.511
R74 VDDD.n1015 VDDD.t878 806.511
R75 VDDD.n1284 VDDD.t1377 806.511
R76 VDDD.t19 VDDD.t1450 790.188
R77 VDDD.t1102 VDDD.t97 790.188
R78 VDDD.t152 VDDD.t662 790.188
R79 VDDD.t209 VDDD.t237 790.188
R80 VDDD.t1403 VDDD.t416 790.188
R81 VDDD.t760 VDDD.t99 790.188
R82 VDDD.t58 VDDD.t235 790.188
R83 VDDD.t833 VDDD.t36 790.188
R84 VDDD.t806 VDDD.t660 790.188
R85 VDDD.t125 VDDD.t1452 790.188
R86 VDDD.t127 VDDD.t249 790.188
R87 VDDD.t1342 VDDD.t358 790.188
R88 VDDD.t865 VDDD.t510 790.188
R89 VDDD.t1255 VDDD.t843 790.188
R90 VDDD.t621 VDDD.t394 790.188
R91 VDDD.t505 VDDD.t1285 790.188
R92 VDDD.t375 VDDD.t1205 790.188
R93 VDDD.t816 VDDD.t353 790.188
R94 VDDD.t733 VDDD.t856 790.188
R95 VDDD.t995 VDDD.t658 790.188
R96 VDDD.t729 VDDD.t973 790.188
R97 VDDD.t1432 VDDD.t1161 790.188
R98 VDDD.t440 VDDD.t533 790.188
R99 VDDD.t1425 VDDD.t0 790.188
R100 VDDD.t245 VDDD.t1289 790.188
R101 VDDD.t1005 VDDD.t669 790.188
R102 VDDD.t596 VDDD.t82 790.188
R103 VDDD.t133 VDDD.t1259 790.188
R104 VDDD.t239 VDDD.t367 790.188
R105 VDDD.t642 VDDD.t121 790.188
R106 VDDD.t1380 VDDD.t30 790.188
R107 VDDD.t1203 VDDD.t364 790.188
R108 VDDD.t948 VDDD.t1037 790.188
R109 VDDD.t1174 VDDD.t705 790.188
R110 VDDD.t274 VDDD.t1120 790.188
R111 VDDD.t1001 VDDD.t707 790.188
R112 VDDD.t752 VDDD.t1122 790.188
R113 VDDD.t308 VDDD.t1118 790.188
R114 VDDD.t591 VDDD.t1039 790.188
R115 VDDD.t773 VDDD.t1185 790.188
R116 VDDD.t6 VDDD.t1041 790.188
R117 VDDD.t922 VDDD.t1183 790.188
R118 VDDD.n1105 VDDD.t1055 675.293
R119 VDDD.n1105 VDDD.t946 675.293
R120 VDDD.n300 VDDD.t1453 667.778
R121 VDDD.n334 VDDD.t661 667.778
R122 VDDD.n369 VDDD.t37 667.778
R123 VDDD.n403 VDDD.t236 667.778
R124 VDDD.n438 VDDD.t100 667.778
R125 VDDD.n472 VDDD.t417 667.778
R126 VDDD.n507 VDDD.t238 667.778
R127 VDDD.n541 VDDD.t663 667.778
R128 VDDD.n576 VDDD.t98 667.778
R129 VDDD.n610 VDDD.t1451 667.778
R130 VDDD.n664 VDDD.t1038 667.778
R131 VDDD.n699 VDDD.t706 667.778
R132 VDDD.n733 VDDD.t1121 667.778
R133 VDDD.n768 VDDD.t708 667.778
R134 VDDD.n802 VDDD.t1123 667.778
R135 VDDD.n837 VDDD.t1119 667.778
R136 VDDD.n871 VDDD.t1040 667.778
R137 VDDD.n906 VDDD.t1186 667.778
R138 VDDD.n940 VDDD.t1042 667.778
R139 VDDD.n975 VDDD.t1184 667.778
R140 VDDD.n2180 VDDD.t1433 667.778
R141 VDDD.n2433 VDDD.t730 667.778
R142 VDDD.n2400 VDDD.t996 667.778
R143 VDDD.n2367 VDDD.t734 667.778
R144 VDDD.n2334 VDDD.t817 667.778
R145 VDDD.n2301 VDDD.t376 667.778
R146 VDDD.n1888 VDDD.t506 667.778
R147 VDDD.n2137 VDDD.t622 667.778
R148 VDDD.n2104 VDDD.t1256 667.778
R149 VDDD.n2071 VDDD.t866 667.778
R150 VDDD.n2038 VDDD.t1343 667.778
R151 VDDD.n2005 VDDD.t128 667.778
R152 VDDD.n1634 VDDD.t534 667.778
R153 VDDD.n1601 VDDD.t1 667.778
R154 VDDD.n1568 VDDD.t1290 667.778
R155 VDDD.n1535 VDDD.t670 667.778
R156 VDDD.n1502 VDDD.t83 667.778
R157 VDDD.n1309 VDDD.t1204 667.778
R158 VDDD.n1791 VDDD.t1381 667.778
R159 VDDD.n1758 VDDD.t643 667.778
R160 VDDD.n1725 VDDD.t240 667.778
R161 VDDD.n1692 VDDD.t134 667.778
R162 VDDD.n321 VDDD.t289 667.751
R163 VDDD.n237 VDDD.t1458 667.751
R164 VDDD.n390 VDDD.t1155 667.751
R165 VDDD.n212 VDDD.t992 667.751
R166 VDDD.n459 VDDD.t551 667.751
R167 VDDD.n187 VDDD.t1160 667.751
R168 VDDD.n528 VDDD.t563 667.751
R169 VDDD.n162 VDDD.t256 667.751
R170 VDDD.n597 VDDD.t932 667.751
R171 VDDD.n138 VDDD.t1111 667.751
R172 VDDD.n643 VDDD.t692 667.751
R173 VDDD.n677 VDDD.t732 667.751
R174 VDDD.n712 VDDD.t581 667.751
R175 VDDD.n746 VDDD.t604 667.751
R176 VDDD.n781 VDDD.t64 667.751
R177 VDDD.n815 VDDD.t302 667.751
R178 VDDD.n850 VDDD.t737 667.751
R179 VDDD.n884 VDDD.t696 667.751
R180 VDDD.n919 VDDD.t1137 667.751
R181 VDDD.n953 VDDD.t75 667.751
R182 VDDD.n2188 VDDD.t1383 667.751
R183 VDDD.n2413 VDDD.t609 667.751
R184 VDDD.n2380 VDDD.t451 667.751
R185 VDDD.n2347 VDDD.t961 667.751
R186 VDDD.n2314 VDDD.t102 667.751
R187 VDDD.n2281 VDDD.t439 667.751
R188 VDDD.n1896 VDDD.t433 667.751
R189 VDDD.n2117 VDDD.t1258 667.751
R190 VDDD.n2084 VDDD.t649 667.751
R191 VDDD.n2051 VDDD.t327 667.751
R192 VDDD.n2018 VDDD.t787 667.751
R193 VDDD.n1985 VDDD.t685 667.751
R194 VDDD.n1614 VDDD.t1397 667.751
R195 VDDD.n1581 VDDD.t800 667.751
R196 VDDD.n1548 VDDD.t1296 667.751
R197 VDDD.n1515 VDDD.t222 667.751
R198 VDDD.n1482 VDDD.t476 667.751
R199 VDDD.n1317 VDDD.t1212 667.751
R200 VDDD.n1771 VDDD.t1135 667.751
R201 VDDD.n1738 VDDD.t1106 667.751
R202 VDDD.n1705 VDDD.t1069 667.751
R203 VDDD.n1672 VDDD.t1240 667.751
R204 VDDD.n1121 VDDD.t254 664.455
R205 VDDD.n1145 VDDD.t163 664.455
R206 VDDD.n1158 VDDD.t393 664.455
R207 VDDD.n1182 VDDD.t228 664.455
R208 VDDD.n1195 VDDD.t1078 664.455
R209 VDDD.n1219 VDDD.t744 664.455
R210 VDDD.n1232 VDDD.t1294 664.455
R211 VDDD.n1256 VDDD.t1194 664.455
R212 VDDD.n1269 VDDD.t954 664.455
R213 VDDD.n1294 VDDD.t789 664.455
R214 VDDD.n1122 VDDD.t1222 663.426
R215 VDDD.n1144 VDDD.t959 663.426
R216 VDDD.n1159 VDDD.t832 663.426
R217 VDDD.n1181 VDDD.t1279 663.426
R218 VDDD.n1196 VDDD.t112 663.426
R219 VDDD.n1218 VDDD.t796 663.426
R220 VDDD.n1233 VDDD.t1389 663.426
R221 VDDD.n1255 VDDD.t43 663.426
R222 VDDD.n1270 VDDD.t1267 663.426
R223 VDDD.n1295 VDDD.t1125 663.426
R224 VDDD.t1110 VDDD.t1371 636.293
R225 VDDD.t931 VDDD.t1144 636.293
R226 VDDD.t255 VDDD.t699 636.293
R227 VDDD.t562 VDDD.t34 636.293
R228 VDDD.t1159 VDDD.t1011 636.293
R229 VDDD.t550 VDDD.t217 636.293
R230 VDDD.t991 VDDD.t90 636.293
R231 VDDD.t1154 VDDD.t1335 636.293
R232 VDDD.t1457 VDDD.t861 636.293
R233 VDDD.t288 VDDD.t1247 636.293
R234 VDDD.t403 VDDD.t684 636.293
R235 VDDD.t52 VDDD.t786 636.293
R236 VDDD.t460 VDDD.t326 636.293
R237 VDDD.t1029 VDDD.t648 636.293
R238 VDDD.t50 VDDD.t1257 636.293
R239 VDDD.t195 VDDD.t432 636.293
R240 VDDD.t231 VDDD.t438 636.293
R241 VDDD.t103 VDDD.t101 636.293
R242 VDDD.t583 VDDD.t960 636.293
R243 VDDD.t1209 VDDD.t450 636.293
R244 VDDD.t554 VDDD.t608 636.293
R245 VDDD.t1353 VDDD.t1382 636.293
R246 VDDD.t1396 VDDD.t962 636.293
R247 VDDD.t799 VDDD.t1045 636.293
R248 VDDD.t1295 VDDD.t1249 636.293
R249 VDDD.t221 VDDD.t1261 636.293
R250 VDDD.t475 VDDD.t88 636.293
R251 VDDD.t1229 VDDD.t1239 636.293
R252 VDDD.t1088 VDDD.t1068 636.293
R253 VDDD.t680 VDDD.t1105 636.293
R254 VDDD.t1365 VDDD.t1134 636.293
R255 VDDD.t229 VDDD.t1211 636.293
R256 VDDD.t691 VDDD.t117 636.293
R257 VDDD.t731 VDDD.t1386 636.293
R258 VDDD.t580 VDDD.t715 636.293
R259 VDDD.t603 VDDD.t770 636.293
R260 VDDD.t63 VDDD.t1031 636.293
R261 VDDD.t301 VDDD.t146 636.293
R262 VDDD.t736 VDDD.t1361 636.293
R263 VDDD.t695 VDDD.t78 636.293
R264 VDDD.t1136 VDDD.t317 636.293
R265 VDDD.t74 VDDD.t599 636.293
R266 VDDD.n1662 VDDD.t321 632.914
R267 VDDD.n252 VDDD.n251 604.457
R268 VDDD.n352 VDDD.n351 604.457
R269 VDDD.n227 VDDD.n226 604.457
R270 VDDD.n421 VDDD.n420 604.457
R271 VDDD.n202 VDDD.n201 604.457
R272 VDDD.n490 VDDD.n489 604.457
R273 VDDD.n177 VDDD.n176 604.457
R274 VDDD.n559 VDDD.n558 604.457
R275 VDDD.n152 VDDD.n151 604.457
R276 VDDD.n628 VDDD.n627 604.457
R277 VDDD.n132 VDDD.n131 604.457
R278 VDDD.n682 VDDD.n121 604.457
R279 VDDD.n107 VDDD.n106 604.457
R280 VDDD.n751 VDDD.n96 604.457
R281 VDDD.n82 VDDD.n81 604.457
R282 VDDD.n820 VDDD.n71 604.457
R283 VDDD.n57 VDDD.n56 604.457
R284 VDDD.n889 VDDD.n46 604.457
R285 VDDD.n32 VDDD.n31 604.457
R286 VDDD.n958 VDDD.n21 604.457
R287 VDDD.n2449 VDDD.n2187 604.457
R288 VDDD.n2201 VDDD.n2200 604.457
R289 VDDD.n2215 VDDD.n2214 604.457
R290 VDDD.n2229 VDDD.n2228 604.457
R291 VDDD.n2243 VDDD.n2242 604.457
R292 VDDD.n2257 VDDD.n2256 604.457
R293 VDDD.n2153 VDDD.n1895 604.457
R294 VDDD.n1909 VDDD.n1908 604.457
R295 VDDD.n1923 VDDD.n1922 604.457
R296 VDDD.n1937 VDDD.n1936 604.457
R297 VDDD.n1951 VDDD.n1950 604.457
R298 VDDD.n1965 VDDD.n1964 604.457
R299 VDDD.n1386 VDDD.n1385 604.457
R300 VDDD.n1400 VDDD.n1399 604.457
R301 VDDD.n1414 VDDD.n1413 604.457
R302 VDDD.n1428 VDDD.n1427 604.457
R303 VDDD.n1442 VDDD.n1441 604.457
R304 VDDD.n1807 VDDD.n1316 604.457
R305 VDDD.n1330 VDDD.n1329 604.457
R306 VDDD.n1344 VDDD.n1343 604.457
R307 VDDD.n1358 VDDD.n1357 604.457
R308 VDDD.n1372 VDDD.n1371 604.457
R309 VDDD.n1086 VDDD.n1085 604.457
R310 VDDD.n1077 VDDD.n1076 604.457
R311 VDDD.n1069 VDDD.n1068 604.457
R312 VDDD.n1060 VDDD.n1059 604.457
R313 VDDD.n1052 VDDD.n1051 604.457
R314 VDDD.n1043 VDDD.n1042 604.457
R315 VDDD.n1035 VDDD.n1034 604.457
R316 VDDD.n1026 VDDD.n1025 604.457
R317 VDDD.n1018 VDDD.n1017 604.457
R318 VDDD.n1293 VDDD.n1292 604.457
R319 VDDD.n295 VDDD.n294 604.394
R320 VDDD.n248 VDDD.n247 604.394
R321 VDDD.n364 VDDD.n363 604.394
R322 VDDD.n223 VDDD.n222 604.394
R323 VDDD.n433 VDDD.n432 604.394
R324 VDDD.n198 VDDD.n197 604.394
R325 VDDD.n502 VDDD.n501 604.394
R326 VDDD.n173 VDDD.n172 604.394
R327 VDDD.n571 VDDD.n570 604.394
R328 VDDD.n148 VDDD.n147 604.394
R329 VDDD.n670 VDDD.n669 604.394
R330 VDDD.n111 VDDD.n110 604.394
R331 VDDD.n739 VDDD.n738 604.394
R332 VDDD.n86 VDDD.n85 604.394
R333 VDDD.n808 VDDD.n807 604.394
R334 VDDD.n61 VDDD.n60 604.394
R335 VDDD.n877 VDDD.n876 604.394
R336 VDDD.n36 VDDD.n35 604.394
R337 VDDD.n946 VDDD.n945 604.394
R338 VDDD.n11 VDDD.n10 604.394
R339 VDDD.n2471 VDDD.n2179 604.394
R340 VDDD.n2438 VDDD.n2192 604.394
R341 VDDD.n2405 VDDD.n2206 604.394
R342 VDDD.n2372 VDDD.n2220 604.394
R343 VDDD.n2339 VDDD.n2234 604.394
R344 VDDD.n2306 VDDD.n2248 604.394
R345 VDDD.n2175 VDDD.n1887 604.394
R346 VDDD.n2142 VDDD.n1900 604.394
R347 VDDD.n2109 VDDD.n1914 604.394
R348 VDDD.n2076 VDDD.n1928 604.394
R349 VDDD.n2043 VDDD.n1942 604.394
R350 VDDD.n2010 VDDD.n1956 604.394
R351 VDDD.n1639 VDDD.n1376 604.394
R352 VDDD.n1606 VDDD.n1390 604.394
R353 VDDD.n1573 VDDD.n1404 604.394
R354 VDDD.n1540 VDDD.n1418 604.394
R355 VDDD.n1507 VDDD.n1432 604.394
R356 VDDD.n1829 VDDD.n1308 604.394
R357 VDDD.n1796 VDDD.n1321 604.394
R358 VDDD.n1763 VDDD.n1335 604.394
R359 VDDD.n1730 VDDD.n1349 604.394
R360 VDDD.n1697 VDDD.n1363 604.394
R361 VDDD.n1301 VDDD.n1010 604.394
R362 VDDD.n1089 VDDD.n1088 604.394
R363 VDDD.n1074 VDDD.n1073 604.394
R364 VDDD.n1072 VDDD.n1071 604.394
R365 VDDD.n1057 VDDD.n1056 604.394
R366 VDDD.n1055 VDDD.n1054 604.394
R367 VDDD.n1040 VDDD.n1039 604.394
R368 VDDD.n1038 VDDD.n1037 604.394
R369 VDDD.n1023 VDDD.n1022 604.394
R370 VDDD.n1021 VDDD.n1020 604.394
R371 VDDD.n308 VDDD.n307 601.679
R372 VDDD.n244 VDDD.n243 601.679
R373 VDDD.n377 VDDD.n376 601.679
R374 VDDD.n219 VDDD.n218 601.679
R375 VDDD.n446 VDDD.n445 601.679
R376 VDDD.n194 VDDD.n193 601.679
R377 VDDD.n515 VDDD.n514 601.679
R378 VDDD.n169 VDDD.n168 601.679
R379 VDDD.n584 VDDD.n583 601.679
R380 VDDD.n144 VDDD.n143 601.679
R381 VDDD.n657 VDDD.n656 601.679
R382 VDDD.n116 VDDD.n115 601.679
R383 VDDD.n726 VDDD.n725 601.679
R384 VDDD.n91 VDDD.n90 601.679
R385 VDDD.n795 VDDD.n794 601.679
R386 VDDD.n66 VDDD.n65 601.679
R387 VDDD.n864 VDDD.n863 601.679
R388 VDDD.n41 VDDD.n40 601.679
R389 VDDD.n933 VDDD.n932 601.679
R390 VDDD.n16 VDDD.n15 601.679
R391 VDDD.n2458 VDDD.n2457 601.679
R392 VDDD.n2426 VDDD.n2197 601.679
R393 VDDD.n2393 VDDD.n2211 601.679
R394 VDDD.n2360 VDDD.n2225 601.679
R395 VDDD.n2327 VDDD.n2239 601.679
R396 VDDD.n2294 VDDD.n2253 601.679
R397 VDDD.n2162 VDDD.n2161 601.679
R398 VDDD.n2130 VDDD.n1905 601.679
R399 VDDD.n2097 VDDD.n1919 601.679
R400 VDDD.n2064 VDDD.n1933 601.679
R401 VDDD.n2031 VDDD.n1947 601.679
R402 VDDD.n1998 VDDD.n1961 601.679
R403 VDDD.n1627 VDDD.n1382 601.679
R404 VDDD.n1594 VDDD.n1396 601.679
R405 VDDD.n1561 VDDD.n1410 601.679
R406 VDDD.n1528 VDDD.n1424 601.679
R407 VDDD.n1495 VDDD.n1438 601.679
R408 VDDD.n1816 VDDD.n1815 601.679
R409 VDDD.n1784 VDDD.n1326 601.679
R410 VDDD.n1751 VDDD.n1340 601.679
R411 VDDD.n1718 VDDD.n1354 601.679
R412 VDDD.n1685 VDDD.n1368 601.679
R413 VDDD.n1083 VDDD.n1082 601.679
R414 VDDD.n1080 VDDD.n1079 601.679
R415 VDDD.n1066 VDDD.n1065 601.679
R416 VDDD.n1063 VDDD.n1062 601.679
R417 VDDD.n1049 VDDD.n1048 601.679
R418 VDDD.n1046 VDDD.n1045 601.679
R419 VDDD.n1032 VDDD.n1031 601.679
R420 VDDD.n1029 VDDD.n1028 601.679
R421 VDDD.n1278 VDDD.n1277 601.679
R422 VDDD.n1286 VDDD.n1285 601.679
R423 VDDD.t269 VDDD 588.942
R424 VDDD.t384 VDDD 588.942
R425 VDDD.t1219 VDDD.t1235 583.023
R426 VDDD.t615 VDDD.t1081 583.023
R427 VDDD.t500 VDDD.t1227 583.023
R428 VDDD.t823 VDDD.t259 583.023
R429 VDDD.t465 VDDD.t1066 583.023
R430 VDDD.t1215 VDDD.t434 583.023
R431 VDDD.t1316 VDDD.t61 583.023
R432 VDDD.t899 VDDD.t1073 583.023
R433 VDDD.t903 VDDD.t458 583.023
R434 VDDD.t630 VDDD.t381 583.023
R435 VDDD.t1169 VDDD.t1322 583.023
R436 VDDD.t15 VDDD.t12 583.023
R437 VDDD.t859 VDDD.t1412 583.023
R438 VDDD.t1166 VDDD.t10 583.023
R439 VDDD.t442 VDDD.t1414 583.023
R440 VDDD.t548 VDDD.t868 583.023
R441 VDDD.t420 VDDD.t776 583.023
R442 VDDD.t682 VDDD.t624 583.023
R443 VDDD.t703 VDDD.t1346 583.023
R444 VDDD.t350 VDDD.t780 583.023
R445 VDDD.t330 VDDD.t1064 583.023
R446 VDDD.t688 VDDD.t181 583.023
R447 VDDD.t265 VDDD.t94 583.023
R448 VDDD.t482 VDDD.t1233 583.023
R449 VDDD.t313 VDDD.t360 583.023
R450 VDDD.t1270 VDDD.t467 583.023
R451 VDDD.t821 VDDD.t1326 583.023
R452 VDDD.t454 VDDD.t907 583.023
R453 VDDD.t517 VDDD.t1302 583.023
R454 VDDD.t213 VDDD.t544 583.023
R455 VDDD.t881 VDDD.t1300 583.023
R456 VDDD.t456 VDDD.t636 583.023
R457 VDDD.t905 VDDD.t1107 583.023
R458 VDDD.t1304 VDDD.t1195 583.023
R459 VDDD.t613 VDDD.t332 583.023
R460 VDDD.t1312 VDDD.t193 583.023
R461 VDDD.t171 VDDD.t594 583.023
R462 VDDD.t634 VDDD.t587 583.023
R463 VDDD.t546 VDDD.t27 583.023
R464 VDDD.t263 VDDD.t723 583.023
R465 VDDD.t901 VDDD.t1282 583.023
R466 VDDD.t1213 VDDD.t845 583.023
R467 VDDD.n2268 VDDD.t323 529.751
R468 VDDD.n1649 VDDD 521.697
R469 VDDD.t964 VDDD 488.318
R470 VDDD.t1075 VDDD 488.318
R471 VDDD.t1251 VDDD 488.318
R472 VDDD.t1331 VDDD 488.318
R473 VDDD.t86 VDDD 488.318
R474 VDDD.t1430 VDDD 420.25
R475 VDDD.t109 VDDD.t540 414.33
R476 VDDD.t1297 VDDD.t611 414.33
R477 VDDD.t151 VDDD.t1298 414.33
R478 VDDD.t1080 VDDD.t835 414.33
R479 VDDD.t1402 VDDD.t1337 414.33
R480 VDDD.t1394 VDDD.t889 414.33
R481 VDDD.t1277 VDDD.t529 414.33
R482 VDDD.t1158 VDDD.t797 414.33
R483 VDDD.t804 VDDD.t1378 414.33
R484 VDDD.t793 VDDD.t1237 414.33
R485 VDDD.n1976 VDDD.t407 414.33
R486 VDDD.t1280 VDDD.t248 414.33
R487 VDDD.t560 VDDD.t357 414.33
R488 VDDD.t919 VDDD.t512 414.33
R489 VDDD.t418 VDDD.t447 414.33
R490 VDDD.t558 VDDD.t772 414.33
R491 VDDD.t673 VDDD.t1171 414.33
R492 VDDD.t135 VDDD.t1330 414.33
R493 VDDD.t646 VDDD.t352 414.33
R494 VDDD.t870 VDDD.t855 414.33
R495 VDDD.t113 VDDD.t657 414.33
R496 VDDD.t709 VDDD.t818 414.33
R497 VDDD.t508 VDDD.t1133 414.33
R498 VDDD.t1328 VDDD.t328 414.33
R499 VDDD.t1427 VDDD.t650 414.33
R500 VDDD.t1263 VDDD.t1097 414.33
R501 VDDD.t362 VDDD.t640 414.33
R502 VDDD.t598 VDDD.t879 414.33
R503 VDDD.t448 VDDD.t504 414.33
R504 VDDD.t1180 VDDD.t369 414.33
R505 VDDD.t257 VDDD.t123 414.33
R506 VDDD.t452 VDDD.t791 414.33
R507 VDDD.t1027 VDDD.t26 414.33
R508 VDDD.t947 VDDD.t1355 414.33
R509 VDDD.t1173 VDDD.t605 414.33
R510 VDDD.t273 VDDD.t808 414.33
R511 VDDD.t1151 VDDD.t999 414.33
R512 VDDD.t750 VDDD.t141 414.33
R513 VDDD.t307 VDDD.t298 414.33
R514 VDDD.t57 VDDD.t745 414.33
R515 VDDD.t775 VDDD.t686 414.33
R516 VDDD.t639 VDDD.t154 414.33
R517 VDDD.t1165 VDDD.t355 414.33
R518 VDDD.n1006 VDDD 413.58
R519 VDDD.t129 VDDD 393.615
R520 VDDD.t1146 VDDD 387.695
R521 VDDD.t754 VDDD 387.695
R522 VDDD.t1384 VDDD 387.695
R523 VDDD.t1423 VDDD 387.695
R524 VDDD.t219 VDDD 387.695
R525 VDDD.t92 VDDD 387.695
R526 VDDD.t1349 VDDD 387.695
R527 VDDD.t748 VDDD 387.695
R528 VDDD.t160 VDDD 387.695
R529 VDDD VDDD.t727 387.695
R530 VDDD VDDD.t158 387.695
R531 VDDD VDDD.t278 387.695
R532 VDDD VDDD.t48 387.695
R533 VDDD VDDD.t197 387.695
R534 VDDD VDDD.t527 387.695
R535 VDDD VDDD.t107 387.695
R536 VDDD VDDD.t936 387.695
R537 VDDD VDDD.t989 387.695
R538 VDDD VDDD.t552 387.695
R539 VDDD VDDD.t1351 387.695
R540 VDDD VDDD.t1084 387.695
R541 VDDD VDDD.t678 387.695
R542 VDDD VDDD.t377 387.695
R543 VDDD VDDD.t1310 387.695
R544 VDDD.t334 VDDD 387.695
R545 VDDD.t713 VDDD 387.695
R546 VDDD.t80 VDDD 387.695
R547 VDDD.t1035 VDDD 387.695
R548 VDDD.t183 VDDD 387.695
R549 VDDD.t1357 VDDD 387.695
R550 VDDD.t863 VDDD 387.695
R551 VDDD.t319 VDDD 387.695
R552 VDDD.t21 VDDD 387.695
R553 VDDD.n1835 VDDD 379.039
R554 VDDD.t619 VDDD 369.938
R555 VDDD.n1836 VDDD.n1832 363.529
R556 VDDD.n1839 VDDD.n1832 363.529
R557 VDDD.n1837 VDDD.n1836 363.529
R558 VDDD.n1977 VDDD.n1970 363.529
R559 VDDD.n1973 VDDD.n1972 363.529
R560 VDDD.n1977 VDDD.n1972 363.529
R561 VDDD.n2269 VDDD.n2262 363.529
R562 VDDD.n2265 VDDD.n2264 363.529
R563 VDDD.n2269 VDDD.n2264 363.529
R564 VDDD.n1650 VDDD.n1643 363.529
R565 VDDD.n1650 VDDD.n1645 363.529
R566 VDDD.n1646 VDDD.n1645 363.529
R567 VDDD.n1663 VDDD.n1656 363.529
R568 VDDD.n1663 VDDD.n1658 363.529
R569 VDDD.n1659 VDDD.n1658 363.529
R570 VDDD.n1097 VDDD.n1094 363.529
R571 VDDD.n1100 VDDD.n1094 363.529
R572 VDDD.n1097 VDDD.n1095 363.529
R573 VDDD.t578 VDDD.t253 360.866
R574 VDDD.t162 VDDD.t520 360.866
R575 VDDD.t654 VDDD.t392 360.866
R576 VDDD.t227 VDDD.t1140 360.866
R577 VDDD.t1243 VDDD.t1077 360.866
R578 VDDD.t743 VDDD.t139 360.866
R579 VDDD.t412 VDDD.t1293 360.866
R580 VDDD.t1193 VDDD.t719 360.866
R581 VDDD.t346 VDDD.t953 360.866
R582 VDDD.t788 VDDD.t814 360.866
R583 VDDD.n323 VDDD.t1248 343.579
R584 VDDD.n357 VDDD.t862 343.579
R585 VDDD.n392 VDDD.t1336 343.579
R586 VDDD.n426 VDDD.t91 343.579
R587 VDDD.n461 VDDD.t218 343.579
R588 VDDD.n495 VDDD.t1012 343.579
R589 VDDD.n530 VDDD.t35 343.579
R590 VDDD.n564 VDDD.t700 343.579
R591 VDDD.n599 VDDD.t1145 343.579
R592 VDDD.n633 VDDD.t1372 343.579
R593 VDDD.n2444 VDDD.t1354 343.579
R594 VDDD.n2411 VDDD.t555 343.579
R595 VDDD.n2378 VDDD.t1210 343.579
R596 VDDD.n2345 VDDD.t584 343.579
R597 VDDD.n2312 VDDD.t104 343.579
R598 VDDD.n2279 VDDD.t232 343.579
R599 VDDD.n2148 VDDD.t196 343.579
R600 VDDD.n2115 VDDD.t51 343.579
R601 VDDD.n2082 VDDD.t1030 343.579
R602 VDDD.n2049 VDDD.t461 343.579
R603 VDDD.n2016 VDDD.t53 343.579
R604 VDDD.n1983 VDDD.t404 343.579
R605 VDDD.n1802 VDDD.t230 343.579
R606 VDDD.n1769 VDDD.t1366 343.579
R607 VDDD.n1736 VDDD.t681 343.579
R608 VDDD.n1703 VDDD.t1089 343.579
R609 VDDD.n1670 VDDD.t1230 343.579
R610 VDDD.n1147 VDDD.t521 343.579
R611 VDDD.n1184 VDDD.t1141 343.579
R612 VDDD.n1221 VDDD.t140 343.579
R613 VDDD.n1258 VDDD.t720 343.579
R614 VDDD.n1300 VDDD.t815 343.579
R615 VDDD.n641 VDDD.t118 343.577
R616 VDDD.n676 VDDD.t1387 343.577
R617 VDDD.n710 VDDD.t716 343.577
R618 VDDD.n745 VDDD.t771 343.577
R619 VDDD.n779 VDDD.t1032 343.577
R620 VDDD.n814 VDDD.t147 343.577
R621 VDDD.n848 VDDD.t1362 343.577
R622 VDDD.n883 VDDD.t79 343.577
R623 VDDD.n917 VDDD.t318 343.577
R624 VDDD.n952 VDDD.t600 343.577
R625 VDDD.n1612 VDDD.t963 343.577
R626 VDDD.n1579 VDDD.t1046 343.577
R627 VDDD.n1546 VDDD.t1250 343.577
R628 VDDD.n1513 VDDD.t1262 343.577
R629 VDDD.n1480 VDDD.t89 343.577
R630 VDDD.n1119 VDDD.t579 343.577
R631 VDDD.n1156 VDDD.t655 343.577
R632 VDDD.n1193 VDDD.t1244 343.577
R633 VDDD.n1230 VDDD.t413 343.577
R634 VDDD.n1267 VDDD.t347 343.577
R635 VDDD.n1848 VDDD.t470 342.377
R636 VDDD.n1854 VDDD.t1431 338.892
R637 VDDD.t542 VDDD 335.69
R638 VDDD.n1109 VDDD.n1108 325.627
R639 VDDD.n1109 VDDD.n1107 325.627
R640 VDDD.n272 VDDD.n270 320.976
R641 VDDD.n269 VDDD.n268 320.976
R642 VDDD.n1846 VDDD.n1845 320.976
R643 VDDD.n1868 VDDD.n1850 320.976
R644 VDDD.n1862 VDDD.n1861 320.976
R645 VDDD.n1860 VDDD.n1853 320.976
R646 VDDD.n5 VDDD.n4 320.976
R647 VDDD.n1004 VDDD.n3 320.976
R648 VDDD.n1474 VDDD.n1446 320.976
R649 VDDD.n1450 VDDD.n1449 320.976
R650 VDDD.t601 VDDD.t488 319.627
R651 VDDD.t897 VDDD.t311 319.627
R652 VDDD.t701 VDDD.t1268 319.627
R653 VDDD.t32 VDDD.t819 319.627
R654 VDDD.t1013 VDDD.t1187 319.627
R655 VDDD.t909 VDDD.t1217 319.627
R656 VDDD.t243 VDDD.t914 319.627
R657 VDDD.t397 VDDD.t486 319.627
R658 VDDD.t928 VDDD.t492 319.627
R659 VDDD.t1245 VDDD.t784 319.627
R660 VDDD.t1416 VDDD.t405 319.627
R661 VDDD.t1197 VDDD.t54 319.627
R662 VDDD.t895 VDDD.t156 319.627
R663 VDDD.t205 VDDD.t276 319.627
R664 VDDD.t1199 VDDD.t44 319.627
R665 VDDD.t303 VDDD.t1398 319.627
R666 VDDD.t179 VDDD.t525 319.627
R667 VDDD.t292 VDDD.t105 319.627
R668 VDDD.t1062 VDDD.t574 319.627
R669 VDDD.t782 VDDD.t987 319.627
R670 VDDD.t1318 VDDD.t556 319.627
R671 VDDD.t294 VDDD.t1129 319.627
R672 VDDD.t966 VDDD.t970 319.627
R673 VDDD.t1043 VDDD.t1071 319.627
R674 VDDD.t1253 VDDD.t617 319.627
R675 VDDD.t1264 VDDD.t115 319.627
R676 VDDD.t1142 VDDD.t169 319.627
R677 VDDD.t515 VDDD.t1231 319.627
R678 VDDD.t849 VDDD.t1086 319.627
R679 VDDD.t632 VDDD.t676 319.627
R680 VDDD.t1272 VDDD.t1367 319.627
R681 VDDD.t968 VDDD.t1308 319.627
R682 VDDD.t1009 VDDD.t463 319.627
R683 VDDD.t336 VDDD.t502 319.627
R684 VDDD.t711 VDDD.t261 319.627
R685 VDDD.t725 VDDD.t851 319.627
R686 VDDD.t1033 VDDD.t1274 319.627
R687 VDDD.t370 VDDD.t490 319.627
R688 VDDD.t1359 VDDD.t1314 319.627
R689 VDDD.t76 VDDD.t513 319.627
R690 VDDD.t315 VDDD.t847 319.627
R691 VDDD.t23 VDDD.t498 319.627
R692 VDDD VDDD.t1306 313.707
R693 VDDD.t323 VDDD 313.707
R694 VDDD.t1324 VDDD.t372 312.192
R695 VDDD.t1320 VDDD.t1408 312.192
R696 VDDD.t1058 VDDD.t893 312.192
R697 VDDD.t199 VDDD.t296 312.192
R698 VDDD.t203 VDDD.t1344 312.192
R699 VDDD.n280 VDDD.n279 310.502
R700 VDDD.n265 VDDD.n264 310.502
R701 VDDD.n287 VDDD.n286 310.502
R702 VDDD.n988 VDDD.n987 310.5
R703 VDDD.n990 VDDD.n989 310.5
R704 VDDD.n997 VDDD.n996 310.5
R705 VDDD.n1467 VDDD.n1451 310.5
R706 VDDD.n1455 VDDD.n1454 310.5
R707 VDDD.n1461 VDDD.n1456 310.5
R708 VDDD.t1235 VDDD.t18 292.991
R709 VDDD.t65 VDDD.t109 292.991
R710 VDDD.t1081 VDDD.t1104 292.991
R711 VDDD.t935 VDDD.t1297 292.991
R712 VDDD.t1227 VDDD.t916 292.991
R713 VDDD.t233 VDDD.t151 292.991
R714 VDDD.t259 VDDD.t1079 292.991
R715 VDDD.t790 VDDD.t1080 292.991
R716 VDDD.t1066 VDDD.t1405 292.991
R717 VDDD.t96 VDDD.t1402 292.991
R718 VDDD.t434 VDDD.t1395 292.991
R719 VDDD.t739 VDDD.t1394 292.991
R720 VDDD.t61 VDDD.t436 292.991
R721 VDDD.t1226 VDDD.t1277 292.991
R722 VDDD.t1073 VDDD.t1157 292.991
R723 VDDD.t767 VDDD.t1158 292.991
R724 VDDD.t458 VDDD.t805 292.991
R725 VDDD.t148 VDDD.t804 292.991
R726 VDDD.t381 VDDD.t794 292.991
R727 VDDD.t145 VDDD.t793 292.991
R728 VDDD.t251 VDDD.t1169 292.991
R729 VDDD.t248 VDDD.t383 292.991
R730 VDDD.t14 VDDD.t15 292.991
R731 VDDD.t357 VDDD.t56 292.991
R732 VDDD.t477 VDDD.t859 292.991
R733 VDDD.t512 VDDD.t675 292.991
R734 VDDD.t1375 VDDD.t1166 292.991
R735 VDDD.t447 VDDD.t437 292.991
R736 VDDD.t396 VDDD.t442 292.991
R737 VDDD.t772 VDDD.t747 292.991
R738 VDDD.t1172 VDDD.t548 292.991
R739 VDDD.t1171 VDDD.t431 292.991
R740 VDDD.t1207 VDDD.t420 292.991
R741 VDDD.t1330 VDDD.t1363 292.991
R742 VDDD.t764 VDDD.t682 292.991
R743 VDDD.t352 VDDD.t532 292.991
R744 VDDD.t1348 VDDD.t703 292.991
R745 VDDD.t855 VDDD.t444 292.991
R746 VDDD.t124 VDDD.t350 292.991
R747 VDDD.t657 VDDD.t1223 292.991
R748 VDDD.t1456 VDDD.t330 292.991
R749 VDDD.t818 VDDD.t17 292.991
R750 VDDD.t589 VDDD.t688 292.991
R751 VDDD.t1133 VDDD.t252 292.991
R752 VDDD.t841 VDDD.t1328 292.991
R753 VDDD.t94 VDDD.t1329 292.991
R754 VDDD.t1096 VDDD.t1427 292.991
R755 VDDD.t1233 VDDD.t697 292.991
R756 VDDD.t985 VDDD.t1263 292.991
R757 VDDD.t360 VDDD.t247 292.991
R758 VDDD.t842 VDDD.t362 292.991
R759 VDDD.t467 VDDD.t363 292.991
R760 VDDD.t1164 VDDD.t598 292.991
R761 VDDD.t1326 VDDD.t1156 292.991
R762 VDDD.t623 VDDD.t454 292.991
R763 VDDD.t504 VDDD.t143 292.991
R764 VDDD.t366 VDDD.t517 292.991
R765 VDDD.t369 VDDD.t60 292.991
R766 VDDD.t571 VDDD.t213 292.991
R767 VDDD.t123 VDDD.t943 292.991
R768 VDDD.t29 VDDD.t881 292.991
R769 VDDD.t791 VDDD.t1339 292.991
R770 VDDD.t25 VDDD.t456 292.991
R771 VDDD.t26 VDDD.t1099 292.991
R772 VDDD.t1107 VDDD.t950 292.991
R773 VDDD.t374 VDDD.t947 292.991
R774 VDDD.t1195 VDDD.t1176 292.991
R775 VDDD.t933 VDDD.t1173 292.991
R776 VDDD.t332 VDDD.t497 292.991
R777 VDDD.t1189 VDDD.t273 292.991
R778 VDDD.t193 VDDD.t1150 292.991
R779 VDDD.t524 VDDD.t1151 292.991
R780 VDDD.t594 VDDD.t751 292.991
R781 VDDD.t564 VDDD.t750 292.991
R782 VDDD.t587 VDDD.t310 292.991
R783 VDDD.t742 VDDD.t307 292.991
R784 VDDD.t27 VDDD.t590 292.991
R785 VDDD.t380 VDDD.t57 292.991
R786 VDDD.t723 VDDD.t494 292.991
R787 VDDD.t981 VDDD.t775 292.991
R788 VDDD.t1282 VDDD.t638 292.991
R789 VDDD.t166 VDDD.t639 292.991
R790 VDDD.t845 VDDD.t921 292.991
R791 VDDD.t998 VDDD.t1165 292.991
R792 VDDD VDDD.t469 290.031
R793 VDDD.t540 VDDD.t1219 287.072
R794 VDDD.t611 VDDD.t615 287.072
R795 VDDD.t1298 VDDD.t500 287.072
R796 VDDD.t835 VDDD.t823 287.072
R797 VDDD.t1337 VDDD.t465 287.072
R798 VDDD.t889 VDDD.t1215 287.072
R799 VDDD.t529 VDDD.t1316 287.072
R800 VDDD.t797 VDDD.t899 287.072
R801 VDDD.t1378 VDDD.t903 287.072
R802 VDDD.t1237 VDDD.t630 287.072
R803 VDDD.t1322 VDDD.t1280 287.072
R804 VDDD.t12 VDDD.t560 287.072
R805 VDDD.t1412 VDDD.t919 287.072
R806 VDDD.t10 VDDD.t418 287.072
R807 VDDD.t1414 VDDD.t558 287.072
R808 VDDD.t868 VDDD.t673 287.072
R809 VDDD.t776 VDDD.t135 287.072
R810 VDDD.t624 VDDD.t646 287.072
R811 VDDD.t1346 VDDD.t870 287.072
R812 VDDD.t780 VDDD.t113 287.072
R813 VDDD.t1064 VDDD.t709 287.072
R814 VDDD.t181 VDDD.t508 287.072
R815 VDDD.t328 VDDD.t265 287.072
R816 VDDD.t650 VDDD.t482 287.072
R817 VDDD.t1097 VDDD.t313 287.072
R818 VDDD.t640 VDDD.t1270 287.072
R819 VDDD.t879 VDDD.t821 287.072
R820 VDDD.t907 VDDD.t448 287.072
R821 VDDD.t1302 VDDD.t1180 287.072
R822 VDDD.t544 VDDD.t257 287.072
R823 VDDD.t1300 VDDD.t452 287.072
R824 VDDD.t636 VDDD.t1027 287.072
R825 VDDD.t1355 VDDD.t905 287.072
R826 VDDD.t605 VDDD.t1304 287.072
R827 VDDD.t808 VDDD.t613 287.072
R828 VDDD.t999 VDDD.t1312 287.072
R829 VDDD.t141 VDDD.t171 287.072
R830 VDDD.t298 VDDD.t634 287.072
R831 VDDD.t745 VDDD.t546 287.072
R832 VDDD.t686 VDDD.t263 287.072
R833 VDDD.t154 VDDD.t901 287.072
R834 VDDD.t355 VDDD.t1213 287.072
R835 VDDD.t1450 VDDD.t65 272.274
R836 VDDD.t97 VDDD.t935 272.274
R837 VDDD.t662 VDDD.t233 272.274
R838 VDDD.t237 VDDD.t790 272.274
R839 VDDD.t416 VDDD.t96 272.274
R840 VDDD.t99 VDDD.t739 272.274
R841 VDDD.t235 VDDD.t1226 272.274
R842 VDDD.t36 VDDD.t767 272.274
R843 VDDD.t660 VDDD.t148 272.274
R844 VDDD.t1452 VDDD.t145 272.274
R845 VDDD.t383 VDDD.t127 272.274
R846 VDDD.t56 VDDD.t1342 272.274
R847 VDDD.t675 VDDD.t865 272.274
R848 VDDD.t437 VDDD.t1255 272.274
R849 VDDD.t747 VDDD.t621 272.274
R850 VDDD.t431 VDDD.t505 272.274
R851 VDDD.t1363 VDDD.t375 272.274
R852 VDDD.t532 VDDD.t816 272.274
R853 VDDD.t444 VDDD.t733 272.274
R854 VDDD.t1223 VDDD.t995 272.274
R855 VDDD.t17 VDDD.t729 272.274
R856 VDDD.t252 VDDD.t1432 272.274
R857 VDDD.t533 VDDD.t841 272.274
R858 VDDD.t0 VDDD.t1096 272.274
R859 VDDD.t1289 VDDD.t985 272.274
R860 VDDD.t669 VDDD.t842 272.274
R861 VDDD.t82 VDDD.t1164 272.274
R862 VDDD.t143 VDDD.t133 272.274
R863 VDDD.t60 VDDD.t239 272.274
R864 VDDD.t943 VDDD.t642 272.274
R865 VDDD.t1339 VDDD.t1380 272.274
R866 VDDD.t1099 VDDD.t1203 272.274
R867 VDDD.t1037 VDDD.t374 272.274
R868 VDDD.t705 VDDD.t933 272.274
R869 VDDD.t1120 VDDD.t1189 272.274
R870 VDDD.t707 VDDD.t524 272.274
R871 VDDD.t1122 VDDD.t564 272.274
R872 VDDD.t1118 VDDD.t742 272.274
R873 VDDD.t1039 VDDD.t380 272.274
R874 VDDD.t1185 VDDD.t981 272.274
R875 VDDD.t1041 VDDD.t166 272.274
R876 VDDD.t1183 VDDD.t998 272.274
R877 VDDD.n1855 VDDD.t1307 260.134
R878 VDDD.n2273 VDDD.t324 255.905
R879 VDDD.n1881 VDDD.t620 255.905
R880 VDDD.t18 VDDD.t858 254.518
R881 VDDD.t1104 VDDD.t934 254.518
R882 VDDD.t916 VDDD.t1182 254.518
R883 VDDD.t1079 VDDD.t610 254.518
R884 VDDD.t1405 VDDD.t740 254.518
R885 VDDD.t1395 VDDD.t738 254.518
R886 VDDD.t436 VDDD.t1225 254.518
R887 VDDD.t1157 VDDD.t593 254.518
R888 VDDD.t805 VDDD.t1128 254.518
R889 VDDD.t794 VDDD.t144 254.518
R890 VDDD.t110 VDDD.t251 254.518
R891 VDDD.t9 VDDD.t14 254.518
R892 VDDD.t972 VDDD.t477 254.518
R893 VDDD.t409 VDDD.t1375 254.518
R894 VDDD.t876 VDDD.t396 254.518
R895 VDDD.t430 VDDD.t1172 254.518
R896 VDDD.t1364 VDDD.t1207 254.518
R897 VDDD.t531 VDDD.t764 254.518
R898 VDDD.t607 VDDD.t1348 254.518
R899 VDDD.t1224 VDDD.t124 254.518
R900 VDDD.t8 VDDD.t1456 254.518
R901 VDDD.t582 VDDD.t589 254.518
R902 VDDD.t1329 VDDD.t840 254.518
R903 VDDD.t697 VDDD.t1095 254.518
R904 VDDD.t247 VDDD.t986 254.518
R905 VDDD.t363 VDDD.t837 254.518
R906 VDDD.t1156 VDDD.t1163 254.518
R907 VDDD.t1208 VDDD.t623 254.518
R908 VDDD.t664 VDDD.t366 254.518
R909 VDDD.t944 VDDD.t571 254.518
R910 VDDD.t690 VDDD.t29 254.518
R911 VDDD.t930 VDDD.t25 254.518
R912 VDDD.t950 VDDD.t234 254.518
R913 VDDD.t1176 VDDD.t519 254.518
R914 VDDD.t497 VDDD.t1190 254.518
R915 VDDD.t1150 VDDD.t735 254.518
R916 VDDD.t751 VDDD.t801 254.518
R917 VDDD.t310 VDDD.t741 254.518
R918 VDDD.t590 VDDD.t379 254.518
R919 VDDD.t494 VDDD.t982 254.518
R920 VDDD.t638 VDDD.t1168 254.518
R921 VDDD.t921 VDDD.t997 254.518
R922 VDDD.n1883 VDDD.t769 252.95
R923 VDDD.n1835 VDDD.n1834 252.213
R924 VDDD.n1976 VDDD.n1975 252.213
R925 VDDD.n2268 VDDD.n2267 252.213
R926 VDDD.n1649 VDDD.n1648 252.213
R927 VDDD.n1662 VDDD.n1661 252.213
R928 VDDD.n1098 VDDD.n1096 252.213
R929 VDDD.n327 VDDD.t161 250.464
R930 VDDD.n235 VDDD.t749 250.464
R931 VDDD.n396 VDDD.t1350 250.464
R932 VDDD.n210 VDDD.t93 250.464
R933 VDDD.n465 VDDD.t220 250.464
R934 VDDD.n185 VDDD.t1424 250.464
R935 VDDD.n534 VDDD.t1385 250.464
R936 VDDD.n160 VDDD.t755 250.464
R937 VDDD.n603 VDDD.t1147 250.464
R938 VDDD.n635 VDDD.t1370 250.464
R939 VDDD.n2190 VDDD.t1352 250.464
R940 VDDD.n2204 VDDD.t553 250.464
R941 VDDD.n2218 VDDD.t990 250.464
R942 VDDD.n2232 VDDD.t937 250.464
R943 VDDD.n2246 VDDD.t108 250.464
R944 VDDD.n2260 VDDD.t528 250.464
R945 VDDD.n1898 VDDD.t198 250.464
R946 VDDD.n1912 VDDD.t49 250.464
R947 VDDD.n1926 VDDD.t279 250.464
R948 VDDD.n1940 VDDD.t159 250.464
R949 VDDD.n1954 VDDD.t728 250.464
R950 VDDD.n1968 VDDD.t408 250.464
R951 VDDD.n1319 VDDD.t1311 250.464
R952 VDDD.n1333 VDDD.t378 250.464
R953 VDDD.n1347 VDDD.t679 250.464
R954 VDDD.n1361 VDDD.t1085 250.464
R955 VDDD.n1375 VDDD.t322 250.464
R956 VDDD.n1302 VDDD.t811 250.464
R957 VDDD.n1151 VDDD.t523 250.464
R958 VDDD.n1188 VDDD.t1139 250.464
R959 VDDD.n1225 VDDD.t138 250.464
R960 VDDD.n1262 VDDD.t281 250.464
R961 VDDD.n637 VDDD.t1008 250.463
R962 VDDD.n123 VDDD.t335 250.463
R963 VDDD.n706 VDDD.t714 250.463
R964 VDDD.n98 VDDD.t81 250.463
R965 VDDD.n775 VDDD.t1036 250.463
R966 VDDD.n73 VDDD.t184 250.463
R967 VDDD.n844 VDDD.t1358 250.463
R968 VDDD.n48 VDDD.t864 250.463
R969 VDDD.n913 VDDD.t320 250.463
R970 VDDD.n23 VDDD.t22 250.463
R971 VDDD.n1389 VDDD.t965 250.463
R972 VDDD.n1403 VDDD.t1076 250.463
R973 VDDD.n1417 VDDD.t1252 250.463
R974 VDDD.n1431 VDDD.t1332 250.463
R975 VDDD.n1445 VDDD.t87 250.463
R976 VDDD.n1115 VDDD.t577 250.463
R977 VDDD.n1152 VDDD.t653 250.463
R978 VDDD.n1189 VDDD.t1242 250.463
R979 VDDD.n1226 VDDD.t803 250.463
R980 VDDD.n1263 VDDD.t349 250.463
R981 VDDD.n1880 VDDD.t192 248.843
R982 VDDD.t1371 VDDD.t1369 248.599
R983 VDDD.t488 VDDD.t1110 248.599
R984 VDDD.t858 VDDD.t601 248.599
R985 VDDD.t284 VDDD.t19 248.599
R986 VDDD.t1144 VDDD.t1146 248.599
R987 VDDD.t311 VDDD.t931 248.599
R988 VDDD.t934 VDDD.t897 248.599
R989 VDDD.t644 VDDD.t1102 248.599
R990 VDDD.t699 VDDD.t754 248.599
R991 VDDD.t1268 VDDD.t255 248.599
R992 VDDD.t1182 VDDD.t701 248.599
R993 VDDD.t983 VDDD.t152 248.599
R994 VDDD.t34 VDDD.t1384 248.599
R995 VDDD.t819 VDDD.t562 248.599
R996 VDDD.t610 VDDD.t32 248.599
R997 VDDD.t131 VDDD.t209 248.599
R998 VDDD.t1011 VDDD.t1423 248.599
R999 VDDD.t1187 VDDD.t1159 248.599
R1000 VDDD.t740 VDDD.t1013 248.599
R1001 VDDD.t537 VDDD.t1403 248.599
R1002 VDDD.t217 VDDD.t219 248.599
R1003 VDDD.t1217 VDDD.t550 248.599
R1004 VDDD.t738 VDDD.t909 248.599
R1005 VDDD.t2 VDDD.t760 248.599
R1006 VDDD.t90 VDDD.t92 248.599
R1007 VDDD.t914 VDDD.t991 248.599
R1008 VDDD.t1225 VDDD.t243 248.599
R1009 VDDD.t1291 VDDD.t58 248.599
R1010 VDDD.t1335 VDDD.t1349 248.599
R1011 VDDD.t486 VDDD.t1154 248.599
R1012 VDDD.t593 VDDD.t397 248.599
R1013 VDDD.t667 VDDD.t833 248.599
R1014 VDDD.t861 VDDD.t748 248.599
R1015 VDDD.t492 VDDD.t1457 248.599
R1016 VDDD.t1128 VDDD.t928 248.599
R1017 VDDD.t84 VDDD.t806 248.599
R1018 VDDD.t1247 VDDD.t160 248.599
R1019 VDDD.t784 VDDD.t288 248.599
R1020 VDDD.t144 VDDD.t1245 248.599
R1021 VDDD.t975 VDDD.t125 248.599
R1022 VDDD.t887 VDDD.t269 248.599
R1023 VDDD.t410 VDDD.t887 248.599
R1024 VDDD.t271 VDDD.t410 248.599
R1025 VDDD.t185 VDDD.t271 248.599
R1026 VDDD.t211 VDDD.t185 248.599
R1027 VDDD.t885 VDDD.t211 248.599
R1028 VDDD.t187 VDDD.t885 248.599
R1029 VDDD.t665 VDDD.t187 248.599
R1030 VDDD.t926 VDDD.t665 248.599
R1031 VDDD.t924 VDDD.t926 248.599
R1032 VDDD.t471 VDDD.t1430 248.599
R1033 VDDD.t173 VDDD.t471 248.599
R1034 VDDD.t1428 VDDD.t173 248.599
R1035 VDDD.t572 VDDD.t1428 248.599
R1036 VDDD.t473 VDDD.t572 248.599
R1037 VDDD.t225 VDDD.t473 248.599
R1038 VDDD.t469 VDDD.t225 248.599
R1039 VDDD.t189 VDDD.t129 248.599
R1040 VDDD.t1003 VDDD.t189 248.599
R1041 VDDD.t191 VDDD.t1003 248.599
R1042 VDDD.t768 VDDD.t619 248.599
R1043 VDDD.t407 VDDD.t403 248.599
R1044 VDDD.t684 VDDD.t1416 248.599
R1045 VDDD.t405 VDDD.t110 248.599
R1046 VDDD.t249 VDDD.t565 248.599
R1047 VDDD.t727 VDDD.t52 248.599
R1048 VDDD.t786 VDDD.t1197 248.599
R1049 VDDD.t54 VDDD.t9 248.599
R1050 VDDD.t358 VDDD.t1112 248.599
R1051 VDDD.t158 VDDD.t460 248.599
R1052 VDDD.t326 VDDD.t895 248.599
R1053 VDDD.t156 VDDD.t972 248.599
R1054 VDDD.t510 VDDD.t1017 248.599
R1055 VDDD.t278 VDDD.t1029 248.599
R1056 VDDD.t648 VDDD.t205 248.599
R1057 VDDD.t276 VDDD.t409 248.599
R1058 VDDD.t843 VDDD.t338 248.599
R1059 VDDD.t48 VDDD.t50 248.599
R1060 VDDD.t1257 VDDD.t1199 248.599
R1061 VDDD.t44 VDDD.t876 248.599
R1062 VDDD.t394 VDDD.t567 248.599
R1063 VDDD.t197 VDDD.t195 248.599
R1064 VDDD.t432 VDDD.t303 248.599
R1065 VDDD.t1398 VDDD.t430 248.599
R1066 VDDD.t1285 VDDD.t1049 248.599
R1067 VDDD.t527 VDDD.t231 248.599
R1068 VDDD.t438 VDDD.t179 248.599
R1069 VDDD.t525 VDDD.t1364 248.599
R1070 VDDD.t1205 VDDD.t340 248.599
R1071 VDDD.t107 VDDD.t103 248.599
R1072 VDDD.t101 VDDD.t292 248.599
R1073 VDDD.t105 VDDD.t531 248.599
R1074 VDDD.t353 VDDD.t1116 248.599
R1075 VDDD.t936 VDDD.t583 248.599
R1076 VDDD.t960 VDDD.t1062 248.599
R1077 VDDD.t574 VDDD.t607 248.599
R1078 VDDD.t856 VDDD.t1019 248.599
R1079 VDDD.t989 VDDD.t1209 248.599
R1080 VDDD.t450 VDDD.t782 248.599
R1081 VDDD.t987 VDDD.t1224 248.599
R1082 VDDD.t658 VDDD.t344 248.599
R1083 VDDD.t552 VDDD.t554 248.599
R1084 VDDD.t608 VDDD.t1318 248.599
R1085 VDDD.t556 VDDD.t8 248.599
R1086 VDDD.t973 VDDD.t342 248.599
R1087 VDDD.t1351 VDDD.t1353 248.599
R1088 VDDD.t1382 VDDD.t294 248.599
R1089 VDDD.t1129 VDDD.t582 248.599
R1090 VDDD.t1161 VDDD.t1025 248.599
R1091 VDDD.t1051 VDDD.t440 248.599
R1092 VDDD.t840 VDDD.t966 248.599
R1093 VDDD.t970 VDDD.t1396 248.599
R1094 VDDD.t962 VDDD.t964 248.599
R1095 VDDD.t829 VDDD.t1425 248.599
R1096 VDDD.t1095 VDDD.t1043 248.599
R1097 VDDD.t1071 VDDD.t799 248.599
R1098 VDDD.t1045 VDDD.t1075 248.599
R1099 VDDD.t1114 VDDD.t245 248.599
R1100 VDDD.t986 VDDD.t1253 248.599
R1101 VDDD.t617 VDDD.t1295 248.599
R1102 VDDD.t1249 VDDD.t1251 248.599
R1103 VDDD.t825 VDDD.t1005 248.599
R1104 VDDD.t837 VDDD.t1264 248.599
R1105 VDDD.t115 VDDD.t221 248.599
R1106 VDDD.t1261 VDDD.t1331 248.599
R1107 VDDD.t693 VDDD.t596 248.599
R1108 VDDD.t1163 VDDD.t1142 248.599
R1109 VDDD.t169 VDDD.t475 248.599
R1110 VDDD.t88 VDDD.t86 248.599
R1111 VDDD.t979 VDDD.t1420 248.599
R1112 VDDD.t1420 VDDD.t422 248.599
R1113 VDDD.t422 VDDD.t1090 248.599
R1114 VDDD.t1090 VDDD.t1440 248.599
R1115 VDDD.t1440 VDDD.t1092 248.599
R1116 VDDD.t1092 VDDD.t1446 248.599
R1117 VDDD.t1446 VDDD.t1442 248.599
R1118 VDDD.t1442 VDDD.t671 248.599
R1119 VDDD.t671 VDDD.t1448 248.599
R1120 VDDD.t1448 VDDD.t1444 248.599
R1121 VDDD.t321 VDDD.t1229 248.599
R1122 VDDD.t1239 VDDD.t515 248.599
R1123 VDDD.t1231 VDDD.t1208 248.599
R1124 VDDD.t1259 VDDD.t1047 248.599
R1125 VDDD.t1084 VDDD.t1088 248.599
R1126 VDDD.t1068 VDDD.t849 248.599
R1127 VDDD.t1086 VDDD.t664 248.599
R1128 VDDD.t367 VDDD.t1023 248.599
R1129 VDDD.t678 VDDD.t680 248.599
R1130 VDDD.t1105 VDDD.t632 248.599
R1131 VDDD.t676 VDDD.t944 248.599
R1132 VDDD.t121 VDDD.t827 248.599
R1133 VDDD.t377 VDDD.t1365 248.599
R1134 VDDD.t1134 VDDD.t1272 248.599
R1135 VDDD.t1367 VDDD.t690 248.599
R1136 VDDD.t30 VDDD.t1021 248.599
R1137 VDDD.t1310 VDDD.t229 248.599
R1138 VDDD.t1211 VDDD.t968 248.599
R1139 VDDD.t1308 VDDD.t930 248.599
R1140 VDDD.t364 VDDD.t1053 248.599
R1141 VDDD.t117 VDDD.t1007 248.599
R1142 VDDD.t463 VDDD.t691 248.599
R1143 VDDD.t234 VDDD.t1009 248.599
R1144 VDDD.t282 VDDD.t948 248.599
R1145 VDDD.t1386 VDDD.t334 248.599
R1146 VDDD.t502 VDDD.t731 248.599
R1147 VDDD.t519 VDDD.t336 248.599
R1148 VDDD.t917 VDDD.t1174 248.599
R1149 VDDD.t715 VDDD.t713 248.599
R1150 VDDD.t261 VDDD.t580 248.599
R1151 VDDD.t1190 VDDD.t711 248.599
R1152 VDDD.t241 VDDD.t274 248.599
R1153 VDDD.t770 VDDD.t80 248.599
R1154 VDDD.t851 VDDD.t603 248.599
R1155 VDDD.t735 VDDD.t725 248.599
R1156 VDDD.t717 VDDD.t1001 248.599
R1157 VDDD.t1031 VDDD.t1035 248.599
R1158 VDDD.t1274 VDDD.t63 248.599
R1159 VDDD.t801 VDDD.t1033 248.599
R1160 VDDD.t535 VDDD.t752 248.599
R1161 VDDD.t146 VDDD.t183 248.599
R1162 VDDD.t490 VDDD.t301 248.599
R1163 VDDD.t741 VDDD.t370 248.599
R1164 VDDD.t4 VDDD.t308 248.599
R1165 VDDD.t1361 VDDD.t1357 248.599
R1166 VDDD.t1314 VDDD.t736 248.599
R1167 VDDD.t379 VDDD.t1359 248.599
R1168 VDDD.t1287 VDDD.t591 248.599
R1169 VDDD.t78 VDDD.t863 248.599
R1170 VDDD.t513 VDDD.t695 248.599
R1171 VDDD.t982 VDDD.t76 248.599
R1172 VDDD.t853 VDDD.t773 248.599
R1173 VDDD.t317 VDDD.t319 248.599
R1174 VDDD.t847 VDDD.t1136 248.599
R1175 VDDD.t1168 VDDD.t315 248.599
R1176 VDDD.t1131 VDDD.t6 248.599
R1177 VDDD.t599 VDDD.t21 248.599
R1178 VDDD.t498 VDDD.t74 248.599
R1179 VDDD.t997 VDDD.t23 248.599
R1180 VDDD.t977 VDDD.t922 248.599
R1181 VDDD.t399 VDDD.t384 248.599
R1182 VDDD.t401 VDDD.t399 248.599
R1183 VDDD.t386 VDDD.t401 248.599
R1184 VDDD.t390 VDDD.t386 248.599
R1185 VDDD.t1454 VDDD.t390 248.599
R1186 VDDD.t267 VDDD.t1454 248.599
R1187 VDDD.t388 VDDD.t267 248.599
R1188 VDDD.t480 VDDD.t388 248.599
R1189 VDDD.t286 VDDD.t480 248.599
R1190 VDDD.t478 VDDD.t286 248.599
R1191 VDDD.n289 VDDD.t270 243.512
R1192 VDDD.n9 VDDD.t385 243.512
R1193 VDDD.n1457 VDDD.t1445 243.512
R1194 VDDD.n1096 VDDD 236.78
R1195 VDDD VDDD.t191 221.964
R1196 VDDD VDDD.t768 198.287
R1197 VDDD VDDD.t284 192.369
R1198 VDDD VDDD.t644 192.369
R1199 VDDD VDDD.t983 192.369
R1200 VDDD VDDD.t131 192.369
R1201 VDDD VDDD.t537 192.369
R1202 VDDD VDDD.t2 192.369
R1203 VDDD VDDD.t1291 192.369
R1204 VDDD VDDD.t667 192.369
R1205 VDDD VDDD.t84 192.369
R1206 VDDD VDDD.t975 192.369
R1207 VDDD.t565 VDDD 192.369
R1208 VDDD.t1112 VDDD 192.369
R1209 VDDD.t1017 VDDD 192.369
R1210 VDDD.t338 VDDD 192.369
R1211 VDDD.t567 VDDD 192.369
R1212 VDDD.t1049 VDDD 192.369
R1213 VDDD.t340 VDDD 192.369
R1214 VDDD.t1116 VDDD 192.369
R1215 VDDD.t1019 VDDD 192.369
R1216 VDDD.t344 VDDD 192.369
R1217 VDDD.t342 VDDD 192.369
R1218 VDDD.t1025 VDDD 192.369
R1219 VDDD.t1047 VDDD 192.369
R1220 VDDD.t1023 VDDD 192.369
R1221 VDDD.t827 VDDD 192.369
R1222 VDDD.t1021 VDDD 192.369
R1223 VDDD.t1053 VDDD 192.369
R1224 VDDD VDDD.t282 192.369
R1225 VDDD VDDD.t917 192.369
R1226 VDDD VDDD.t241 192.369
R1227 VDDD VDDD.t717 192.369
R1228 VDDD VDDD.t535 192.369
R1229 VDDD VDDD.t4 192.369
R1230 VDDD VDDD.t1287 192.369
R1231 VDDD VDDD.t853 192.369
R1232 VDDD VDDD.t1131 192.369
R1233 VDDD VDDD.t977 192.369
R1234 VDDD VDDD.t924 189.409
R1235 VDDD VDDD.t478 189.409
R1236 VDDD.n1840 VDDD.n1839 185
R1237 VDDD.n1837 VDDD.n1833 185
R1238 VDDD.n1836 VDDD.n1831 185
R1239 VDDD.n1836 VDDD.n1835 185
R1240 VDDD.n1841 VDDD.n1832 185
R1241 VDDD.n1834 VDDD.n1832 185
R1242 VDDD.n1978 VDDD.n1977 185
R1243 VDDD.n1977 VDDD.n1976 185
R1244 VDDD.n1972 VDDD.n1971 185
R1245 VDDD.n1975 VDDD.n1972 185
R1246 VDDD.n1973 VDDD.n1969 185
R1247 VDDD.n1979 VDDD.n1970 185
R1248 VDDD.n2270 VDDD.n2269 185
R1249 VDDD.n2269 VDDD.n2268 185
R1250 VDDD.n2264 VDDD.n2263 185
R1251 VDDD.n2267 VDDD.n2264 185
R1252 VDDD.n2265 VDDD.n2261 185
R1253 VDDD.n2271 VDDD.n2262 185
R1254 VDDD.n1646 VDDD.n1642 185
R1255 VDDD.n1652 VDDD.n1643 185
R1256 VDDD.n1651 VDDD.n1650 185
R1257 VDDD.n1650 VDDD.n1649 185
R1258 VDDD.n1645 VDDD.n1644 185
R1259 VDDD.n1648 VDDD.n1645 185
R1260 VDDD.n1659 VDDD.n1655 185
R1261 VDDD.n1665 VDDD.n1656 185
R1262 VDDD.n1664 VDDD.n1663 185
R1263 VDDD.n1663 VDDD.n1662 185
R1264 VDDD.n1658 VDDD.n1657 185
R1265 VDDD.n1661 VDDD.n1658 185
R1266 VDDD.n1097 VDDD.n1093 185
R1267 VDDD.n1098 VDDD.n1097 185
R1268 VDDD.n1095 VDDD.n1092 185
R1269 VDDD.n1101 VDDD.n1100 185
R1270 VDDD.n1102 VDDD.n1094 185
R1271 VDDD.n1096 VDDD.n1094 185
R1272 VDDD.t912 VDDD.t542 181.273
R1273 VDDD.n1839 VDDD.n1838 161.239
R1274 VDDD.n1974 VDDD.n1973 161.239
R1275 VDDD.n2266 VDDD.n2265 161.239
R1276 VDDD.n1647 VDDD.n1646 161.239
R1277 VDDD.n1660 VDDD.n1659 161.239
R1278 VDDD.n1099 VDDD.n1095 161.239
R1279 VDDD.t951 VDDD.t462 144.346
R1280 VDDD.t38 VDDD.t569 144.346
R1281 VDDD.t40 VDDD.t119 144.346
R1282 VDDD.t485 VDDD.t1284 144.346
R1283 VDDD.t1400 VDDD.t759 144.346
R1284 VDDD.t956 VDDD.t1333 144.346
R1285 VDDD.t585 VDDD.t1056 144.346
R1286 VDDD.t867 VDDD.t1192 144.346
R1287 VDDD.t911 VDDD.t424 144.346
R1288 VDDD.t872 VDDD.t428 144.346
R1289 VDDD.t762 VDDD.t891 144.346
R1290 VDDD.t1374 VDDD.t874 144.346
R1291 VDDD.t539 VDDD.t938 144.346
R1292 VDDD.t46 VDDD.t1015 144.346
R1293 VDDD.t164 VDDD.t215 144.346
R1294 VDDD.t629 VDDD.t1083 144.346
R1295 VDDD.t698 VDDD.t72 144.346
R1296 VDDD.t993 VDDD.t877 144.346
R1297 VDDD.t1376 VDDD.t1126 144.346
R1298 VDDD.t1179 VDDD.t207 144.346
R1299 VDDD.t945 VDDD.t912 140.989
R1300 VDDD.t576 VDDD.t167 127.562
R1301 VDDD.t883 VDDD.t522 127.562
R1302 VDDD.t652 VDDD.t765 127.562
R1303 VDDD.t757 VDDD.t1138 127.562
R1304 VDDD.t1241 VDDD.t445 127.562
R1305 VDDD.t425 VDDD.t137 127.562
R1306 VDDD.t802 VDDD.t1148 127.562
R1307 VDDD.t939 VDDD.t280 127.562
R1308 VDDD.t348 VDDD.t1177 127.562
R1309 VDDD.t70 VDDD.t810 127.562
R1310 VDDD.n251 VDDD.t1246 119.608
R1311 VDDD.n351 VDDD.t929 119.608
R1312 VDDD.n226 VDDD.t398 119.608
R1313 VDDD.n420 VDDD.t244 119.608
R1314 VDDD.n201 VDDD.t910 119.608
R1315 VDDD.n489 VDDD.t1014 119.608
R1316 VDDD.n176 VDDD.t33 119.608
R1317 VDDD.n558 VDDD.t702 119.608
R1318 VDDD.n151 VDDD.t898 119.608
R1319 VDDD.n627 VDDD.t602 119.608
R1320 VDDD.n131 VDDD.t1010 119.608
R1321 VDDD.n121 VDDD.t337 119.608
R1322 VDDD.n106 VDDD.t712 119.608
R1323 VDDD.n96 VDDD.t726 119.608
R1324 VDDD.n81 VDDD.t1034 119.608
R1325 VDDD.n71 VDDD.t371 119.608
R1326 VDDD.n56 VDDD.t1360 119.608
R1327 VDDD.n46 VDDD.t77 119.608
R1328 VDDD.n31 VDDD.t316 119.608
R1329 VDDD.n21 VDDD.t24 119.608
R1330 VDDD.n2187 VDDD.t1130 119.608
R1331 VDDD.n2200 VDDD.t557 119.608
R1332 VDDD.n2214 VDDD.t988 119.608
R1333 VDDD.n2228 VDDD.t575 119.608
R1334 VDDD.n2242 VDDD.t106 119.608
R1335 VDDD.n2256 VDDD.t526 119.608
R1336 VDDD.n1895 VDDD.t1399 119.608
R1337 VDDD.n1908 VDDD.t45 119.608
R1338 VDDD.n1922 VDDD.t277 119.608
R1339 VDDD.n1936 VDDD.t157 119.608
R1340 VDDD.n1950 VDDD.t55 119.608
R1341 VDDD.n1964 VDDD.t406 119.608
R1342 VDDD.n1385 VDDD.t967 119.608
R1343 VDDD.n1399 VDDD.t1044 119.608
R1344 VDDD.n1413 VDDD.t1254 119.608
R1345 VDDD.n1427 VDDD.t1265 119.608
R1346 VDDD.n1441 VDDD.t1143 119.608
R1347 VDDD.n1316 VDDD.t1309 119.608
R1348 VDDD.n1329 VDDD.t1368 119.608
R1349 VDDD.n1343 VDDD.t677 119.608
R1350 VDDD.n1357 VDDD.t1087 119.608
R1351 VDDD.n1371 VDDD.t1232 119.608
R1352 VDDD.n1085 VDDD.t942 119.608
R1353 VDDD.n1076 VDDD.t150 119.608
R1354 VDDD.n1068 VDDD.t291 119.608
R1355 VDDD.n1059 VDDD.t306 119.608
R1356 VDDD.n1051 VDDD.t496 119.608
R1357 VDDD.n1042 VDDD.t839 119.608
R1358 VDDD.n1034 VDDD.t415 119.608
R1359 VDDD.n1025 VDDD.t722 119.608
R1360 VDDD.n1017 VDDD.t1101 119.608
R1361 VDDD.n1292 VDDD.t813 119.608
R1362 VDDD.n1107 VDDD.t913 116.341
R1363 VDDD.n1108 VDDD.t1070 116.341
R1364 VDDD VDDD.t945 112.457
R1365 VDDD.t1152 VDDD 109.1
R1366 VDDD.t1438 VDDD 109.1
R1367 VDDD.t1436 VDDD 109.1
R1368 VDDD.t66 VDDD 109.1
R1369 VDDD.t68 VDDD 109.1
R1370 VDDD.t300 VDDD.t941 93.9934
R1371 VDDD.t149 VDDD.t952 93.9934
R1372 VDDD.t1191 VDDD.t290 93.9934
R1373 VDDD.t305 VDDD.t1401 93.9934
R1374 VDDD.t875 VDDD.t495 93.9934
R1375 VDDD.t838 VDDD.t792 93.9934
R1376 VDDD.t1422 VDDD.t414 93.9934
R1377 VDDD.t721 VDDD.t1109 93.9934
R1378 VDDD.t208 VDDD.t1100 93.9934
R1379 VDDD.t812 VDDD.t1276 93.9934
R1380 VDDD.n307 VDDD.t1238 93.81
R1381 VDDD.n243 VDDD.t1379 93.81
R1382 VDDD.n376 VDDD.t798 93.81
R1383 VDDD.n218 VDDD.t530 93.81
R1384 VDDD.n445 VDDD.t890 93.81
R1385 VDDD.n193 VDDD.t1338 93.81
R1386 VDDD.n514 VDDD.t836 93.81
R1387 VDDD.n168 VDDD.t1299 93.81
R1388 VDDD.n583 VDDD.t612 93.81
R1389 VDDD.n143 VDDD.t541 93.81
R1390 VDDD.n656 VDDD.t1356 93.81
R1391 VDDD.n115 VDDD.t606 93.81
R1392 VDDD.n725 VDDD.t809 93.81
R1393 VDDD.n90 VDDD.t1000 93.81
R1394 VDDD.n794 VDDD.t142 93.81
R1395 VDDD.n65 VDDD.t299 93.81
R1396 VDDD.n863 VDDD.t746 93.81
R1397 VDDD.n40 VDDD.t687 93.81
R1398 VDDD.n932 VDDD.t155 93.81
R1399 VDDD.n15 VDDD.t356 93.81
R1400 VDDD.n2457 VDDD.t509 93.81
R1401 VDDD.n2197 VDDD.t710 93.81
R1402 VDDD.n2211 VDDD.t114 93.81
R1403 VDDD.n2225 VDDD.t871 93.81
R1404 VDDD.n2239 VDDD.t647 93.81
R1405 VDDD.n2253 VDDD.t136 93.81
R1406 VDDD.n2161 VDDD.t674 93.81
R1407 VDDD.n1905 VDDD.t559 93.81
R1408 VDDD.n1919 VDDD.t419 93.81
R1409 VDDD.n1933 VDDD.t920 93.81
R1410 VDDD.n1947 VDDD.t561 93.81
R1411 VDDD.n1961 VDDD.t1281 93.81
R1412 VDDD.n1382 VDDD.t329 93.81
R1413 VDDD.n1396 VDDD.t651 93.81
R1414 VDDD.n1410 VDDD.t1098 93.81
R1415 VDDD.n1424 VDDD.t641 93.81
R1416 VDDD.n1438 VDDD.t880 93.81
R1417 VDDD.n1815 VDDD.t1028 93.81
R1418 VDDD.n1326 VDDD.t453 93.81
R1419 VDDD.n1340 VDDD.t258 93.81
R1420 VDDD.n1354 VDDD.t1181 93.81
R1421 VDDD.n1368 VDDD.t449 93.81
R1422 VDDD.n1082 VDDD.t39 93.81
R1423 VDDD.n1079 VDDD.t120 93.81
R1424 VDDD.n1065 VDDD.t957 93.81
R1425 VDDD.n1062 VDDD.t1057 93.81
R1426 VDDD.n1048 VDDD.t873 93.81
R1427 VDDD.n1045 VDDD.t892 93.81
R1428 VDDD.n1031 VDDD.t47 93.81
R1429 VDDD.n1028 VDDD.t216 93.81
R1430 VDDD.n1277 VDDD.t994 93.81
R1431 VDDD.n1285 VDDD.t1127 93.81
R1432 VDDD VDDD.t1051 91.745
R1433 VDDD VDDD.t829 91.745
R1434 VDDD VDDD.t1114 91.745
R1435 VDDD VDDD.t825 91.745
R1436 VDDD VDDD.t693 91.745
R1437 VDDD VDDD.t979 88.7855
R1438 VDDD.t626 VDDD.t300 87.2797
R1439 VDDD.t952 VDDD.t1410 87.2797
R1440 VDDD.t1406 VDDD.t1191 87.2797
R1441 VDDD.t1401 VDDD.t177 87.2797
R1442 VDDD.t175 VDDD.t875 87.2797
R1443 VDDD.t792 VDDD.t1060 87.2797
R1444 VDDD.t778 VDDD.t1422 87.2797
R1445 VDDD.t1109 VDDD.t201 87.2797
R1446 VDDD.t1418 VDDD.t208 87.2797
R1447 VDDD.t1276 VDDD.t1201 87.2797
R1448 VDDD.n1838 VDDD.n1834 82.0552
R1449 VDDD.n1975 VDDD.n1974 82.0552
R1450 VDDD.n2267 VDDD.n2266 82.0552
R1451 VDDD.n1648 VDDD.n1647 82.0552
R1452 VDDD.n1661 VDDD.n1660 82.0552
R1453 VDDD.n1099 VDDD.n1098 82.0552
R1454 VDDD.t253 VDDD.t1221 73.8521
R1455 VDDD.t958 VDDD.t162 73.8521
R1456 VDDD.t392 VDDD.t831 73.8521
R1457 VDDD.t1278 VDDD.t227 73.8521
R1458 VDDD.t1077 VDDD.t111 73.8521
R1459 VDDD.t795 VDDD.t743 73.8521
R1460 VDDD.t1293 VDDD.t1388 73.8521
R1461 VDDD.t42 VDDD.t1193 73.8521
R1462 VDDD.t953 VDDD.t1266 73.8521
R1463 VDDD.t1124 VDDD.t788 73.8521
R1464 VDDD.t941 VDDD.t484 72.1736
R1465 VDDD.t325 VDDD.t149 72.1736
R1466 VDDD.t290 VDDD.t955 72.1736
R1467 VDDD.t756 VDDD.t305 72.1736
R1468 VDDD.t495 VDDD.t1373 72.1736
R1469 VDDD.t427 VDDD.t838 72.1736
R1470 VDDD.t414 VDDD.t628 72.1736
R1471 VDDD.t507 VDDD.t721 72.1736
R1472 VDDD.t1100 VDDD.t1094 72.1736
R1473 VDDD.t73 VDDD.t812 72.1736
R1474 VDDD.t484 VDDD.t951 68.8168
R1475 VDDD.t1284 VDDD.t325 68.8168
R1476 VDDD.t955 VDDD.t1400 68.8168
R1477 VDDD.t1192 VDDD.t756 68.8168
R1478 VDDD.t1373 VDDD.t911 68.8168
R1479 VDDD.t874 VDDD.t427 68.8168
R1480 VDDD.t628 VDDD.t539 68.8168
R1481 VDDD.t1083 VDDD.t507 68.8168
R1482 VDDD.t1094 VDDD.t698 68.8168
R1483 VDDD.t207 VDDD.t73 68.8168
R1484 VDDD.n1838 VDDD.n1837 68.2267
R1485 VDDD.n1974 VDDD.n1970 68.2267
R1486 VDDD.n2266 VDDD.n2262 68.2267
R1487 VDDD.n1647 VDDD.n1643 68.2267
R1488 VDDD.n1660 VDDD.n1656 68.2267
R1489 VDDD.n1100 VDDD.n1099 68.2267
R1490 VDDD.t1221 VDDD.t626 67.1383
R1491 VDDD.t1410 VDDD.t958 67.1383
R1492 VDDD.t831 VDDD.t1406 67.1383
R1493 VDDD.t177 VDDD.t1278 67.1383
R1494 VDDD.t111 VDDD.t175 67.1383
R1495 VDDD.t1060 VDDD.t795 67.1383
R1496 VDDD.t1388 VDDD.t778 67.1383
R1497 VDDD.t201 VDDD.t42 67.1383
R1498 VDDD.t1266 VDDD.t1418 67.1383
R1499 VDDD.t1201 VDDD.t1124 67.1383
R1500 VDDD.n307 VDDD.t631 63.3219
R1501 VDDD.n251 VDDD.t785 63.3219
R1502 VDDD.n243 VDDD.t904 63.3219
R1503 VDDD.n351 VDDD.t493 63.3219
R1504 VDDD.n376 VDDD.t900 63.3219
R1505 VDDD.n226 VDDD.t487 63.3219
R1506 VDDD.n218 VDDD.t1317 63.3219
R1507 VDDD.n420 VDDD.t915 63.3219
R1508 VDDD.n445 VDDD.t1216 63.3219
R1509 VDDD.n201 VDDD.t1218 63.3219
R1510 VDDD.n193 VDDD.t466 63.3219
R1511 VDDD.n489 VDDD.t1188 63.3219
R1512 VDDD.n514 VDDD.t824 63.3219
R1513 VDDD.n176 VDDD.t820 63.3219
R1514 VDDD.n168 VDDD.t501 63.3219
R1515 VDDD.n558 VDDD.t1269 63.3219
R1516 VDDD.n583 VDDD.t616 63.3219
R1517 VDDD.n151 VDDD.t312 63.3219
R1518 VDDD.n143 VDDD.t1220 63.3219
R1519 VDDD.n627 VDDD.t489 63.3219
R1520 VDDD.n131 VDDD.t464 63.3219
R1521 VDDD.n656 VDDD.t906 63.3219
R1522 VDDD.n121 VDDD.t503 63.3219
R1523 VDDD.n115 VDDD.t1305 63.3219
R1524 VDDD.n106 VDDD.t262 63.3219
R1525 VDDD.n725 VDDD.t614 63.3219
R1526 VDDD.n96 VDDD.t852 63.3219
R1527 VDDD.n90 VDDD.t1313 63.3219
R1528 VDDD.n81 VDDD.t1275 63.3219
R1529 VDDD.n794 VDDD.t172 63.3219
R1530 VDDD.n71 VDDD.t491 63.3219
R1531 VDDD.n65 VDDD.t635 63.3219
R1532 VDDD.n56 VDDD.t1315 63.3219
R1533 VDDD.n863 VDDD.t547 63.3219
R1534 VDDD.n46 VDDD.t514 63.3219
R1535 VDDD.n40 VDDD.t264 63.3219
R1536 VDDD.n31 VDDD.t848 63.3219
R1537 VDDD.n932 VDDD.t902 63.3219
R1538 VDDD.n21 VDDD.t499 63.3219
R1539 VDDD.n15 VDDD.t1214 63.3219
R1540 VDDD.n2457 VDDD.t182 63.3219
R1541 VDDD.n2187 VDDD.t295 63.3219
R1542 VDDD.n2197 VDDD.t1065 63.3219
R1543 VDDD.n2200 VDDD.t1319 63.3219
R1544 VDDD.n2211 VDDD.t781 63.3219
R1545 VDDD.n2214 VDDD.t783 63.3219
R1546 VDDD.n2225 VDDD.t1347 63.3219
R1547 VDDD.n2228 VDDD.t1063 63.3219
R1548 VDDD.n2239 VDDD.t625 63.3219
R1549 VDDD.n2242 VDDD.t293 63.3219
R1550 VDDD.n2253 VDDD.t777 63.3219
R1551 VDDD.n2256 VDDD.t180 63.3219
R1552 VDDD.n2161 VDDD.t869 63.3219
R1553 VDDD.n1895 VDDD.t304 63.3219
R1554 VDDD.n1905 VDDD.t1415 63.3219
R1555 VDDD.n1908 VDDD.t1200 63.3219
R1556 VDDD.n1919 VDDD.t11 63.3219
R1557 VDDD.n1922 VDDD.t206 63.3219
R1558 VDDD.n1933 VDDD.t1413 63.3219
R1559 VDDD.n1936 VDDD.t896 63.3219
R1560 VDDD.n1947 VDDD.t13 63.3219
R1561 VDDD.n1950 VDDD.t1198 63.3219
R1562 VDDD.n1961 VDDD.t1323 63.3219
R1563 VDDD.n1964 VDDD.t1417 63.3219
R1564 VDDD.n1382 VDDD.t266 63.3219
R1565 VDDD.n1385 VDDD.t971 63.3219
R1566 VDDD.n1396 VDDD.t483 63.3219
R1567 VDDD.n1399 VDDD.t1072 63.3219
R1568 VDDD.n1410 VDDD.t314 63.3219
R1569 VDDD.n1413 VDDD.t618 63.3219
R1570 VDDD.n1424 VDDD.t1271 63.3219
R1571 VDDD.n1427 VDDD.t116 63.3219
R1572 VDDD.n1438 VDDD.t822 63.3219
R1573 VDDD.n1441 VDDD.t170 63.3219
R1574 VDDD.n1815 VDDD.t637 63.3219
R1575 VDDD.n1316 VDDD.t969 63.3219
R1576 VDDD.n1326 VDDD.t1301 63.3219
R1577 VDDD.n1329 VDDD.t1273 63.3219
R1578 VDDD.n1340 VDDD.t545 63.3219
R1579 VDDD.n1343 VDDD.t633 63.3219
R1580 VDDD.n1354 VDDD.t1303 63.3219
R1581 VDDD.n1357 VDDD.t850 63.3219
R1582 VDDD.n1368 VDDD.t908 63.3219
R1583 VDDD.n1371 VDDD.t516 63.3219
R1584 VDDD.n1085 VDDD.t627 63.3219
R1585 VDDD.n1082 VDDD.t1325 63.3219
R1586 VDDD.n1079 VDDD.t373 63.3219
R1587 VDDD.n1076 VDDD.t1411 63.3219
R1588 VDDD.n1068 VDDD.t1407 63.3219
R1589 VDDD.n1065 VDDD.t1321 63.3219
R1590 VDDD.n1062 VDDD.t1409 63.3219
R1591 VDDD.n1059 VDDD.t178 63.3219
R1592 VDDD.n1051 VDDD.t176 63.3219
R1593 VDDD.n1048 VDDD.t1059 63.3219
R1594 VDDD.n1045 VDDD.t894 63.3219
R1595 VDDD.n1042 VDDD.t1061 63.3219
R1596 VDDD.n1034 VDDD.t779 63.3219
R1597 VDDD.n1031 VDDD.t200 63.3219
R1598 VDDD.n1028 VDDD.t297 63.3219
R1599 VDDD.n1025 VDDD.t202 63.3219
R1600 VDDD.n1017 VDDD.t1419 63.3219
R1601 VDDD.n1277 VDDD.t204 63.3219
R1602 VDDD.n1285 VDDD.t1345 63.3219
R1603 VDDD.n1292 VDDD.t1202 63.3219
R1604 VDDD VDDD.t1390 52.0323
R1605 VDDD VDDD.t223 52.0323
R1606 VDDD VDDD.t1434 52.0323
R1607 VDDD VDDD.t1340 52.0323
R1608 VDDD VDDD.t1392 52.0323
R1609 VDDD.n272 VDDD.n271 43.1829
R1610 VDDD.n1005 VDDD.n1004 43.1829
R1611 VDDD.n294 VDDD.t126 41.5552
R1612 VDDD.n294 VDDD.t976 41.5552
R1613 VDDD.n247 VDDD.t807 41.5552
R1614 VDDD.n247 VDDD.t85 41.5552
R1615 VDDD.n363 VDDD.t834 41.5552
R1616 VDDD.n363 VDDD.t668 41.5552
R1617 VDDD.n222 VDDD.t59 41.5552
R1618 VDDD.n222 VDDD.t1292 41.5552
R1619 VDDD.n432 VDDD.t761 41.5552
R1620 VDDD.n432 VDDD.t3 41.5552
R1621 VDDD.n197 VDDD.t1404 41.5552
R1622 VDDD.n197 VDDD.t538 41.5552
R1623 VDDD.n501 VDDD.t210 41.5552
R1624 VDDD.n501 VDDD.t132 41.5552
R1625 VDDD.n172 VDDD.t153 41.5552
R1626 VDDD.n172 VDDD.t984 41.5552
R1627 VDDD.n570 VDDD.t1103 41.5552
R1628 VDDD.n570 VDDD.t645 41.5552
R1629 VDDD.n147 VDDD.t20 41.5552
R1630 VDDD.n147 VDDD.t285 41.5552
R1631 VDDD.n669 VDDD.t949 41.5552
R1632 VDDD.n669 VDDD.t283 41.5552
R1633 VDDD.n110 VDDD.t1175 41.5552
R1634 VDDD.n110 VDDD.t918 41.5552
R1635 VDDD.n738 VDDD.t275 41.5552
R1636 VDDD.n738 VDDD.t242 41.5552
R1637 VDDD.n85 VDDD.t1002 41.5552
R1638 VDDD.n85 VDDD.t718 41.5552
R1639 VDDD.n807 VDDD.t753 41.5552
R1640 VDDD.n807 VDDD.t536 41.5552
R1641 VDDD.n60 VDDD.t309 41.5552
R1642 VDDD.n60 VDDD.t5 41.5552
R1643 VDDD.n876 VDDD.t592 41.5552
R1644 VDDD.n876 VDDD.t1288 41.5552
R1645 VDDD.n35 VDDD.t774 41.5552
R1646 VDDD.n35 VDDD.t854 41.5552
R1647 VDDD.n945 VDDD.t7 41.5552
R1648 VDDD.n945 VDDD.t1132 41.5552
R1649 VDDD.n10 VDDD.t923 41.5552
R1650 VDDD.n10 VDDD.t978 41.5552
R1651 VDDD.n2179 VDDD.t1162 41.5552
R1652 VDDD.n2179 VDDD.t1026 41.5552
R1653 VDDD.n2192 VDDD.t974 41.5552
R1654 VDDD.n2192 VDDD.t343 41.5552
R1655 VDDD.n2206 VDDD.t659 41.5552
R1656 VDDD.n2206 VDDD.t345 41.5552
R1657 VDDD.n2220 VDDD.t857 41.5552
R1658 VDDD.n2220 VDDD.t1020 41.5552
R1659 VDDD.n2234 VDDD.t354 41.5552
R1660 VDDD.n2234 VDDD.t1117 41.5552
R1661 VDDD.n2248 VDDD.t1206 41.5552
R1662 VDDD.n2248 VDDD.t341 41.5552
R1663 VDDD.n1887 VDDD.t1286 41.5552
R1664 VDDD.n1887 VDDD.t1050 41.5552
R1665 VDDD.n1900 VDDD.t395 41.5552
R1666 VDDD.n1900 VDDD.t568 41.5552
R1667 VDDD.n1914 VDDD.t844 41.5552
R1668 VDDD.n1914 VDDD.t339 41.5552
R1669 VDDD.n1928 VDDD.t511 41.5552
R1670 VDDD.n1928 VDDD.t1018 41.5552
R1671 VDDD.n1942 VDDD.t359 41.5552
R1672 VDDD.n1942 VDDD.t1113 41.5552
R1673 VDDD.n1956 VDDD.t250 41.5552
R1674 VDDD.n1956 VDDD.t566 41.5552
R1675 VDDD.n1376 VDDD.t1052 41.5552
R1676 VDDD.n1376 VDDD.t441 41.5552
R1677 VDDD.n1390 VDDD.t830 41.5552
R1678 VDDD.n1390 VDDD.t1426 41.5552
R1679 VDDD.n1404 VDDD.t1115 41.5552
R1680 VDDD.n1404 VDDD.t246 41.5552
R1681 VDDD.n1418 VDDD.t826 41.5552
R1682 VDDD.n1418 VDDD.t1006 41.5552
R1683 VDDD.n1432 VDDD.t694 41.5552
R1684 VDDD.n1432 VDDD.t597 41.5552
R1685 VDDD.n1308 VDDD.t365 41.5552
R1686 VDDD.n1308 VDDD.t1054 41.5552
R1687 VDDD.n1321 VDDD.t31 41.5552
R1688 VDDD.n1321 VDDD.t1022 41.5552
R1689 VDDD.n1335 VDDD.t122 41.5552
R1690 VDDD.n1335 VDDD.t828 41.5552
R1691 VDDD.n1349 VDDD.t368 41.5552
R1692 VDDD.n1349 VDDD.t1024 41.5552
R1693 VDDD.n1363 VDDD.t1260 41.5552
R1694 VDDD.n1363 VDDD.t1048 41.5552
R1695 VDDD.n1010 VDDD.t71 41.5552
R1696 VDDD.n1010 VDDD.t69 41.5552
R1697 VDDD.n1088 VDDD.t1391 41.5552
R1698 VDDD.n1088 VDDD.t168 41.5552
R1699 VDDD.n1073 VDDD.t884 41.5552
R1700 VDDD.n1073 VDDD.t1153 41.5552
R1701 VDDD.n1071 VDDD.t224 41.5552
R1702 VDDD.n1071 VDDD.t766 41.5552
R1703 VDDD.n1056 VDDD.t758 41.5552
R1704 VDDD.n1056 VDDD.t1439 41.5552
R1705 VDDD.n1054 VDDD.t1435 41.5552
R1706 VDDD.n1054 VDDD.t446 41.5552
R1707 VDDD.n1039 VDDD.t426 41.5552
R1708 VDDD.n1039 VDDD.t1437 41.5552
R1709 VDDD.n1037 VDDD.t1341 41.5552
R1710 VDDD.n1037 VDDD.t1149 41.5552
R1711 VDDD.n1022 VDDD.t940 41.5552
R1712 VDDD.n1022 VDDD.t67 41.5552
R1713 VDDD.n1020 VDDD.t1393 41.5552
R1714 VDDD.n1020 VDDD.t1178 41.5552
R1715 VDDD.n1841 VDDD.n1840 38.777
R1716 VDDD.n1840 VDDD.n1833 38.777
R1717 VDDD.n1833 VDDD.n1831 38.777
R1718 VDDD.n1841 VDDD.n1831 38.777
R1719 VDDD.n1979 VDDD.n1978 38.777
R1720 VDDD.n1978 VDDD.n1971 38.777
R1721 VDDD.n1971 VDDD.n1969 38.777
R1722 VDDD.n1979 VDDD.n1969 38.777
R1723 VDDD.n2271 VDDD.n2270 38.777
R1724 VDDD.n2270 VDDD.n2263 38.777
R1725 VDDD.n2263 VDDD.n2261 38.777
R1726 VDDD.n2271 VDDD.n2261 38.777
R1727 VDDD.n1652 VDDD.n1642 38.777
R1728 VDDD.n1644 VDDD.n1642 38.777
R1729 VDDD.n1652 VDDD.n1651 38.777
R1730 VDDD.n1651 VDDD.n1644 38.777
R1731 VDDD.n1665 VDDD.n1655 38.777
R1732 VDDD.n1657 VDDD.n1655 38.777
R1733 VDDD.n1665 VDDD.n1664 38.777
R1734 VDDD.n1664 VDDD.n1657 38.777
R1735 VDDD.n1093 VDDD.n1092 38.777
R1736 VDDD.n1102 VDDD.n1093 38.777
R1737 VDDD.n1101 VDDD.n1092 38.777
R1738 VDDD.n1102 VDDD.n1101 38.777
R1739 VDDD.n278 VDDD.n266 34.6358
R1740 VDDD.n274 VDDD.n273 34.6358
R1741 VDDD.n282 VDDD.n281 34.6358
R1742 VDDD.n293 VDDD.n260 34.6358
R1743 VDDD.n296 VDDD.n258 34.6358
R1744 VDDD.n306 VDDD.n256 34.6358
R1745 VDDD.n302 VDDD.n256 34.6358
R1746 VDDD.n302 VDDD.n301 34.6358
R1747 VDDD.n310 VDDD.n309 34.6358
R1748 VDDD.n316 VDDD.n315 34.6358
R1749 VDDD.n315 VDDD.n314 34.6358
R1750 VDDD.n333 VDDD.n332 34.6358
R1751 VDDD.n340 VDDD.n339 34.6358
R1752 VDDD.n339 VDDD.n338 34.6358
R1753 VDDD.n338 VDDD.n245 34.6358
R1754 VDDD.n344 VDDD.n241 34.6358
R1755 VDDD.n350 VDDD.n239 34.6358
R1756 VDDD.n346 VDDD.n239 34.6358
R1757 VDDD.n365 VDDD.n233 34.6358
R1758 VDDD.n375 VDDD.n231 34.6358
R1759 VDDD.n371 VDDD.n231 34.6358
R1760 VDDD.n371 VDDD.n370 34.6358
R1761 VDDD.n379 VDDD.n378 34.6358
R1762 VDDD.n385 VDDD.n384 34.6358
R1763 VDDD.n384 VDDD.n383 34.6358
R1764 VDDD.n402 VDDD.n401 34.6358
R1765 VDDD.n409 VDDD.n408 34.6358
R1766 VDDD.n408 VDDD.n407 34.6358
R1767 VDDD.n407 VDDD.n220 34.6358
R1768 VDDD.n413 VDDD.n216 34.6358
R1769 VDDD.n419 VDDD.n214 34.6358
R1770 VDDD.n415 VDDD.n214 34.6358
R1771 VDDD.n434 VDDD.n208 34.6358
R1772 VDDD.n444 VDDD.n206 34.6358
R1773 VDDD.n440 VDDD.n206 34.6358
R1774 VDDD.n440 VDDD.n439 34.6358
R1775 VDDD.n448 VDDD.n447 34.6358
R1776 VDDD.n454 VDDD.n453 34.6358
R1777 VDDD.n453 VDDD.n452 34.6358
R1778 VDDD.n471 VDDD.n470 34.6358
R1779 VDDD.n478 VDDD.n477 34.6358
R1780 VDDD.n477 VDDD.n476 34.6358
R1781 VDDD.n476 VDDD.n195 34.6358
R1782 VDDD.n482 VDDD.n191 34.6358
R1783 VDDD.n488 VDDD.n189 34.6358
R1784 VDDD.n484 VDDD.n189 34.6358
R1785 VDDD.n503 VDDD.n183 34.6358
R1786 VDDD.n513 VDDD.n181 34.6358
R1787 VDDD.n509 VDDD.n181 34.6358
R1788 VDDD.n509 VDDD.n508 34.6358
R1789 VDDD.n517 VDDD.n516 34.6358
R1790 VDDD.n523 VDDD.n522 34.6358
R1791 VDDD.n522 VDDD.n521 34.6358
R1792 VDDD.n540 VDDD.n539 34.6358
R1793 VDDD.n547 VDDD.n546 34.6358
R1794 VDDD.n546 VDDD.n545 34.6358
R1795 VDDD.n545 VDDD.n170 34.6358
R1796 VDDD.n551 VDDD.n166 34.6358
R1797 VDDD.n557 VDDD.n164 34.6358
R1798 VDDD.n553 VDDD.n164 34.6358
R1799 VDDD.n572 VDDD.n158 34.6358
R1800 VDDD.n582 VDDD.n156 34.6358
R1801 VDDD.n578 VDDD.n156 34.6358
R1802 VDDD.n578 VDDD.n577 34.6358
R1803 VDDD.n586 VDDD.n585 34.6358
R1804 VDDD.n592 VDDD.n591 34.6358
R1805 VDDD.n591 VDDD.n590 34.6358
R1806 VDDD.n609 VDDD.n608 34.6358
R1807 VDDD.n616 VDDD.n615 34.6358
R1808 VDDD.n615 VDDD.n614 34.6358
R1809 VDDD.n614 VDDD.n145 34.6358
R1810 VDDD.n620 VDDD.n141 34.6358
R1811 VDDD.n626 VDDD.n139 34.6358
R1812 VDDD.n622 VDDD.n139 34.6358
R1813 VDDD.n649 VDDD.n648 34.6358
R1814 VDDD.n650 VDDD.n649 34.6358
R1815 VDDD.n655 VDDD.n654 34.6358
R1816 VDDD.n658 VDDD.n127 34.6358
R1817 VDDD.n662 VDDD.n127 34.6358
R1818 VDDD.n663 VDDD.n662 34.6358
R1819 VDDD.n668 VDDD.n125 34.6358
R1820 VDDD.n684 VDDD.n683 34.6358
R1821 VDDD.n684 VDDD.n118 34.6358
R1822 VDDD.n690 VDDD.n689 34.6358
R1823 VDDD.n694 VDDD.n693 34.6358
R1824 VDDD.n695 VDDD.n694 34.6358
R1825 VDDD.n695 VDDD.n113 34.6358
R1826 VDDD.n701 VDDD.n700 34.6358
R1827 VDDD.n718 VDDD.n717 34.6358
R1828 VDDD.n719 VDDD.n718 34.6358
R1829 VDDD.n724 VDDD.n723 34.6358
R1830 VDDD.n727 VDDD.n102 34.6358
R1831 VDDD.n731 VDDD.n102 34.6358
R1832 VDDD.n732 VDDD.n731 34.6358
R1833 VDDD.n737 VDDD.n100 34.6358
R1834 VDDD.n753 VDDD.n752 34.6358
R1835 VDDD.n753 VDDD.n93 34.6358
R1836 VDDD.n759 VDDD.n758 34.6358
R1837 VDDD.n763 VDDD.n762 34.6358
R1838 VDDD.n764 VDDD.n763 34.6358
R1839 VDDD.n764 VDDD.n88 34.6358
R1840 VDDD.n770 VDDD.n769 34.6358
R1841 VDDD.n787 VDDD.n786 34.6358
R1842 VDDD.n788 VDDD.n787 34.6358
R1843 VDDD.n793 VDDD.n792 34.6358
R1844 VDDD.n796 VDDD.n77 34.6358
R1845 VDDD.n800 VDDD.n77 34.6358
R1846 VDDD.n801 VDDD.n800 34.6358
R1847 VDDD.n806 VDDD.n75 34.6358
R1848 VDDD.n822 VDDD.n821 34.6358
R1849 VDDD.n822 VDDD.n68 34.6358
R1850 VDDD.n828 VDDD.n827 34.6358
R1851 VDDD.n832 VDDD.n831 34.6358
R1852 VDDD.n833 VDDD.n832 34.6358
R1853 VDDD.n833 VDDD.n63 34.6358
R1854 VDDD.n839 VDDD.n838 34.6358
R1855 VDDD.n856 VDDD.n855 34.6358
R1856 VDDD.n857 VDDD.n856 34.6358
R1857 VDDD.n862 VDDD.n861 34.6358
R1858 VDDD.n865 VDDD.n52 34.6358
R1859 VDDD.n869 VDDD.n52 34.6358
R1860 VDDD.n870 VDDD.n869 34.6358
R1861 VDDD.n875 VDDD.n50 34.6358
R1862 VDDD.n891 VDDD.n890 34.6358
R1863 VDDD.n891 VDDD.n43 34.6358
R1864 VDDD.n897 VDDD.n896 34.6358
R1865 VDDD.n901 VDDD.n900 34.6358
R1866 VDDD.n902 VDDD.n901 34.6358
R1867 VDDD.n902 VDDD.n38 34.6358
R1868 VDDD.n908 VDDD.n907 34.6358
R1869 VDDD.n925 VDDD.n924 34.6358
R1870 VDDD.n926 VDDD.n925 34.6358
R1871 VDDD.n931 VDDD.n930 34.6358
R1872 VDDD.n934 VDDD.n27 34.6358
R1873 VDDD.n938 VDDD.n27 34.6358
R1874 VDDD.n939 VDDD.n938 34.6358
R1875 VDDD.n944 VDDD.n25 34.6358
R1876 VDDD.n960 VDDD.n959 34.6358
R1877 VDDD.n960 VDDD.n18 34.6358
R1878 VDDD.n966 VDDD.n965 34.6358
R1879 VDDD.n970 VDDD.n969 34.6358
R1880 VDDD.n971 VDDD.n970 34.6358
R1881 VDDD.n971 VDDD.n13 34.6358
R1882 VDDD.n977 VDDD.n976 34.6358
R1883 VDDD.n982 VDDD.n981 34.6358
R1884 VDDD.n995 VDDD.n7 34.6358
R1885 VDDD.n999 VDDD.n998 34.6358
R1886 VDDD.n1003 VDDD.n1002 34.6358
R1887 VDDD.n2470 VDDD.n2469 34.6358
R1888 VDDD.n2463 VDDD.n2182 34.6358
R1889 VDDD.n2464 VDDD.n2463 34.6358
R1890 VDDD.n2465 VDDD.n2464 34.6358
R1891 VDDD.n2459 VDDD.n2456 34.6358
R1892 VDDD.n2450 VDDD.n2185 34.6358
R1893 VDDD.n2454 VDDD.n2185 34.6358
R1894 VDDD.n2437 VDDD.n2193 34.6358
R1895 VDDD.n2427 VDDD.n2195 34.6358
R1896 VDDD.n2431 VDDD.n2195 34.6358
R1897 VDDD.n2432 VDDD.n2431 34.6358
R1898 VDDD.n2425 VDDD.n2424 34.6358
R1899 VDDD.n2419 VDDD.n2418 34.6358
R1900 VDDD.n2420 VDDD.n2419 34.6358
R1901 VDDD.n2404 VDDD.n2207 34.6358
R1902 VDDD.n2394 VDDD.n2209 34.6358
R1903 VDDD.n2398 VDDD.n2209 34.6358
R1904 VDDD.n2399 VDDD.n2398 34.6358
R1905 VDDD.n2392 VDDD.n2391 34.6358
R1906 VDDD.n2386 VDDD.n2385 34.6358
R1907 VDDD.n2387 VDDD.n2386 34.6358
R1908 VDDD.n2371 VDDD.n2221 34.6358
R1909 VDDD.n2361 VDDD.n2223 34.6358
R1910 VDDD.n2365 VDDD.n2223 34.6358
R1911 VDDD.n2366 VDDD.n2365 34.6358
R1912 VDDD.n2359 VDDD.n2358 34.6358
R1913 VDDD.n2353 VDDD.n2352 34.6358
R1914 VDDD.n2354 VDDD.n2353 34.6358
R1915 VDDD.n2338 VDDD.n2235 34.6358
R1916 VDDD.n2328 VDDD.n2237 34.6358
R1917 VDDD.n2332 VDDD.n2237 34.6358
R1918 VDDD.n2333 VDDD.n2332 34.6358
R1919 VDDD.n2326 VDDD.n2325 34.6358
R1920 VDDD.n2320 VDDD.n2319 34.6358
R1921 VDDD.n2321 VDDD.n2320 34.6358
R1922 VDDD.n2305 VDDD.n2249 34.6358
R1923 VDDD.n2295 VDDD.n2251 34.6358
R1924 VDDD.n2299 VDDD.n2251 34.6358
R1925 VDDD.n2300 VDDD.n2299 34.6358
R1926 VDDD.n2293 VDDD.n2292 34.6358
R1927 VDDD.n2287 VDDD.n2286 34.6358
R1928 VDDD.n2288 VDDD.n2287 34.6358
R1929 VDDD.n1875 VDDD.n1846 34.6358
R1930 VDDD.n1879 VDDD.n1846 34.6358
R1931 VDDD.n1859 VDDD.n1858 34.6358
R1932 VDDD.n1867 VDDD.n1851 34.6358
R1933 VDDD.n1870 VDDD.n1869 34.6358
R1934 VDDD.n2174 VDDD.n2173 34.6358
R1935 VDDD.n2167 VDDD.n1890 34.6358
R1936 VDDD.n2168 VDDD.n2167 34.6358
R1937 VDDD.n2169 VDDD.n2168 34.6358
R1938 VDDD.n2163 VDDD.n2160 34.6358
R1939 VDDD.n2154 VDDD.n1893 34.6358
R1940 VDDD.n2158 VDDD.n1893 34.6358
R1941 VDDD.n2141 VDDD.n1901 34.6358
R1942 VDDD.n2131 VDDD.n1903 34.6358
R1943 VDDD.n2135 VDDD.n1903 34.6358
R1944 VDDD.n2136 VDDD.n2135 34.6358
R1945 VDDD.n2129 VDDD.n2128 34.6358
R1946 VDDD.n2123 VDDD.n2122 34.6358
R1947 VDDD.n2124 VDDD.n2123 34.6358
R1948 VDDD.n2108 VDDD.n1915 34.6358
R1949 VDDD.n2098 VDDD.n1917 34.6358
R1950 VDDD.n2102 VDDD.n1917 34.6358
R1951 VDDD.n2103 VDDD.n2102 34.6358
R1952 VDDD.n2096 VDDD.n2095 34.6358
R1953 VDDD.n2090 VDDD.n2089 34.6358
R1954 VDDD.n2091 VDDD.n2090 34.6358
R1955 VDDD.n2075 VDDD.n1929 34.6358
R1956 VDDD.n2065 VDDD.n1931 34.6358
R1957 VDDD.n2069 VDDD.n1931 34.6358
R1958 VDDD.n2070 VDDD.n2069 34.6358
R1959 VDDD.n2063 VDDD.n2062 34.6358
R1960 VDDD.n2057 VDDD.n2056 34.6358
R1961 VDDD.n2058 VDDD.n2057 34.6358
R1962 VDDD.n2042 VDDD.n1943 34.6358
R1963 VDDD.n2032 VDDD.n1945 34.6358
R1964 VDDD.n2036 VDDD.n1945 34.6358
R1965 VDDD.n2037 VDDD.n2036 34.6358
R1966 VDDD.n2030 VDDD.n2029 34.6358
R1967 VDDD.n2024 VDDD.n2023 34.6358
R1968 VDDD.n2025 VDDD.n2024 34.6358
R1969 VDDD.n2009 VDDD.n1957 34.6358
R1970 VDDD.n1999 VDDD.n1959 34.6358
R1971 VDDD.n2003 VDDD.n1959 34.6358
R1972 VDDD.n2004 VDDD.n2003 34.6358
R1973 VDDD.n1997 VDDD.n1996 34.6358
R1974 VDDD.n1991 VDDD.n1990 34.6358
R1975 VDDD.n1992 VDDD.n1991 34.6358
R1976 VDDD.n1638 VDDD.n1378 34.6358
R1977 VDDD.n1633 VDDD.n1632 34.6358
R1978 VDDD.n1632 VDDD.n1380 34.6358
R1979 VDDD.n1628 VDDD.n1380 34.6358
R1980 VDDD.n1626 VDDD.n1625 34.6358
R1981 VDDD.n1621 VDDD.n1620 34.6358
R1982 VDDD.n1620 VDDD.n1619 34.6358
R1983 VDDD.n1605 VDDD.n1392 34.6358
R1984 VDDD.n1600 VDDD.n1599 34.6358
R1985 VDDD.n1599 VDDD.n1394 34.6358
R1986 VDDD.n1595 VDDD.n1394 34.6358
R1987 VDDD.n1593 VDDD.n1592 34.6358
R1988 VDDD.n1588 VDDD.n1587 34.6358
R1989 VDDD.n1587 VDDD.n1586 34.6358
R1990 VDDD.n1572 VDDD.n1406 34.6358
R1991 VDDD.n1567 VDDD.n1566 34.6358
R1992 VDDD.n1566 VDDD.n1408 34.6358
R1993 VDDD.n1562 VDDD.n1408 34.6358
R1994 VDDD.n1560 VDDD.n1559 34.6358
R1995 VDDD.n1555 VDDD.n1554 34.6358
R1996 VDDD.n1554 VDDD.n1553 34.6358
R1997 VDDD.n1539 VDDD.n1420 34.6358
R1998 VDDD.n1534 VDDD.n1533 34.6358
R1999 VDDD.n1533 VDDD.n1422 34.6358
R2000 VDDD.n1529 VDDD.n1422 34.6358
R2001 VDDD.n1527 VDDD.n1526 34.6358
R2002 VDDD.n1522 VDDD.n1521 34.6358
R2003 VDDD.n1521 VDDD.n1520 34.6358
R2004 VDDD.n1506 VDDD.n1434 34.6358
R2005 VDDD.n1501 VDDD.n1500 34.6358
R2006 VDDD.n1500 VDDD.n1436 34.6358
R2007 VDDD.n1496 VDDD.n1436 34.6358
R2008 VDDD.n1494 VDDD.n1493 34.6358
R2009 VDDD.n1489 VDDD.n1488 34.6358
R2010 VDDD.n1488 VDDD.n1487 34.6358
R2011 VDDD.n1473 VDDD.n1447 34.6358
R2012 VDDD.n1469 VDDD.n1468 34.6358
R2013 VDDD.n1466 VDDD.n1452 34.6358
R2014 VDDD.n1828 VDDD.n1827 34.6358
R2015 VDDD.n1821 VDDD.n1311 34.6358
R2016 VDDD.n1822 VDDD.n1821 34.6358
R2017 VDDD.n1823 VDDD.n1822 34.6358
R2018 VDDD.n1817 VDDD.n1814 34.6358
R2019 VDDD.n1808 VDDD.n1314 34.6358
R2020 VDDD.n1812 VDDD.n1314 34.6358
R2021 VDDD.n1795 VDDD.n1322 34.6358
R2022 VDDD.n1785 VDDD.n1324 34.6358
R2023 VDDD.n1789 VDDD.n1324 34.6358
R2024 VDDD.n1790 VDDD.n1789 34.6358
R2025 VDDD.n1783 VDDD.n1782 34.6358
R2026 VDDD.n1777 VDDD.n1776 34.6358
R2027 VDDD.n1778 VDDD.n1777 34.6358
R2028 VDDD.n1762 VDDD.n1336 34.6358
R2029 VDDD.n1752 VDDD.n1338 34.6358
R2030 VDDD.n1756 VDDD.n1338 34.6358
R2031 VDDD.n1757 VDDD.n1756 34.6358
R2032 VDDD.n1750 VDDD.n1749 34.6358
R2033 VDDD.n1744 VDDD.n1743 34.6358
R2034 VDDD.n1745 VDDD.n1744 34.6358
R2035 VDDD.n1729 VDDD.n1350 34.6358
R2036 VDDD.n1719 VDDD.n1352 34.6358
R2037 VDDD.n1723 VDDD.n1352 34.6358
R2038 VDDD.n1724 VDDD.n1723 34.6358
R2039 VDDD.n1717 VDDD.n1716 34.6358
R2040 VDDD.n1711 VDDD.n1710 34.6358
R2041 VDDD.n1712 VDDD.n1711 34.6358
R2042 VDDD.n1696 VDDD.n1364 34.6358
R2043 VDDD.n1686 VDDD.n1366 34.6358
R2044 VDDD.n1690 VDDD.n1366 34.6358
R2045 VDDD.n1691 VDDD.n1690 34.6358
R2046 VDDD.n1684 VDDD.n1683 34.6358
R2047 VDDD.n1678 VDDD.n1677 34.6358
R2048 VDDD.n1679 VDDD.n1678 34.6358
R2049 VDDD.n1110 VDDD.n1106 34.6358
R2050 VDDD.n1114 VDDD.n1090 34.6358
R2051 VDDD.n1128 VDDD.n1127 34.6358
R2052 VDDD.n1129 VDDD.n1128 34.6358
R2053 VDDD.n1138 VDDD.n1137 34.6358
R2054 VDDD.n1139 VDDD.n1138 34.6358
R2055 VDDD.n1165 VDDD.n1164 34.6358
R2056 VDDD.n1166 VDDD.n1165 34.6358
R2057 VDDD.n1175 VDDD.n1174 34.6358
R2058 VDDD.n1176 VDDD.n1175 34.6358
R2059 VDDD.n1202 VDDD.n1201 34.6358
R2060 VDDD.n1203 VDDD.n1202 34.6358
R2061 VDDD.n1212 VDDD.n1211 34.6358
R2062 VDDD.n1213 VDDD.n1212 34.6358
R2063 VDDD.n1239 VDDD.n1238 34.6358
R2064 VDDD.n1240 VDDD.n1239 34.6358
R2065 VDDD.n1249 VDDD.n1248 34.6358
R2066 VDDD.n1250 VDDD.n1249 34.6358
R2067 VDDD.n1276 VDDD.n1275 34.6358
R2068 VDDD.n1279 VDDD.n1276 34.6358
R2069 VDDD.n1287 VDDD.n1013 34.6358
R2070 VDDD.n1291 VDDD.n1013 34.6358
R2071 VDDD.n1475 VDDD.n1474 33.8829
R2072 VDDD.n2478 VDDD 32.5497
R2073 VDDD.n301 VDDD.n300 32.377
R2074 VDDD.n334 VDDD.n245 32.377
R2075 VDDD.n370 VDDD.n369 32.377
R2076 VDDD.n403 VDDD.n220 32.377
R2077 VDDD.n439 VDDD.n438 32.377
R2078 VDDD.n472 VDDD.n195 32.377
R2079 VDDD.n508 VDDD.n507 32.377
R2080 VDDD.n541 VDDD.n170 32.377
R2081 VDDD.n577 VDDD.n576 32.377
R2082 VDDD.n610 VDDD.n145 32.377
R2083 VDDD.n664 VDDD.n663 32.377
R2084 VDDD.n699 VDDD.n113 32.377
R2085 VDDD.n733 VDDD.n732 32.377
R2086 VDDD.n768 VDDD.n88 32.377
R2087 VDDD.n802 VDDD.n801 32.377
R2088 VDDD.n837 VDDD.n63 32.377
R2089 VDDD.n871 VDDD.n870 32.377
R2090 VDDD.n906 VDDD.n38 32.377
R2091 VDDD.n940 VDDD.n939 32.377
R2092 VDDD.n975 VDDD.n13 32.377
R2093 VDDD.n2465 VDDD.n2180 32.377
R2094 VDDD.n2433 VDDD.n2432 32.377
R2095 VDDD.n2400 VDDD.n2399 32.377
R2096 VDDD.n2367 VDDD.n2366 32.377
R2097 VDDD.n2334 VDDD.n2333 32.377
R2098 VDDD.n2301 VDDD.n2300 32.377
R2099 VDDD.n2169 VDDD.n1888 32.377
R2100 VDDD.n2137 VDDD.n2136 32.377
R2101 VDDD.n2104 VDDD.n2103 32.377
R2102 VDDD.n2071 VDDD.n2070 32.377
R2103 VDDD.n2038 VDDD.n2037 32.377
R2104 VDDD.n2005 VDDD.n2004 32.377
R2105 VDDD.n1634 VDDD.n1633 32.377
R2106 VDDD.n1601 VDDD.n1600 32.377
R2107 VDDD.n1568 VDDD.n1567 32.377
R2108 VDDD.n1535 VDDD.n1534 32.377
R2109 VDDD.n1502 VDDD.n1501 32.377
R2110 VDDD.n1823 VDDD.n1309 32.377
R2111 VDDD.n1791 VDDD.n1790 32.377
R2112 VDDD.n1758 VDDD.n1757 32.377
R2113 VDDD.n1725 VDDD.n1724 32.377
R2114 VDDD.n1692 VDDD.n1691 32.377
R2115 VDDD.n287 VDDD.n262 32.0005
R2116 VDDD.n314 VDDD.n254 32.0005
R2117 VDDD.n346 VDDD.n345 32.0005
R2118 VDDD.n383 VDDD.n229 32.0005
R2119 VDDD.n415 VDDD.n414 32.0005
R2120 VDDD.n452 VDDD.n204 32.0005
R2121 VDDD.n484 VDDD.n483 32.0005
R2122 VDDD.n521 VDDD.n179 32.0005
R2123 VDDD.n553 VDDD.n552 32.0005
R2124 VDDD.n590 VDDD.n154 32.0005
R2125 VDDD.n622 VDDD.n621 32.0005
R2126 VDDD.n650 VDDD.n129 32.0005
R2127 VDDD.n688 VDDD.n118 32.0005
R2128 VDDD.n719 VDDD.n104 32.0005
R2129 VDDD.n757 VDDD.n93 32.0005
R2130 VDDD.n788 VDDD.n79 32.0005
R2131 VDDD.n826 VDDD.n68 32.0005
R2132 VDDD.n857 VDDD.n54 32.0005
R2133 VDDD.n895 VDDD.n43 32.0005
R2134 VDDD.n926 VDDD.n29 32.0005
R2135 VDDD.n964 VDDD.n18 32.0005
R2136 VDDD.n991 VDDD.n988 32.0005
R2137 VDDD.n2455 VDDD.n2454 32.0005
R2138 VDDD.n2420 VDDD.n2198 32.0005
R2139 VDDD.n2387 VDDD.n2212 32.0005
R2140 VDDD.n2354 VDDD.n2226 32.0005
R2141 VDDD.n2321 VDDD.n2240 32.0005
R2142 VDDD.n2288 VDDD.n2254 32.0005
R2143 VDDD.n1863 VDDD.n1862 32.0005
R2144 VDDD.n2159 VDDD.n2158 32.0005
R2145 VDDD.n2124 VDDD.n1906 32.0005
R2146 VDDD.n2091 VDDD.n1920 32.0005
R2147 VDDD.n2058 VDDD.n1934 32.0005
R2148 VDDD.n2025 VDDD.n1948 32.0005
R2149 VDDD.n1992 VDDD.n1962 32.0005
R2150 VDDD.n1621 VDDD.n1383 32.0005
R2151 VDDD.n1588 VDDD.n1397 32.0005
R2152 VDDD.n1555 VDDD.n1411 32.0005
R2153 VDDD.n1522 VDDD.n1425 32.0005
R2154 VDDD.n1489 VDDD.n1439 32.0005
R2155 VDDD.n1462 VDDD.n1461 32.0005
R2156 VDDD.n1813 VDDD.n1812 32.0005
R2157 VDDD.n1778 VDDD.n1327 32.0005
R2158 VDDD.n1745 VDDD.n1341 32.0005
R2159 VDDD.n1712 VDDD.n1355 32.0005
R2160 VDDD.n1679 VDDD.n1369 32.0005
R2161 VDDD.n1874 VDDD.n1873 31.2476
R2162 VDDD.n1863 VDDD.n1860 31.2476
R2163 VDDD.n1640 VDDD.n1639 30.7593
R2164 VDDD.n1123 VDDD.n1086 30.1181
R2165 VDDD.n1143 VDDD.n1077 30.1181
R2166 VDDD.n1160 VDDD.n1069 30.1181
R2167 VDDD.n1180 VDDD.n1060 30.1181
R2168 VDDD.n1197 VDDD.n1052 30.1181
R2169 VDDD.n1217 VDDD.n1043 30.1181
R2170 VDDD.n1234 VDDD.n1035 30.1181
R2171 VDDD.n1254 VDDD.n1026 30.1181
R2172 VDDD.n1271 VDDD.n1018 30.1181
R2173 VDDD.n1296 VDDD.n1293 30.1181
R2174 VDDD.n320 VDDD.n252 30.1181
R2175 VDDD.n353 VDDD.n352 30.1181
R2176 VDDD.n389 VDDD.n227 30.1181
R2177 VDDD.n422 VDDD.n421 30.1181
R2178 VDDD.n458 VDDD.n202 30.1181
R2179 VDDD.n491 VDDD.n490 30.1181
R2180 VDDD.n527 VDDD.n177 30.1181
R2181 VDDD.n560 VDDD.n559 30.1181
R2182 VDDD.n596 VDDD.n152 30.1181
R2183 VDDD.n629 VDDD.n628 30.1181
R2184 VDDD.n644 VDDD.n132 30.1181
R2185 VDDD.n682 VDDD.n120 30.1181
R2186 VDDD.n713 VDDD.n107 30.1181
R2187 VDDD.n751 VDDD.n95 30.1181
R2188 VDDD.n782 VDDD.n82 30.1181
R2189 VDDD.n820 VDDD.n70 30.1181
R2190 VDDD.n851 VDDD.n57 30.1181
R2191 VDDD.n889 VDDD.n45 30.1181
R2192 VDDD.n920 VDDD.n32 30.1181
R2193 VDDD.n958 VDDD.n20 30.1181
R2194 VDDD.n2449 VDDD.n2448 30.1181
R2195 VDDD.n2414 VDDD.n2201 30.1181
R2196 VDDD.n2381 VDDD.n2215 30.1181
R2197 VDDD.n2348 VDDD.n2229 30.1181
R2198 VDDD.n2315 VDDD.n2243 30.1181
R2199 VDDD.n2282 VDDD.n2257 30.1181
R2200 VDDD.n2153 VDDD.n2152 30.1181
R2201 VDDD.n2118 VDDD.n1909 30.1181
R2202 VDDD.n2085 VDDD.n1923 30.1181
R2203 VDDD.n2052 VDDD.n1937 30.1181
R2204 VDDD.n2019 VDDD.n1951 30.1181
R2205 VDDD.n1986 VDDD.n1965 30.1181
R2206 VDDD.n1615 VDDD.n1386 30.1181
R2207 VDDD.n1582 VDDD.n1400 30.1181
R2208 VDDD.n1549 VDDD.n1414 30.1181
R2209 VDDD.n1516 VDDD.n1428 30.1181
R2210 VDDD.n1483 VDDD.n1442 30.1181
R2211 VDDD.n1807 VDDD.n1806 30.1181
R2212 VDDD.n1772 VDDD.n1330 30.1181
R2213 VDDD.n1739 VDDD.n1344 30.1181
R2214 VDDD.n1706 VDDD.n1358 30.1181
R2215 VDDD.n1673 VDDD.n1372 30.1181
R2216 VDDD.n1855 VDDD.n1854 30.0041
R2217 VDDD.n1107 VDDD.t656 28.4453
R2218 VDDD.n1108 VDDD.t543 28.4453
R2219 VDDD.n274 VDDD.n269 27.8593
R2220 VDDD.n1002 VDDD.n5 27.8593
R2221 VDDD.n1450 VDDD.n1447 27.8593
R2222 VDDD.n328 VDDD.n327 27.4829
R2223 VDDD.n362 VDDD.n235 27.4829
R2224 VDDD.n397 VDDD.n396 27.4829
R2225 VDDD.n431 VDDD.n210 27.4829
R2226 VDDD.n466 VDDD.n465 27.4829
R2227 VDDD.n500 VDDD.n185 27.4829
R2228 VDDD.n535 VDDD.n534 27.4829
R2229 VDDD.n569 VDDD.n160 27.4829
R2230 VDDD.n604 VDDD.n603 27.4829
R2231 VDDD.n671 VDDD.n123 27.4829
R2232 VDDD.n706 VDDD.n705 27.4829
R2233 VDDD.n740 VDDD.n98 27.4829
R2234 VDDD.n775 VDDD.n774 27.4829
R2235 VDDD.n809 VDDD.n73 27.4829
R2236 VDDD.n844 VDDD.n843 27.4829
R2237 VDDD.n878 VDDD.n48 27.4829
R2238 VDDD.n913 VDDD.n912 27.4829
R2239 VDDD.n947 VDDD.n23 27.4829
R2240 VDDD.n2439 VDDD.n2190 27.4829
R2241 VDDD.n2406 VDDD.n2204 27.4829
R2242 VDDD.n2373 VDDD.n2218 27.4829
R2243 VDDD.n2340 VDDD.n2232 27.4829
R2244 VDDD.n2307 VDDD.n2246 27.4829
R2245 VDDD.n2274 VDDD.n2260 27.4829
R2246 VDDD.n2143 VDDD.n1898 27.4829
R2247 VDDD.n2110 VDDD.n1912 27.4829
R2248 VDDD.n2077 VDDD.n1926 27.4829
R2249 VDDD.n2044 VDDD.n1940 27.4829
R2250 VDDD.n2011 VDDD.n1954 27.4829
R2251 VDDD.n1607 VDDD.n1389 27.4829
R2252 VDDD.n1574 VDDD.n1403 27.4829
R2253 VDDD.n1541 VDDD.n1417 27.4829
R2254 VDDD.n1508 VDDD.n1431 27.4829
R2255 VDDD.n1797 VDDD.n1319 27.4829
R2256 VDDD.n1764 VDDD.n1333 27.4829
R2257 VDDD.n1731 VDDD.n1347 27.4829
R2258 VDDD.n1698 VDDD.n1361 27.4829
R2259 VDDD.n1475 VDDD.n1445 27.1064
R2260 VDDD.n1115 VDDD.n1114 27.1064
R2261 VDDD.n270 VDDD.t927 26.5955
R2262 VDDD.n270 VDDD.t925 26.5955
R2263 VDDD.n268 VDDD.t188 26.5955
R2264 VDDD.n268 VDDD.t666 26.5955
R2265 VDDD.n279 VDDD.t212 26.5955
R2266 VDDD.n279 VDDD.t886 26.5955
R2267 VDDD.n264 VDDD.t272 26.5955
R2268 VDDD.n264 VDDD.t186 26.5955
R2269 VDDD.n286 VDDD.t888 26.5955
R2270 VDDD.n286 VDDD.t411 26.5955
R2271 VDDD.n987 VDDD.t400 26.5955
R2272 VDDD.n987 VDDD.t402 26.5955
R2273 VDDD.n989 VDDD.t387 26.5955
R2274 VDDD.n989 VDDD.t391 26.5955
R2275 VDDD.n996 VDDD.t1455 26.5955
R2276 VDDD.n996 VDDD.t268 26.5955
R2277 VDDD.n4 VDDD.t389 26.5955
R2278 VDDD.n4 VDDD.t481 26.5955
R2279 VDDD.n3 VDDD.t287 26.5955
R2280 VDDD.n3 VDDD.t479 26.5955
R2281 VDDD.n1845 VDDD.t190 26.5955
R2282 VDDD.n1845 VDDD.t1004 26.5955
R2283 VDDD.n1850 VDDD.t474 26.5955
R2284 VDDD.n1850 VDDD.t226 26.5955
R2285 VDDD.n1861 VDDD.t1429 26.5955
R2286 VDDD.n1861 VDDD.t573 26.5955
R2287 VDDD.n1853 VDDD.t472 26.5955
R2288 VDDD.n1853 VDDD.t174 26.5955
R2289 VDDD.n1446 VDDD.t980 26.5955
R2290 VDDD.n1446 VDDD.t1421 26.5955
R2291 VDDD.n1449 VDDD.t423 26.5955
R2292 VDDD.n1449 VDDD.t1091 26.5955
R2293 VDDD.n1451 VDDD.t1441 26.5955
R2294 VDDD.n1451 VDDD.t1093 26.5955
R2295 VDDD.n1454 VDDD.t1447 26.5955
R2296 VDDD.n1454 VDDD.t1443 26.5955
R2297 VDDD.n1456 VDDD.t672 26.5955
R2298 VDDD.n1456 VDDD.t1449 26.5955
R2299 VDDD.n289 VDDD.n288 25.977
R2300 VDDD.n986 VDDD.n9 25.977
R2301 VDDD.n1868 VDDD.n1867 25.977
R2302 VDDD.n1460 VDDD.n1457 25.977
R2303 VDDD.n1882 VDDD.n1881 25.224
R2304 VDDD.n1883 VDDD.n1882 25.224
R2305 VDDD.n323 VDDD.n322 24.8476
R2306 VDDD.n357 VDDD.n356 24.8476
R2307 VDDD.n392 VDDD.n391 24.8476
R2308 VDDD.n426 VDDD.n425 24.8476
R2309 VDDD.n461 VDDD.n460 24.8476
R2310 VDDD.n495 VDDD.n494 24.8476
R2311 VDDD.n530 VDDD.n529 24.8476
R2312 VDDD.n564 VDDD.n563 24.8476
R2313 VDDD.n599 VDDD.n598 24.8476
R2314 VDDD.n633 VDDD.n136 24.8476
R2315 VDDD.n642 VDDD.n641 24.8476
R2316 VDDD.n678 VDDD.n676 24.8476
R2317 VDDD.n711 VDDD.n710 24.8476
R2318 VDDD.n747 VDDD.n745 24.8476
R2319 VDDD.n780 VDDD.n779 24.8476
R2320 VDDD.n816 VDDD.n814 24.8476
R2321 VDDD.n849 VDDD.n848 24.8476
R2322 VDDD.n885 VDDD.n883 24.8476
R2323 VDDD.n918 VDDD.n917 24.8476
R2324 VDDD.n954 VDDD.n952 24.8476
R2325 VDDD.n2445 VDDD.n2444 24.8476
R2326 VDDD.n2412 VDDD.n2411 24.8476
R2327 VDDD.n2379 VDDD.n2378 24.8476
R2328 VDDD.n2346 VDDD.n2345 24.8476
R2329 VDDD.n2313 VDDD.n2312 24.8476
R2330 VDDD.n2280 VDDD.n2279 24.8476
R2331 VDDD.n2149 VDDD.n2148 24.8476
R2332 VDDD.n2116 VDDD.n2115 24.8476
R2333 VDDD.n2083 VDDD.n2082 24.8476
R2334 VDDD.n2050 VDDD.n2049 24.8476
R2335 VDDD.n2017 VDDD.n2016 24.8476
R2336 VDDD.n1984 VDDD.n1983 24.8476
R2337 VDDD.n1613 VDDD.n1612 24.8476
R2338 VDDD.n1580 VDDD.n1579 24.8476
R2339 VDDD.n1547 VDDD.n1546 24.8476
R2340 VDDD.n1514 VDDD.n1513 24.8476
R2341 VDDD.n1481 VDDD.n1480 24.8476
R2342 VDDD.n1803 VDDD.n1802 24.8476
R2343 VDDD.n1770 VDDD.n1769 24.8476
R2344 VDDD.n1737 VDDD.n1736 24.8476
R2345 VDDD.n1704 VDDD.n1703 24.8476
R2346 VDDD.n1671 VDDD.n1670 24.8476
R2347 VDDD.n1120 VDDD.n1119 24.8476
R2348 VDDD.n1147 VDDD.n1146 24.8476
R2349 VDDD.n1157 VDDD.n1156 24.8476
R2350 VDDD.n1184 VDDD.n1183 24.8476
R2351 VDDD.n1194 VDDD.n1193 24.8476
R2352 VDDD.n1221 VDDD.n1220 24.8476
R2353 VDDD.n1231 VDDD.n1230 24.8476
R2354 VDDD.n1258 VDDD.n1257 24.8476
R2355 VDDD.n1268 VDDD.n1267 24.8476
R2356 VDDD.n1300 VDDD.n1011 24.8476
R2357 VDDD.n296 VDDD.n295 22.9652
R2358 VDDD.n327 VDDD.n249 22.9652
R2359 VDDD.n332 VDDD.n248 22.9652
R2360 VDDD.n358 VDDD.n235 22.9652
R2361 VDDD.n365 VDDD.n364 22.9652
R2362 VDDD.n396 VDDD.n224 22.9652
R2363 VDDD.n401 VDDD.n223 22.9652
R2364 VDDD.n427 VDDD.n210 22.9652
R2365 VDDD.n434 VDDD.n433 22.9652
R2366 VDDD.n465 VDDD.n199 22.9652
R2367 VDDD.n470 VDDD.n198 22.9652
R2368 VDDD.n496 VDDD.n185 22.9652
R2369 VDDD.n503 VDDD.n502 22.9652
R2370 VDDD.n534 VDDD.n174 22.9652
R2371 VDDD.n539 VDDD.n173 22.9652
R2372 VDDD.n565 VDDD.n160 22.9652
R2373 VDDD.n572 VDDD.n571 22.9652
R2374 VDDD.n603 VDDD.n149 22.9652
R2375 VDDD.n608 VDDD.n148 22.9652
R2376 VDDD.n635 VDDD.n634 22.9652
R2377 VDDD.n637 VDDD.n134 22.9652
R2378 VDDD.n670 VDDD.n668 22.9652
R2379 VDDD.n675 VDDD.n123 22.9652
R2380 VDDD.n701 VDDD.n111 22.9652
R2381 VDDD.n706 VDDD.n109 22.9652
R2382 VDDD.n739 VDDD.n737 22.9652
R2383 VDDD.n744 VDDD.n98 22.9652
R2384 VDDD.n770 VDDD.n86 22.9652
R2385 VDDD.n775 VDDD.n84 22.9652
R2386 VDDD.n808 VDDD.n806 22.9652
R2387 VDDD.n813 VDDD.n73 22.9652
R2388 VDDD.n839 VDDD.n61 22.9652
R2389 VDDD.n844 VDDD.n59 22.9652
R2390 VDDD.n877 VDDD.n875 22.9652
R2391 VDDD.n882 VDDD.n48 22.9652
R2392 VDDD.n908 VDDD.n36 22.9652
R2393 VDDD.n913 VDDD.n34 22.9652
R2394 VDDD.n946 VDDD.n944 22.9652
R2395 VDDD.n951 VDDD.n23 22.9652
R2396 VDDD.n977 VDDD.n11 22.9652
R2397 VDDD.n2471 VDDD.n2470 22.9652
R2398 VDDD.n2443 VDDD.n2190 22.9652
R2399 VDDD.n2438 VDDD.n2437 22.9652
R2400 VDDD.n2410 VDDD.n2204 22.9652
R2401 VDDD.n2405 VDDD.n2404 22.9652
R2402 VDDD.n2377 VDDD.n2218 22.9652
R2403 VDDD.n2372 VDDD.n2371 22.9652
R2404 VDDD.n2344 VDDD.n2232 22.9652
R2405 VDDD.n2339 VDDD.n2338 22.9652
R2406 VDDD.n2311 VDDD.n2246 22.9652
R2407 VDDD.n2306 VDDD.n2305 22.9652
R2408 VDDD.n2278 VDDD.n2260 22.9652
R2409 VDDD.n2175 VDDD.n2174 22.9652
R2410 VDDD.n2147 VDDD.n1898 22.9652
R2411 VDDD.n2142 VDDD.n2141 22.9652
R2412 VDDD.n2114 VDDD.n1912 22.9652
R2413 VDDD.n2109 VDDD.n2108 22.9652
R2414 VDDD.n2081 VDDD.n1926 22.9652
R2415 VDDD.n2076 VDDD.n2075 22.9652
R2416 VDDD.n2048 VDDD.n1940 22.9652
R2417 VDDD.n2043 VDDD.n2042 22.9652
R2418 VDDD.n2015 VDDD.n1954 22.9652
R2419 VDDD.n2010 VDDD.n2009 22.9652
R2420 VDDD.n1982 VDDD.n1968 22.9652
R2421 VDDD.n1639 VDDD.n1638 22.9652
R2422 VDDD.n1611 VDDD.n1389 22.9652
R2423 VDDD.n1606 VDDD.n1605 22.9652
R2424 VDDD.n1578 VDDD.n1403 22.9652
R2425 VDDD.n1573 VDDD.n1572 22.9652
R2426 VDDD.n1545 VDDD.n1417 22.9652
R2427 VDDD.n1540 VDDD.n1539 22.9652
R2428 VDDD.n1512 VDDD.n1431 22.9652
R2429 VDDD.n1507 VDDD.n1506 22.9652
R2430 VDDD.n1479 VDDD.n1445 22.9652
R2431 VDDD.n1829 VDDD.n1828 22.9652
R2432 VDDD.n1801 VDDD.n1319 22.9652
R2433 VDDD.n1796 VDDD.n1795 22.9652
R2434 VDDD.n1768 VDDD.n1333 22.9652
R2435 VDDD.n1763 VDDD.n1762 22.9652
R2436 VDDD.n1735 VDDD.n1347 22.9652
R2437 VDDD.n1730 VDDD.n1729 22.9652
R2438 VDDD.n1702 VDDD.n1361 22.9652
R2439 VDDD.n1697 VDDD.n1696 22.9652
R2440 VDDD.n1669 VDDD.n1375 22.9652
R2441 VDDD.n1875 VDDD.n1874 22.2123
R2442 VDDD.n1880 VDDD.n1879 22.2123
R2443 VDDD.t462 VDDD.t38 21.8203
R2444 VDDD.t119 VDDD.t485 21.8203
R2445 VDDD.t759 VDDD.t956 21.8203
R2446 VDDD.t1056 VDDD.t867 21.8203
R2447 VDDD.t424 VDDD.t872 21.8203
R2448 VDDD.t891 VDDD.t1374 21.8203
R2449 VDDD.t938 VDDD.t46 21.8203
R2450 VDDD.t215 VDDD.t629 21.8203
R2451 VDDD.t72 VDDD.t993 21.8203
R2452 VDDD.t1126 VDDD.t1179 21.8203
R2453 VDDD.n295 VDDD.n293 21.4593
R2454 VDDD.n323 VDDD.n249 21.4593
R2455 VDDD.n328 VDDD.n248 21.4593
R2456 VDDD.n358 VDDD.n357 21.4593
R2457 VDDD.n364 VDDD.n362 21.4593
R2458 VDDD.n392 VDDD.n224 21.4593
R2459 VDDD.n397 VDDD.n223 21.4593
R2460 VDDD.n427 VDDD.n426 21.4593
R2461 VDDD.n433 VDDD.n431 21.4593
R2462 VDDD.n461 VDDD.n199 21.4593
R2463 VDDD.n466 VDDD.n198 21.4593
R2464 VDDD.n496 VDDD.n495 21.4593
R2465 VDDD.n502 VDDD.n500 21.4593
R2466 VDDD.n530 VDDD.n174 21.4593
R2467 VDDD.n535 VDDD.n173 21.4593
R2468 VDDD.n565 VDDD.n564 21.4593
R2469 VDDD.n571 VDDD.n569 21.4593
R2470 VDDD.n599 VDDD.n149 21.4593
R2471 VDDD.n604 VDDD.n148 21.4593
R2472 VDDD.n634 VDDD.n633 21.4593
R2473 VDDD.n641 VDDD.n134 21.4593
R2474 VDDD.n671 VDDD.n670 21.4593
R2475 VDDD.n676 VDDD.n675 21.4593
R2476 VDDD.n705 VDDD.n111 21.4593
R2477 VDDD.n710 VDDD.n109 21.4593
R2478 VDDD.n740 VDDD.n739 21.4593
R2479 VDDD.n745 VDDD.n744 21.4593
R2480 VDDD.n774 VDDD.n86 21.4593
R2481 VDDD.n779 VDDD.n84 21.4593
R2482 VDDD.n809 VDDD.n808 21.4593
R2483 VDDD.n814 VDDD.n813 21.4593
R2484 VDDD.n843 VDDD.n61 21.4593
R2485 VDDD.n848 VDDD.n59 21.4593
R2486 VDDD.n878 VDDD.n877 21.4593
R2487 VDDD.n883 VDDD.n882 21.4593
R2488 VDDD.n912 VDDD.n36 21.4593
R2489 VDDD.n917 VDDD.n34 21.4593
R2490 VDDD.n947 VDDD.n946 21.4593
R2491 VDDD.n952 VDDD.n951 21.4593
R2492 VDDD.n981 VDDD.n11 21.4593
R2493 VDDD.n2444 VDDD.n2443 21.4593
R2494 VDDD.n2439 VDDD.n2438 21.4593
R2495 VDDD.n2411 VDDD.n2410 21.4593
R2496 VDDD.n2406 VDDD.n2405 21.4593
R2497 VDDD.n2378 VDDD.n2377 21.4593
R2498 VDDD.n2373 VDDD.n2372 21.4593
R2499 VDDD.n2345 VDDD.n2344 21.4593
R2500 VDDD.n2340 VDDD.n2339 21.4593
R2501 VDDD.n2312 VDDD.n2311 21.4593
R2502 VDDD.n2307 VDDD.n2306 21.4593
R2503 VDDD.n2279 VDDD.n2278 21.4593
R2504 VDDD.n2148 VDDD.n2147 21.4593
R2505 VDDD.n2143 VDDD.n2142 21.4593
R2506 VDDD.n2115 VDDD.n2114 21.4593
R2507 VDDD.n2110 VDDD.n2109 21.4593
R2508 VDDD.n2082 VDDD.n2081 21.4593
R2509 VDDD.n2077 VDDD.n2076 21.4593
R2510 VDDD.n2049 VDDD.n2048 21.4593
R2511 VDDD.n2044 VDDD.n2043 21.4593
R2512 VDDD.n2016 VDDD.n2015 21.4593
R2513 VDDD.n2011 VDDD.n2010 21.4593
R2514 VDDD.n1983 VDDD.n1982 21.4593
R2515 VDDD.n1612 VDDD.n1611 21.4593
R2516 VDDD.n1607 VDDD.n1606 21.4593
R2517 VDDD.n1579 VDDD.n1578 21.4593
R2518 VDDD.n1574 VDDD.n1573 21.4593
R2519 VDDD.n1546 VDDD.n1545 21.4593
R2520 VDDD.n1541 VDDD.n1540 21.4593
R2521 VDDD.n1513 VDDD.n1512 21.4593
R2522 VDDD.n1508 VDDD.n1507 21.4593
R2523 VDDD.n1480 VDDD.n1479 21.4593
R2524 VDDD.n1802 VDDD.n1801 21.4593
R2525 VDDD.n1797 VDDD.n1796 21.4593
R2526 VDDD.n1769 VDDD.n1768 21.4593
R2527 VDDD.n1764 VDDD.n1763 21.4593
R2528 VDDD.n1736 VDDD.n1735 21.4593
R2529 VDDD.n1731 VDDD.n1730 21.4593
R2530 VDDD.n1703 VDDD.n1702 21.4593
R2531 VDDD.n1698 VDDD.n1697 21.4593
R2532 VDDD.n1670 VDDD.n1669 21.4593
R2533 VDDD.n1881 VDDD.n1880 20.7064
R2534 VDDD.n316 VDDD.n252 20.3299
R2535 VDDD.n352 VDDD.n350 20.3299
R2536 VDDD.n385 VDDD.n227 20.3299
R2537 VDDD.n421 VDDD.n419 20.3299
R2538 VDDD.n454 VDDD.n202 20.3299
R2539 VDDD.n490 VDDD.n488 20.3299
R2540 VDDD.n523 VDDD.n177 20.3299
R2541 VDDD.n559 VDDD.n557 20.3299
R2542 VDDD.n592 VDDD.n152 20.3299
R2543 VDDD.n628 VDDD.n626 20.3299
R2544 VDDD.n648 VDDD.n132 20.3299
R2545 VDDD.n683 VDDD.n682 20.3299
R2546 VDDD.n717 VDDD.n107 20.3299
R2547 VDDD.n752 VDDD.n751 20.3299
R2548 VDDD.n786 VDDD.n82 20.3299
R2549 VDDD.n821 VDDD.n820 20.3299
R2550 VDDD.n855 VDDD.n57 20.3299
R2551 VDDD.n890 VDDD.n889 20.3299
R2552 VDDD.n924 VDDD.n32 20.3299
R2553 VDDD.n959 VDDD.n958 20.3299
R2554 VDDD.n2450 VDDD.n2449 20.3299
R2555 VDDD.n2418 VDDD.n2201 20.3299
R2556 VDDD.n2385 VDDD.n2215 20.3299
R2557 VDDD.n2352 VDDD.n2229 20.3299
R2558 VDDD.n2319 VDDD.n2243 20.3299
R2559 VDDD.n2286 VDDD.n2257 20.3299
R2560 VDDD.n2154 VDDD.n2153 20.3299
R2561 VDDD.n2122 VDDD.n1909 20.3299
R2562 VDDD.n2089 VDDD.n1923 20.3299
R2563 VDDD.n2056 VDDD.n1937 20.3299
R2564 VDDD.n2023 VDDD.n1951 20.3299
R2565 VDDD.n1990 VDDD.n1965 20.3299
R2566 VDDD.n1619 VDDD.n1386 20.3299
R2567 VDDD.n1586 VDDD.n1400 20.3299
R2568 VDDD.n1553 VDDD.n1414 20.3299
R2569 VDDD.n1520 VDDD.n1428 20.3299
R2570 VDDD.n1487 VDDD.n1442 20.3299
R2571 VDDD.n1808 VDDD.n1807 20.3299
R2572 VDDD.n1776 VDDD.n1330 20.3299
R2573 VDDD.n1743 VDDD.n1344 20.3299
R2574 VDDD.n1710 VDDD.n1358 20.3299
R2575 VDDD.n1677 VDDD.n1372 20.3299
R2576 VDDD.n1127 VDDD.n1086 20.3299
R2577 VDDD.n1139 VDDD.n1077 20.3299
R2578 VDDD.n1152 VDDD.n1151 20.3299
R2579 VDDD.n1164 VDDD.n1069 20.3299
R2580 VDDD.n1176 VDDD.n1060 20.3299
R2581 VDDD.n1189 VDDD.n1188 20.3299
R2582 VDDD.n1201 VDDD.n1052 20.3299
R2583 VDDD.n1213 VDDD.n1043 20.3299
R2584 VDDD.n1226 VDDD.n1225 20.3299
R2585 VDDD.n1238 VDDD.n1035 20.3299
R2586 VDDD.n1250 VDDD.n1026 20.3299
R2587 VDDD.n1263 VDDD.n1262 20.3299
R2588 VDDD.n1275 VDDD.n1018 20.3299
R2589 VDDD.n1293 VDDD.n1291 20.3299
R2590 VDDD.n1304 VDDD 19.8156
R2591 VDDD.n2481 VDDD 18.9706
R2592 VDDD.n1858 VDDD.n1854 18.824
R2593 VDDD.t569 VDDD.t1324 18.4634
R2594 VDDD.t372 VDDD.t40 18.4634
R2595 VDDD.t1333 VDDD.t1320 18.4634
R2596 VDDD.t1408 VDDD.t585 18.4634
R2597 VDDD.t428 VDDD.t1058 18.4634
R2598 VDDD.t893 VDDD.t762 18.4634
R2599 VDDD.t1015 VDDD.t199 18.4634
R2600 VDDD.t296 VDDD.t164 18.4634
R2601 VDDD.t877 VDDD.t203 18.4634
R2602 VDDD.t1344 VDDD.t1376 18.4634
R2603 VDDD.n289 VDDD.n260 18.4476
R2604 VDDD.n982 VDDD.n9 18.4476
R2605 VDDD.n2273 VDDD.n2272 18.2003
R2606 VDDD.n300 VDDD.n258 18.0711
R2607 VDDD.n334 VDDD.n333 18.0711
R2608 VDDD.n369 VDDD.n233 18.0711
R2609 VDDD.n403 VDDD.n402 18.0711
R2610 VDDD.n438 VDDD.n208 18.0711
R2611 VDDD.n472 VDDD.n471 18.0711
R2612 VDDD.n507 VDDD.n183 18.0711
R2613 VDDD.n541 VDDD.n540 18.0711
R2614 VDDD.n576 VDDD.n158 18.0711
R2615 VDDD.n610 VDDD.n609 18.0711
R2616 VDDD.n664 VDDD.n125 18.0711
R2617 VDDD.n700 VDDD.n699 18.0711
R2618 VDDD.n733 VDDD.n100 18.0711
R2619 VDDD.n769 VDDD.n768 18.0711
R2620 VDDD.n802 VDDD.n75 18.0711
R2621 VDDD.n838 VDDD.n837 18.0711
R2622 VDDD.n871 VDDD.n50 18.0711
R2623 VDDD.n907 VDDD.n906 18.0711
R2624 VDDD.n940 VDDD.n25 18.0711
R2625 VDDD.n976 VDDD.n975 18.0711
R2626 VDDD.n2469 VDDD.n2180 18.0711
R2627 VDDD.n2433 VDDD.n2193 18.0711
R2628 VDDD.n2400 VDDD.n2207 18.0711
R2629 VDDD.n2367 VDDD.n2221 18.0711
R2630 VDDD.n2334 VDDD.n2235 18.0711
R2631 VDDD.n2301 VDDD.n2249 18.0711
R2632 VDDD.n2173 VDDD.n1888 18.0711
R2633 VDDD.n2137 VDDD.n1901 18.0711
R2634 VDDD.n2104 VDDD.n1915 18.0711
R2635 VDDD.n2071 VDDD.n1929 18.0711
R2636 VDDD.n2038 VDDD.n1943 18.0711
R2637 VDDD.n2005 VDDD.n1957 18.0711
R2638 VDDD.n1634 VDDD.n1378 18.0711
R2639 VDDD.n1601 VDDD.n1392 18.0711
R2640 VDDD.n1568 VDDD.n1406 18.0711
R2641 VDDD.n1535 VDDD.n1420 18.0711
R2642 VDDD.n1502 VDDD.n1434 18.0711
R2643 VDDD.n1827 VDDD.n1309 18.0711
R2644 VDDD.n1791 VDDD.n1322 18.0711
R2645 VDDD.n1758 VDDD.n1336 18.0711
R2646 VDDD.n1725 VDDD.n1350 18.0711
R2647 VDDD.n1692 VDDD.n1364 18.0711
R2648 VDDD.n2474 VDDD 17.7752
R2649 VDDD.n1122 VDDD.n1121 14.3064
R2650 VDDD.n1145 VDDD.n1144 14.3064
R2651 VDDD.n1159 VDDD.n1158 14.3064
R2652 VDDD.n1182 VDDD.n1181 14.3064
R2653 VDDD.n1196 VDDD.n1195 14.3064
R2654 VDDD.n1219 VDDD.n1218 14.3064
R2655 VDDD.n1233 VDDD.n1232 14.3064
R2656 VDDD.n1256 VDDD.n1255 14.3064
R2657 VDDD.n1270 VDDD.n1269 14.3064
R2658 VDDD.n1295 VDDD.n1294 14.3064
R2659 VDDD.n1870 VDDD.n1848 13.5534
R2660 VDDD.n1105 VDDD.n1104 13.4417
R2661 VDDD.t1390 VDDD.t576 13.4281
R2662 VDDD.t167 VDDD.t578 13.4281
R2663 VDDD.t520 VDDD.t883 13.4281
R2664 VDDD.t522 VDDD.t1152 13.4281
R2665 VDDD.t223 VDDD.t652 13.4281
R2666 VDDD.t765 VDDD.t654 13.4281
R2667 VDDD.t1140 VDDD.t757 13.4281
R2668 VDDD.t1138 VDDD.t1438 13.4281
R2669 VDDD.t1434 VDDD.t1241 13.4281
R2670 VDDD.t445 VDDD.t1243 13.4281
R2671 VDDD.t139 VDDD.t425 13.4281
R2672 VDDD.t137 VDDD.t1436 13.4281
R2673 VDDD.t1340 VDDD.t802 13.4281
R2674 VDDD.t1148 VDDD.t412 13.4281
R2675 VDDD.t719 VDDD.t939 13.4281
R2676 VDDD.t280 VDDD.t66 13.4281
R2677 VDDD.t1392 VDDD.t348 13.4281
R2678 VDDD.t1177 VDDD.t346 13.4281
R2679 VDDD.t814 VDDD.t70 13.4281
R2680 VDDD.t810 VDDD.t68 13.4281
R2681 VDDD.n1121 VDDD.n1120 13.177
R2682 VDDD.n1146 VDDD.n1145 13.177
R2683 VDDD.n1158 VDDD.n1157 13.177
R2684 VDDD.n1183 VDDD.n1182 13.177
R2685 VDDD.n1195 VDDD.n1194 13.177
R2686 VDDD.n1220 VDDD.n1219 13.177
R2687 VDDD.n1232 VDDD.n1231 13.177
R2688 VDDD.n1257 VDDD.n1256 13.177
R2689 VDDD.n1269 VDDD.n1268 13.177
R2690 VDDD.n1294 VDDD.n1011 13.177
R2691 VDDD.n288 VDDD.n287 12.424
R2692 VDDD.n988 VDDD.n986 12.424
R2693 VDDD.n1461 VDDD.n1460 12.424
R2694 VDDD.n2492 VDDD.n2491 11
R2695 VDDD.n2475 VDDD.n1305 10.7339
R2696 VDDD.n2476 VDDD.n2475 10.2118
R2697 VDDD.n1302 VDDD.n1301 9.78874
R2698 VDDD.n1115 VDDD.n1089 9.78874
R2699 VDDD.n1119 VDDD.n1089 9.78874
R2700 VDDD.n1147 VDDD.n1074 9.78874
R2701 VDDD.n1151 VDDD.n1074 9.78874
R2702 VDDD.n1152 VDDD.n1072 9.78874
R2703 VDDD.n1156 VDDD.n1072 9.78874
R2704 VDDD.n1184 VDDD.n1057 9.78874
R2705 VDDD.n1188 VDDD.n1057 9.78874
R2706 VDDD.n1189 VDDD.n1055 9.78874
R2707 VDDD.n1193 VDDD.n1055 9.78874
R2708 VDDD.n1221 VDDD.n1040 9.78874
R2709 VDDD.n1225 VDDD.n1040 9.78874
R2710 VDDD.n1226 VDDD.n1038 9.78874
R2711 VDDD.n1230 VDDD.n1038 9.78874
R2712 VDDD.n1258 VDDD.n1023 9.78874
R2713 VDDD.n1262 VDDD.n1023 9.78874
R2714 VDDD.n1263 VDDD.n1021 9.78874
R2715 VDDD.n1267 VDDD.n1021 9.78874
R2716 VDDD.n1301 VDDD.n1300 9.78874
R2717 VDDD.n2272 VDDD.n2271 9.65395
R2718 VDDD.n1980 VDDD.n1979 9.54619
R2719 VDDD.n1103 VDDD.n1092 9.45675
R2720 VDDD.n280 VDDD.n278 9.41227
R2721 VDDD.n310 VDDD.n254 9.41227
R2722 VDDD.n345 VDDD.n344 9.41227
R2723 VDDD.n379 VDDD.n229 9.41227
R2724 VDDD.n414 VDDD.n413 9.41227
R2725 VDDD.n448 VDDD.n204 9.41227
R2726 VDDD.n483 VDDD.n482 9.41227
R2727 VDDD.n517 VDDD.n179 9.41227
R2728 VDDD.n552 VDDD.n551 9.41227
R2729 VDDD.n586 VDDD.n154 9.41227
R2730 VDDD.n621 VDDD.n620 9.41227
R2731 VDDD.n654 VDDD.n129 9.41227
R2732 VDDD.n689 VDDD.n688 9.41227
R2733 VDDD.n723 VDDD.n104 9.41227
R2734 VDDD.n758 VDDD.n757 9.41227
R2735 VDDD.n792 VDDD.n79 9.41227
R2736 VDDD.n827 VDDD.n826 9.41227
R2737 VDDD.n861 VDDD.n54 9.41227
R2738 VDDD.n896 VDDD.n895 9.41227
R2739 VDDD.n930 VDDD.n29 9.41227
R2740 VDDD.n965 VDDD.n964 9.41227
R2741 VDDD.n998 VDDD.n997 9.41227
R2742 VDDD.n2456 VDDD.n2455 9.41227
R2743 VDDD.n2424 VDDD.n2198 9.41227
R2744 VDDD.n2391 VDDD.n2212 9.41227
R2745 VDDD.n2358 VDDD.n2226 9.41227
R2746 VDDD.n2325 VDDD.n2240 9.41227
R2747 VDDD.n2292 VDDD.n2254 9.41227
R2748 VDDD.n2160 VDDD.n2159 9.41227
R2749 VDDD.n2128 VDDD.n1906 9.41227
R2750 VDDD.n2095 VDDD.n1920 9.41227
R2751 VDDD.n2062 VDDD.n1934 9.41227
R2752 VDDD.n2029 VDDD.n1948 9.41227
R2753 VDDD.n1996 VDDD.n1962 9.41227
R2754 VDDD.n1625 VDDD.n1383 9.41227
R2755 VDDD.n1592 VDDD.n1397 9.41227
R2756 VDDD.n1559 VDDD.n1411 9.41227
R2757 VDDD.n1526 VDDD.n1425 9.41227
R2758 VDDD.n1493 VDDD.n1439 9.41227
R2759 VDDD.n1468 VDDD.n1467 9.41227
R2760 VDDD.n1814 VDDD.n1813 9.41227
R2761 VDDD.n1782 VDDD.n1327 9.41227
R2762 VDDD.n1749 VDDD.n1341 9.41227
R2763 VDDD.n1716 VDDD.n1355 9.41227
R2764 VDDD.n1683 VDDD.n1369 9.41227
R2765 VDDD.n1106 VDDD.n1105 9.41227
R2766 VDDD.n1133 VDDD.n1132 9.41227
R2767 VDDD.n1134 VDDD.n1133 9.41227
R2768 VDDD.n1170 VDDD.n1169 9.41227
R2769 VDDD.n1171 VDDD.n1170 9.41227
R2770 VDDD.n1207 VDDD.n1206 9.41227
R2771 VDDD.n1208 VDDD.n1207 9.41227
R2772 VDDD.n1244 VDDD.n1243 9.41227
R2773 VDDD.n1245 VDDD.n1244 9.41227
R2774 VDDD.n1283 VDDD.n1015 9.41227
R2775 VDDD.n1284 VDDD.n1283 9.41227
R2776 VDDD.n1885 VDDD.n1841 9.32421
R2777 VDDD.n1856 VDDD.n1854 9.3005
R2778 VDDD.n1858 VDDD.n1857 9.3005
R2779 VDDD.n1859 VDDD.n1852 9.3005
R2780 VDDD.n1864 VDDD.n1863 9.3005
R2781 VDDD.n1865 VDDD.n1851 9.3005
R2782 VDDD.n1867 VDDD.n1866 9.3005
R2783 VDDD.n1869 VDDD.n1849 9.3005
R2784 VDDD.n1871 VDDD.n1870 9.3005
R2785 VDDD.n1873 VDDD.n1872 9.3005
R2786 VDDD.n1874 VDDD.n1847 9.3005
R2787 VDDD.n1876 VDDD.n1875 9.3005
R2788 VDDD.n1877 VDDD.n1846 9.3005
R2789 VDDD.n1879 VDDD.n1878 9.3005
R2790 VDDD.n1880 VDDD.n1844 9.3005
R2791 VDDD.n1881 VDDD.n1843 9.3005
R2792 VDDD.n1882 VDDD.n1842 9.3005
R2793 VDDD.n1884 VDDD.n1883 9.3005
R2794 VDDD.n1980 VDDD.n1968 9.3005
R2795 VDDD.n1982 VDDD.n1981 9.3005
R2796 VDDD.n1983 VDDD.n1967 9.3005
R2797 VDDD.n1984 VDDD.n1966 9.3005
R2798 VDDD.n1987 VDDD.n1986 9.3005
R2799 VDDD.n1988 VDDD.n1965 9.3005
R2800 VDDD.n1990 VDDD.n1989 9.3005
R2801 VDDD.n1991 VDDD.n1963 9.3005
R2802 VDDD.n1993 VDDD.n1992 9.3005
R2803 VDDD.n1994 VDDD.n1962 9.3005
R2804 VDDD.n1996 VDDD.n1995 9.3005
R2805 VDDD.n1997 VDDD.n1960 9.3005
R2806 VDDD.n2000 VDDD.n1999 9.3005
R2807 VDDD.n2001 VDDD.n1959 9.3005
R2808 VDDD.n2003 VDDD.n2002 9.3005
R2809 VDDD.n2004 VDDD.n1958 9.3005
R2810 VDDD.n2006 VDDD.n2005 9.3005
R2811 VDDD.n2007 VDDD.n1957 9.3005
R2812 VDDD.n2009 VDDD.n2008 9.3005
R2813 VDDD.n2010 VDDD.n1955 9.3005
R2814 VDDD.n2012 VDDD.n2011 9.3005
R2815 VDDD.n2013 VDDD.n1954 9.3005
R2816 VDDD.n2015 VDDD.n2014 9.3005
R2817 VDDD.n2016 VDDD.n1953 9.3005
R2818 VDDD.n2017 VDDD.n1952 9.3005
R2819 VDDD.n2020 VDDD.n2019 9.3005
R2820 VDDD.n2021 VDDD.n1951 9.3005
R2821 VDDD.n2023 VDDD.n2022 9.3005
R2822 VDDD.n2024 VDDD.n1949 9.3005
R2823 VDDD.n2026 VDDD.n2025 9.3005
R2824 VDDD.n2027 VDDD.n1948 9.3005
R2825 VDDD.n2029 VDDD.n2028 9.3005
R2826 VDDD.n2030 VDDD.n1946 9.3005
R2827 VDDD.n2033 VDDD.n2032 9.3005
R2828 VDDD.n2034 VDDD.n1945 9.3005
R2829 VDDD.n2036 VDDD.n2035 9.3005
R2830 VDDD.n2037 VDDD.n1944 9.3005
R2831 VDDD.n2039 VDDD.n2038 9.3005
R2832 VDDD.n2040 VDDD.n1943 9.3005
R2833 VDDD.n2042 VDDD.n2041 9.3005
R2834 VDDD.n2043 VDDD.n1941 9.3005
R2835 VDDD.n2045 VDDD.n2044 9.3005
R2836 VDDD.n2046 VDDD.n1940 9.3005
R2837 VDDD.n2048 VDDD.n2047 9.3005
R2838 VDDD.n2049 VDDD.n1939 9.3005
R2839 VDDD.n2050 VDDD.n1938 9.3005
R2840 VDDD.n2053 VDDD.n2052 9.3005
R2841 VDDD.n2054 VDDD.n1937 9.3005
R2842 VDDD.n2056 VDDD.n2055 9.3005
R2843 VDDD.n2057 VDDD.n1935 9.3005
R2844 VDDD.n2059 VDDD.n2058 9.3005
R2845 VDDD.n2060 VDDD.n1934 9.3005
R2846 VDDD.n2062 VDDD.n2061 9.3005
R2847 VDDD.n2063 VDDD.n1932 9.3005
R2848 VDDD.n2066 VDDD.n2065 9.3005
R2849 VDDD.n2067 VDDD.n1931 9.3005
R2850 VDDD.n2069 VDDD.n2068 9.3005
R2851 VDDD.n2070 VDDD.n1930 9.3005
R2852 VDDD.n2072 VDDD.n2071 9.3005
R2853 VDDD.n2073 VDDD.n1929 9.3005
R2854 VDDD.n2075 VDDD.n2074 9.3005
R2855 VDDD.n2076 VDDD.n1927 9.3005
R2856 VDDD.n2078 VDDD.n2077 9.3005
R2857 VDDD.n2079 VDDD.n1926 9.3005
R2858 VDDD.n2081 VDDD.n2080 9.3005
R2859 VDDD.n2082 VDDD.n1925 9.3005
R2860 VDDD.n2083 VDDD.n1924 9.3005
R2861 VDDD.n2086 VDDD.n2085 9.3005
R2862 VDDD.n2087 VDDD.n1923 9.3005
R2863 VDDD.n2089 VDDD.n2088 9.3005
R2864 VDDD.n2090 VDDD.n1921 9.3005
R2865 VDDD.n2092 VDDD.n2091 9.3005
R2866 VDDD.n2093 VDDD.n1920 9.3005
R2867 VDDD.n2095 VDDD.n2094 9.3005
R2868 VDDD.n2096 VDDD.n1918 9.3005
R2869 VDDD.n2099 VDDD.n2098 9.3005
R2870 VDDD.n2100 VDDD.n1917 9.3005
R2871 VDDD.n2102 VDDD.n2101 9.3005
R2872 VDDD.n2103 VDDD.n1916 9.3005
R2873 VDDD.n2105 VDDD.n2104 9.3005
R2874 VDDD.n2106 VDDD.n1915 9.3005
R2875 VDDD.n2108 VDDD.n2107 9.3005
R2876 VDDD.n2109 VDDD.n1913 9.3005
R2877 VDDD.n2111 VDDD.n2110 9.3005
R2878 VDDD.n2112 VDDD.n1912 9.3005
R2879 VDDD.n2114 VDDD.n2113 9.3005
R2880 VDDD.n2115 VDDD.n1911 9.3005
R2881 VDDD.n2116 VDDD.n1910 9.3005
R2882 VDDD.n2119 VDDD.n2118 9.3005
R2883 VDDD.n2120 VDDD.n1909 9.3005
R2884 VDDD.n2122 VDDD.n2121 9.3005
R2885 VDDD.n2123 VDDD.n1907 9.3005
R2886 VDDD.n2125 VDDD.n2124 9.3005
R2887 VDDD.n2126 VDDD.n1906 9.3005
R2888 VDDD.n2128 VDDD.n2127 9.3005
R2889 VDDD.n2129 VDDD.n1904 9.3005
R2890 VDDD.n2132 VDDD.n2131 9.3005
R2891 VDDD.n2133 VDDD.n1903 9.3005
R2892 VDDD.n2135 VDDD.n2134 9.3005
R2893 VDDD.n2136 VDDD.n1902 9.3005
R2894 VDDD.n2138 VDDD.n2137 9.3005
R2895 VDDD.n2139 VDDD.n1901 9.3005
R2896 VDDD.n2141 VDDD.n2140 9.3005
R2897 VDDD.n2142 VDDD.n1899 9.3005
R2898 VDDD.n2144 VDDD.n2143 9.3005
R2899 VDDD.n2145 VDDD.n1898 9.3005
R2900 VDDD.n2147 VDDD.n2146 9.3005
R2901 VDDD.n2148 VDDD.n1897 9.3005
R2902 VDDD.n2150 VDDD.n2149 9.3005
R2903 VDDD.n2152 VDDD.n2151 9.3005
R2904 VDDD.n2153 VDDD.n1894 9.3005
R2905 VDDD.n2155 VDDD.n2154 9.3005
R2906 VDDD.n2156 VDDD.n1893 9.3005
R2907 VDDD.n2158 VDDD.n2157 9.3005
R2908 VDDD.n2159 VDDD.n1892 9.3005
R2909 VDDD.n2160 VDDD.n1891 9.3005
R2910 VDDD.n2164 VDDD.n2163 9.3005
R2911 VDDD.n2165 VDDD.n1890 9.3005
R2912 VDDD.n2167 VDDD.n2166 9.3005
R2913 VDDD.n2168 VDDD.n1889 9.3005
R2914 VDDD.n2170 VDDD.n2169 9.3005
R2915 VDDD.n2171 VDDD.n1888 9.3005
R2916 VDDD.n2173 VDDD.n2172 9.3005
R2917 VDDD.n2174 VDDD.n1886 9.3005
R2918 VDDD.n2275 VDDD.n2274 9.3005
R2919 VDDD.n2276 VDDD.n2260 9.3005
R2920 VDDD.n2278 VDDD.n2277 9.3005
R2921 VDDD.n2279 VDDD.n2259 9.3005
R2922 VDDD.n2280 VDDD.n2258 9.3005
R2923 VDDD.n2283 VDDD.n2282 9.3005
R2924 VDDD.n2284 VDDD.n2257 9.3005
R2925 VDDD.n2286 VDDD.n2285 9.3005
R2926 VDDD.n2287 VDDD.n2255 9.3005
R2927 VDDD.n2289 VDDD.n2288 9.3005
R2928 VDDD.n2290 VDDD.n2254 9.3005
R2929 VDDD.n2292 VDDD.n2291 9.3005
R2930 VDDD.n2293 VDDD.n2252 9.3005
R2931 VDDD.n2296 VDDD.n2295 9.3005
R2932 VDDD.n2297 VDDD.n2251 9.3005
R2933 VDDD.n2299 VDDD.n2298 9.3005
R2934 VDDD.n2300 VDDD.n2250 9.3005
R2935 VDDD.n2302 VDDD.n2301 9.3005
R2936 VDDD.n2303 VDDD.n2249 9.3005
R2937 VDDD.n2305 VDDD.n2304 9.3005
R2938 VDDD.n2306 VDDD.n2247 9.3005
R2939 VDDD.n2308 VDDD.n2307 9.3005
R2940 VDDD.n2309 VDDD.n2246 9.3005
R2941 VDDD.n2311 VDDD.n2310 9.3005
R2942 VDDD.n2312 VDDD.n2245 9.3005
R2943 VDDD.n2313 VDDD.n2244 9.3005
R2944 VDDD.n2316 VDDD.n2315 9.3005
R2945 VDDD.n2317 VDDD.n2243 9.3005
R2946 VDDD.n2319 VDDD.n2318 9.3005
R2947 VDDD.n2320 VDDD.n2241 9.3005
R2948 VDDD.n2322 VDDD.n2321 9.3005
R2949 VDDD.n2323 VDDD.n2240 9.3005
R2950 VDDD.n2325 VDDD.n2324 9.3005
R2951 VDDD.n2326 VDDD.n2238 9.3005
R2952 VDDD.n2329 VDDD.n2328 9.3005
R2953 VDDD.n2330 VDDD.n2237 9.3005
R2954 VDDD.n2332 VDDD.n2331 9.3005
R2955 VDDD.n2333 VDDD.n2236 9.3005
R2956 VDDD.n2335 VDDD.n2334 9.3005
R2957 VDDD.n2336 VDDD.n2235 9.3005
R2958 VDDD.n2338 VDDD.n2337 9.3005
R2959 VDDD.n2339 VDDD.n2233 9.3005
R2960 VDDD.n2341 VDDD.n2340 9.3005
R2961 VDDD.n2342 VDDD.n2232 9.3005
R2962 VDDD.n2344 VDDD.n2343 9.3005
R2963 VDDD.n2345 VDDD.n2231 9.3005
R2964 VDDD.n2346 VDDD.n2230 9.3005
R2965 VDDD.n2349 VDDD.n2348 9.3005
R2966 VDDD.n2350 VDDD.n2229 9.3005
R2967 VDDD.n2352 VDDD.n2351 9.3005
R2968 VDDD.n2353 VDDD.n2227 9.3005
R2969 VDDD.n2355 VDDD.n2354 9.3005
R2970 VDDD.n2356 VDDD.n2226 9.3005
R2971 VDDD.n2358 VDDD.n2357 9.3005
R2972 VDDD.n2359 VDDD.n2224 9.3005
R2973 VDDD.n2362 VDDD.n2361 9.3005
R2974 VDDD.n2363 VDDD.n2223 9.3005
R2975 VDDD.n2365 VDDD.n2364 9.3005
R2976 VDDD.n2366 VDDD.n2222 9.3005
R2977 VDDD.n2368 VDDD.n2367 9.3005
R2978 VDDD.n2369 VDDD.n2221 9.3005
R2979 VDDD.n2371 VDDD.n2370 9.3005
R2980 VDDD.n2372 VDDD.n2219 9.3005
R2981 VDDD.n2374 VDDD.n2373 9.3005
R2982 VDDD.n2375 VDDD.n2218 9.3005
R2983 VDDD.n2377 VDDD.n2376 9.3005
R2984 VDDD.n2378 VDDD.n2217 9.3005
R2985 VDDD.n2379 VDDD.n2216 9.3005
R2986 VDDD.n2382 VDDD.n2381 9.3005
R2987 VDDD.n2383 VDDD.n2215 9.3005
R2988 VDDD.n2385 VDDD.n2384 9.3005
R2989 VDDD.n2386 VDDD.n2213 9.3005
R2990 VDDD.n2388 VDDD.n2387 9.3005
R2991 VDDD.n2389 VDDD.n2212 9.3005
R2992 VDDD.n2391 VDDD.n2390 9.3005
R2993 VDDD.n2392 VDDD.n2210 9.3005
R2994 VDDD.n2395 VDDD.n2394 9.3005
R2995 VDDD.n2396 VDDD.n2209 9.3005
R2996 VDDD.n2398 VDDD.n2397 9.3005
R2997 VDDD.n2399 VDDD.n2208 9.3005
R2998 VDDD.n2401 VDDD.n2400 9.3005
R2999 VDDD.n2402 VDDD.n2207 9.3005
R3000 VDDD.n2404 VDDD.n2403 9.3005
R3001 VDDD.n2405 VDDD.n2205 9.3005
R3002 VDDD.n2407 VDDD.n2406 9.3005
R3003 VDDD.n2408 VDDD.n2204 9.3005
R3004 VDDD.n2410 VDDD.n2409 9.3005
R3005 VDDD.n2411 VDDD.n2203 9.3005
R3006 VDDD.n2412 VDDD.n2202 9.3005
R3007 VDDD.n2415 VDDD.n2414 9.3005
R3008 VDDD.n2416 VDDD.n2201 9.3005
R3009 VDDD.n2418 VDDD.n2417 9.3005
R3010 VDDD.n2419 VDDD.n2199 9.3005
R3011 VDDD.n2421 VDDD.n2420 9.3005
R3012 VDDD.n2422 VDDD.n2198 9.3005
R3013 VDDD.n2424 VDDD.n2423 9.3005
R3014 VDDD.n2425 VDDD.n2196 9.3005
R3015 VDDD.n2428 VDDD.n2427 9.3005
R3016 VDDD.n2429 VDDD.n2195 9.3005
R3017 VDDD.n2431 VDDD.n2430 9.3005
R3018 VDDD.n2432 VDDD.n2194 9.3005
R3019 VDDD.n2434 VDDD.n2433 9.3005
R3020 VDDD.n2435 VDDD.n2193 9.3005
R3021 VDDD.n2437 VDDD.n2436 9.3005
R3022 VDDD.n2438 VDDD.n2191 9.3005
R3023 VDDD.n2440 VDDD.n2439 9.3005
R3024 VDDD.n2441 VDDD.n2190 9.3005
R3025 VDDD.n2443 VDDD.n2442 9.3005
R3026 VDDD.n2444 VDDD.n2189 9.3005
R3027 VDDD.n2446 VDDD.n2445 9.3005
R3028 VDDD.n2448 VDDD.n2447 9.3005
R3029 VDDD.n2449 VDDD.n2186 9.3005
R3030 VDDD.n2451 VDDD.n2450 9.3005
R3031 VDDD.n2452 VDDD.n2185 9.3005
R3032 VDDD.n2454 VDDD.n2453 9.3005
R3033 VDDD.n2455 VDDD.n2184 9.3005
R3034 VDDD.n2456 VDDD.n2183 9.3005
R3035 VDDD.n2460 VDDD.n2459 9.3005
R3036 VDDD.n2461 VDDD.n2182 9.3005
R3037 VDDD.n2463 VDDD.n2462 9.3005
R3038 VDDD.n2464 VDDD.n2181 9.3005
R3039 VDDD.n2466 VDDD.n2465 9.3005
R3040 VDDD.n2467 VDDD.n2180 9.3005
R3041 VDDD.n2469 VDDD.n2468 9.3005
R3042 VDDD.n2470 VDDD.n2178 9.3005
R3043 VDDD.n1667 VDDD.n1375 9.3005
R3044 VDDD.n1669 VDDD.n1668 9.3005
R3045 VDDD.n1670 VDDD.n1374 9.3005
R3046 VDDD.n1671 VDDD.n1373 9.3005
R3047 VDDD.n1674 VDDD.n1673 9.3005
R3048 VDDD.n1675 VDDD.n1372 9.3005
R3049 VDDD.n1677 VDDD.n1676 9.3005
R3050 VDDD.n1678 VDDD.n1370 9.3005
R3051 VDDD.n1680 VDDD.n1679 9.3005
R3052 VDDD.n1681 VDDD.n1369 9.3005
R3053 VDDD.n1683 VDDD.n1682 9.3005
R3054 VDDD.n1684 VDDD.n1367 9.3005
R3055 VDDD.n1687 VDDD.n1686 9.3005
R3056 VDDD.n1688 VDDD.n1366 9.3005
R3057 VDDD.n1690 VDDD.n1689 9.3005
R3058 VDDD.n1691 VDDD.n1365 9.3005
R3059 VDDD.n1693 VDDD.n1692 9.3005
R3060 VDDD.n1694 VDDD.n1364 9.3005
R3061 VDDD.n1696 VDDD.n1695 9.3005
R3062 VDDD.n1697 VDDD.n1362 9.3005
R3063 VDDD.n1699 VDDD.n1698 9.3005
R3064 VDDD.n1700 VDDD.n1361 9.3005
R3065 VDDD.n1702 VDDD.n1701 9.3005
R3066 VDDD.n1703 VDDD.n1360 9.3005
R3067 VDDD.n1704 VDDD.n1359 9.3005
R3068 VDDD.n1707 VDDD.n1706 9.3005
R3069 VDDD.n1708 VDDD.n1358 9.3005
R3070 VDDD.n1710 VDDD.n1709 9.3005
R3071 VDDD.n1711 VDDD.n1356 9.3005
R3072 VDDD.n1713 VDDD.n1712 9.3005
R3073 VDDD.n1714 VDDD.n1355 9.3005
R3074 VDDD.n1716 VDDD.n1715 9.3005
R3075 VDDD.n1717 VDDD.n1353 9.3005
R3076 VDDD.n1720 VDDD.n1719 9.3005
R3077 VDDD.n1721 VDDD.n1352 9.3005
R3078 VDDD.n1723 VDDD.n1722 9.3005
R3079 VDDD.n1724 VDDD.n1351 9.3005
R3080 VDDD.n1726 VDDD.n1725 9.3005
R3081 VDDD.n1727 VDDD.n1350 9.3005
R3082 VDDD.n1729 VDDD.n1728 9.3005
R3083 VDDD.n1730 VDDD.n1348 9.3005
R3084 VDDD.n1732 VDDD.n1731 9.3005
R3085 VDDD.n1733 VDDD.n1347 9.3005
R3086 VDDD.n1735 VDDD.n1734 9.3005
R3087 VDDD.n1736 VDDD.n1346 9.3005
R3088 VDDD.n1737 VDDD.n1345 9.3005
R3089 VDDD.n1740 VDDD.n1739 9.3005
R3090 VDDD.n1741 VDDD.n1344 9.3005
R3091 VDDD.n1743 VDDD.n1742 9.3005
R3092 VDDD.n1744 VDDD.n1342 9.3005
R3093 VDDD.n1746 VDDD.n1745 9.3005
R3094 VDDD.n1747 VDDD.n1341 9.3005
R3095 VDDD.n1749 VDDD.n1748 9.3005
R3096 VDDD.n1750 VDDD.n1339 9.3005
R3097 VDDD.n1753 VDDD.n1752 9.3005
R3098 VDDD.n1754 VDDD.n1338 9.3005
R3099 VDDD.n1756 VDDD.n1755 9.3005
R3100 VDDD.n1757 VDDD.n1337 9.3005
R3101 VDDD.n1759 VDDD.n1758 9.3005
R3102 VDDD.n1760 VDDD.n1336 9.3005
R3103 VDDD.n1762 VDDD.n1761 9.3005
R3104 VDDD.n1763 VDDD.n1334 9.3005
R3105 VDDD.n1765 VDDD.n1764 9.3005
R3106 VDDD.n1766 VDDD.n1333 9.3005
R3107 VDDD.n1768 VDDD.n1767 9.3005
R3108 VDDD.n1769 VDDD.n1332 9.3005
R3109 VDDD.n1770 VDDD.n1331 9.3005
R3110 VDDD.n1773 VDDD.n1772 9.3005
R3111 VDDD.n1774 VDDD.n1330 9.3005
R3112 VDDD.n1776 VDDD.n1775 9.3005
R3113 VDDD.n1777 VDDD.n1328 9.3005
R3114 VDDD.n1779 VDDD.n1778 9.3005
R3115 VDDD.n1780 VDDD.n1327 9.3005
R3116 VDDD.n1782 VDDD.n1781 9.3005
R3117 VDDD.n1783 VDDD.n1325 9.3005
R3118 VDDD.n1786 VDDD.n1785 9.3005
R3119 VDDD.n1787 VDDD.n1324 9.3005
R3120 VDDD.n1789 VDDD.n1788 9.3005
R3121 VDDD.n1790 VDDD.n1323 9.3005
R3122 VDDD.n1792 VDDD.n1791 9.3005
R3123 VDDD.n1793 VDDD.n1322 9.3005
R3124 VDDD.n1795 VDDD.n1794 9.3005
R3125 VDDD.n1796 VDDD.n1320 9.3005
R3126 VDDD.n1798 VDDD.n1797 9.3005
R3127 VDDD.n1799 VDDD.n1319 9.3005
R3128 VDDD.n1801 VDDD.n1800 9.3005
R3129 VDDD.n1802 VDDD.n1318 9.3005
R3130 VDDD.n1804 VDDD.n1803 9.3005
R3131 VDDD.n1806 VDDD.n1805 9.3005
R3132 VDDD.n1807 VDDD.n1315 9.3005
R3133 VDDD.n1809 VDDD.n1808 9.3005
R3134 VDDD.n1810 VDDD.n1314 9.3005
R3135 VDDD.n1812 VDDD.n1811 9.3005
R3136 VDDD.n1813 VDDD.n1313 9.3005
R3137 VDDD.n1814 VDDD.n1312 9.3005
R3138 VDDD.n1818 VDDD.n1817 9.3005
R3139 VDDD.n1819 VDDD.n1311 9.3005
R3140 VDDD.n1821 VDDD.n1820 9.3005
R3141 VDDD.n1822 VDDD.n1310 9.3005
R3142 VDDD.n1824 VDDD.n1823 9.3005
R3143 VDDD.n1825 VDDD.n1309 9.3005
R3144 VDDD.n1827 VDDD.n1826 9.3005
R3145 VDDD.n1828 VDDD.n1307 9.3005
R3146 VDDD.n1657 VDDD.n1654 9.3005
R3147 VDDD.n1666 VDDD.n1665 9.3005
R3148 VDDD.n1644 VDDD.n1641 9.3005
R3149 VDDD.n1653 VDDD.n1652 9.3005
R3150 VDDD.n1639 VDDD.n1377 9.3005
R3151 VDDD.n1638 VDDD.n1637 9.3005
R3152 VDDD.n1636 VDDD.n1378 9.3005
R3153 VDDD.n1635 VDDD.n1634 9.3005
R3154 VDDD.n1633 VDDD.n1379 9.3005
R3155 VDDD.n1632 VDDD.n1631 9.3005
R3156 VDDD.n1630 VDDD.n1380 9.3005
R3157 VDDD.n1629 VDDD.n1628 9.3005
R3158 VDDD.n1626 VDDD.n1381 9.3005
R3159 VDDD.n1625 VDDD.n1624 9.3005
R3160 VDDD.n1623 VDDD.n1383 9.3005
R3161 VDDD.n1622 VDDD.n1621 9.3005
R3162 VDDD.n1620 VDDD.n1384 9.3005
R3163 VDDD.n1619 VDDD.n1618 9.3005
R3164 VDDD.n1617 VDDD.n1386 9.3005
R3165 VDDD.n1616 VDDD.n1615 9.3005
R3166 VDDD.n1613 VDDD.n1387 9.3005
R3167 VDDD.n1612 VDDD.n1388 9.3005
R3168 VDDD.n1611 VDDD.n1610 9.3005
R3169 VDDD.n1609 VDDD.n1389 9.3005
R3170 VDDD.n1608 VDDD.n1607 9.3005
R3171 VDDD.n1606 VDDD.n1391 9.3005
R3172 VDDD.n1605 VDDD.n1604 9.3005
R3173 VDDD.n1603 VDDD.n1392 9.3005
R3174 VDDD.n1602 VDDD.n1601 9.3005
R3175 VDDD.n1600 VDDD.n1393 9.3005
R3176 VDDD.n1599 VDDD.n1598 9.3005
R3177 VDDD.n1597 VDDD.n1394 9.3005
R3178 VDDD.n1596 VDDD.n1595 9.3005
R3179 VDDD.n1593 VDDD.n1395 9.3005
R3180 VDDD.n1592 VDDD.n1591 9.3005
R3181 VDDD.n1590 VDDD.n1397 9.3005
R3182 VDDD.n1589 VDDD.n1588 9.3005
R3183 VDDD.n1587 VDDD.n1398 9.3005
R3184 VDDD.n1586 VDDD.n1585 9.3005
R3185 VDDD.n1584 VDDD.n1400 9.3005
R3186 VDDD.n1583 VDDD.n1582 9.3005
R3187 VDDD.n1580 VDDD.n1401 9.3005
R3188 VDDD.n1579 VDDD.n1402 9.3005
R3189 VDDD.n1578 VDDD.n1577 9.3005
R3190 VDDD.n1576 VDDD.n1403 9.3005
R3191 VDDD.n1575 VDDD.n1574 9.3005
R3192 VDDD.n1573 VDDD.n1405 9.3005
R3193 VDDD.n1572 VDDD.n1571 9.3005
R3194 VDDD.n1570 VDDD.n1406 9.3005
R3195 VDDD.n1569 VDDD.n1568 9.3005
R3196 VDDD.n1567 VDDD.n1407 9.3005
R3197 VDDD.n1566 VDDD.n1565 9.3005
R3198 VDDD.n1564 VDDD.n1408 9.3005
R3199 VDDD.n1563 VDDD.n1562 9.3005
R3200 VDDD.n1560 VDDD.n1409 9.3005
R3201 VDDD.n1559 VDDD.n1558 9.3005
R3202 VDDD.n1557 VDDD.n1411 9.3005
R3203 VDDD.n1556 VDDD.n1555 9.3005
R3204 VDDD.n1554 VDDD.n1412 9.3005
R3205 VDDD.n1553 VDDD.n1552 9.3005
R3206 VDDD.n1551 VDDD.n1414 9.3005
R3207 VDDD.n1550 VDDD.n1549 9.3005
R3208 VDDD.n1547 VDDD.n1415 9.3005
R3209 VDDD.n1546 VDDD.n1416 9.3005
R3210 VDDD.n1545 VDDD.n1544 9.3005
R3211 VDDD.n1543 VDDD.n1417 9.3005
R3212 VDDD.n1542 VDDD.n1541 9.3005
R3213 VDDD.n1540 VDDD.n1419 9.3005
R3214 VDDD.n1539 VDDD.n1538 9.3005
R3215 VDDD.n1537 VDDD.n1420 9.3005
R3216 VDDD.n1536 VDDD.n1535 9.3005
R3217 VDDD.n1534 VDDD.n1421 9.3005
R3218 VDDD.n1533 VDDD.n1532 9.3005
R3219 VDDD.n1531 VDDD.n1422 9.3005
R3220 VDDD.n1530 VDDD.n1529 9.3005
R3221 VDDD.n1527 VDDD.n1423 9.3005
R3222 VDDD.n1526 VDDD.n1525 9.3005
R3223 VDDD.n1524 VDDD.n1425 9.3005
R3224 VDDD.n1523 VDDD.n1522 9.3005
R3225 VDDD.n1521 VDDD.n1426 9.3005
R3226 VDDD.n1520 VDDD.n1519 9.3005
R3227 VDDD.n1518 VDDD.n1428 9.3005
R3228 VDDD.n1517 VDDD.n1516 9.3005
R3229 VDDD.n1514 VDDD.n1429 9.3005
R3230 VDDD.n1513 VDDD.n1430 9.3005
R3231 VDDD.n1512 VDDD.n1511 9.3005
R3232 VDDD.n1510 VDDD.n1431 9.3005
R3233 VDDD.n1509 VDDD.n1508 9.3005
R3234 VDDD.n1507 VDDD.n1433 9.3005
R3235 VDDD.n1506 VDDD.n1505 9.3005
R3236 VDDD.n1504 VDDD.n1434 9.3005
R3237 VDDD.n1503 VDDD.n1502 9.3005
R3238 VDDD.n1501 VDDD.n1435 9.3005
R3239 VDDD.n1500 VDDD.n1499 9.3005
R3240 VDDD.n1498 VDDD.n1436 9.3005
R3241 VDDD.n1497 VDDD.n1496 9.3005
R3242 VDDD.n1494 VDDD.n1437 9.3005
R3243 VDDD.n1493 VDDD.n1492 9.3005
R3244 VDDD.n1491 VDDD.n1439 9.3005
R3245 VDDD.n1490 VDDD.n1489 9.3005
R3246 VDDD.n1488 VDDD.n1440 9.3005
R3247 VDDD.n1487 VDDD.n1486 9.3005
R3248 VDDD.n1485 VDDD.n1442 9.3005
R3249 VDDD.n1484 VDDD.n1483 9.3005
R3250 VDDD.n1481 VDDD.n1443 9.3005
R3251 VDDD.n1480 VDDD.n1444 9.3005
R3252 VDDD.n1479 VDDD.n1478 9.3005
R3253 VDDD.n1477 VDDD.n1445 9.3005
R3254 VDDD.n1476 VDDD.n1475 9.3005
R3255 VDDD.n1473 VDDD.n1472 9.3005
R3256 VDDD.n1471 VDDD.n1447 9.3005
R3257 VDDD.n1470 VDDD.n1469 9.3005
R3258 VDDD.n1468 VDDD.n1448 9.3005
R3259 VDDD.n1466 VDDD.n1465 9.3005
R3260 VDDD.n1464 VDDD.n1452 9.3005
R3261 VDDD.n1463 VDDD.n1462 9.3005
R3262 VDDD.n1461 VDDD.n1453 9.3005
R3263 VDDD.n1460 VDDD.n1459 9.3005
R3264 VDDD.n1300 VDDD.n1299 9.3005
R3265 VDDD.n1303 VDDD.n1302 9.3005
R3266 VDDD.n1301 VDDD.n1009 9.3005
R3267 VDDD.n1298 VDDD.n1011 9.3005
R3268 VDDD.n1297 VDDD.n1296 9.3005
R3269 VDDD.n1293 VDDD.n1012 9.3005
R3270 VDDD.n1291 VDDD.n1290 9.3005
R3271 VDDD.n1289 VDDD.n1013 9.3005
R3272 VDDD.n1288 VDDD.n1287 9.3005
R3273 VDDD.n1284 VDDD.n1014 9.3005
R3274 VDDD.n1283 VDDD.n1282 9.3005
R3275 VDDD.n1281 VDDD.n1015 9.3005
R3276 VDDD.n1280 VDDD.n1279 9.3005
R3277 VDDD.n1276 VDDD.n1016 9.3005
R3278 VDDD.n1275 VDDD.n1274 9.3005
R3279 VDDD.n1273 VDDD.n1018 9.3005
R3280 VDDD.n1272 VDDD.n1271 9.3005
R3281 VDDD.n1268 VDDD.n1019 9.3005
R3282 VDDD.n1267 VDDD.n1266 9.3005
R3283 VDDD.n1106 VDDD.n1091 9.3005
R3284 VDDD.n1111 VDDD.n1110 9.3005
R3285 VDDD.n1112 VDDD.n1090 9.3005
R3286 VDDD.n1114 VDDD.n1113 9.3005
R3287 VDDD.n1116 VDDD.n1115 9.3005
R3288 VDDD.n1117 VDDD.n1089 9.3005
R3289 VDDD.n1119 VDDD.n1118 9.3005
R3290 VDDD.n1120 VDDD.n1087 9.3005
R3291 VDDD.n1124 VDDD.n1123 9.3005
R3292 VDDD.n1125 VDDD.n1086 9.3005
R3293 VDDD.n1127 VDDD.n1126 9.3005
R3294 VDDD.n1128 VDDD.n1084 9.3005
R3295 VDDD.n1130 VDDD.n1129 9.3005
R3296 VDDD.n1132 VDDD.n1131 9.3005
R3297 VDDD.n1133 VDDD.n1081 9.3005
R3298 VDDD.n1135 VDDD.n1134 9.3005
R3299 VDDD.n1137 VDDD.n1136 9.3005
R3300 VDDD.n1138 VDDD.n1078 9.3005
R3301 VDDD.n1140 VDDD.n1139 9.3005
R3302 VDDD.n1141 VDDD.n1077 9.3005
R3303 VDDD.n1143 VDDD.n1142 9.3005
R3304 VDDD.n1146 VDDD.n1075 9.3005
R3305 VDDD.n1148 VDDD.n1147 9.3005
R3306 VDDD.n1149 VDDD.n1074 9.3005
R3307 VDDD.n1151 VDDD.n1150 9.3005
R3308 VDDD.n1153 VDDD.n1152 9.3005
R3309 VDDD.n1154 VDDD.n1072 9.3005
R3310 VDDD.n1156 VDDD.n1155 9.3005
R3311 VDDD.n1157 VDDD.n1070 9.3005
R3312 VDDD.n1161 VDDD.n1160 9.3005
R3313 VDDD.n1162 VDDD.n1069 9.3005
R3314 VDDD.n1164 VDDD.n1163 9.3005
R3315 VDDD.n1165 VDDD.n1067 9.3005
R3316 VDDD.n1167 VDDD.n1166 9.3005
R3317 VDDD.n1169 VDDD.n1168 9.3005
R3318 VDDD.n1170 VDDD.n1064 9.3005
R3319 VDDD.n1172 VDDD.n1171 9.3005
R3320 VDDD.n1174 VDDD.n1173 9.3005
R3321 VDDD.n1175 VDDD.n1061 9.3005
R3322 VDDD.n1177 VDDD.n1176 9.3005
R3323 VDDD.n1178 VDDD.n1060 9.3005
R3324 VDDD.n1180 VDDD.n1179 9.3005
R3325 VDDD.n1183 VDDD.n1058 9.3005
R3326 VDDD.n1185 VDDD.n1184 9.3005
R3327 VDDD.n1186 VDDD.n1057 9.3005
R3328 VDDD.n1188 VDDD.n1187 9.3005
R3329 VDDD.n1190 VDDD.n1189 9.3005
R3330 VDDD.n1191 VDDD.n1055 9.3005
R3331 VDDD.n1193 VDDD.n1192 9.3005
R3332 VDDD.n1194 VDDD.n1053 9.3005
R3333 VDDD.n1198 VDDD.n1197 9.3005
R3334 VDDD.n1199 VDDD.n1052 9.3005
R3335 VDDD.n1201 VDDD.n1200 9.3005
R3336 VDDD.n1202 VDDD.n1050 9.3005
R3337 VDDD.n1204 VDDD.n1203 9.3005
R3338 VDDD.n1206 VDDD.n1205 9.3005
R3339 VDDD.n1207 VDDD.n1047 9.3005
R3340 VDDD.n1209 VDDD.n1208 9.3005
R3341 VDDD.n1211 VDDD.n1210 9.3005
R3342 VDDD.n1212 VDDD.n1044 9.3005
R3343 VDDD.n1214 VDDD.n1213 9.3005
R3344 VDDD.n1215 VDDD.n1043 9.3005
R3345 VDDD.n1217 VDDD.n1216 9.3005
R3346 VDDD.n1220 VDDD.n1041 9.3005
R3347 VDDD.n1222 VDDD.n1221 9.3005
R3348 VDDD.n1223 VDDD.n1040 9.3005
R3349 VDDD.n1225 VDDD.n1224 9.3005
R3350 VDDD.n1227 VDDD.n1226 9.3005
R3351 VDDD.n1228 VDDD.n1038 9.3005
R3352 VDDD.n1230 VDDD.n1229 9.3005
R3353 VDDD.n1231 VDDD.n1036 9.3005
R3354 VDDD.n1235 VDDD.n1234 9.3005
R3355 VDDD.n1236 VDDD.n1035 9.3005
R3356 VDDD.n1238 VDDD.n1237 9.3005
R3357 VDDD.n1239 VDDD.n1033 9.3005
R3358 VDDD.n1241 VDDD.n1240 9.3005
R3359 VDDD.n1243 VDDD.n1242 9.3005
R3360 VDDD.n1244 VDDD.n1030 9.3005
R3361 VDDD.n1246 VDDD.n1245 9.3005
R3362 VDDD.n1248 VDDD.n1247 9.3005
R3363 VDDD.n1249 VDDD.n1027 9.3005
R3364 VDDD.n1251 VDDD.n1250 9.3005
R3365 VDDD.n1252 VDDD.n1026 9.3005
R3366 VDDD.n1254 VDDD.n1253 9.3005
R3367 VDDD.n1257 VDDD.n1024 9.3005
R3368 VDDD.n1259 VDDD.n1258 9.3005
R3369 VDDD.n1260 VDDD.n1023 9.3005
R3370 VDDD.n1262 VDDD.n1261 9.3005
R3371 VDDD.n1264 VDDD.n1263 9.3005
R3372 VDDD.n1265 VDDD.n1021 9.3005
R3373 VDDD.n1103 VDDD.n1102 9.3005
R3374 VDDD.n1003 VDDD.n2 9.3005
R3375 VDDD.n1002 VDDD.n1001 9.3005
R3376 VDDD.n1000 VDDD.n999 9.3005
R3377 VDDD.n998 VDDD.n6 9.3005
R3378 VDDD.n995 VDDD.n994 9.3005
R3379 VDDD.n993 VDDD.n7 9.3005
R3380 VDDD.n992 VDDD.n991 9.3005
R3381 VDDD.n988 VDDD.n8 9.3005
R3382 VDDD.n986 VDDD.n985 9.3005
R3383 VDDD.n984 VDDD.n9 9.3005
R3384 VDDD.n638 VDDD.n637 9.3005
R3385 VDDD.n639 VDDD.n134 9.3005
R3386 VDDD.n641 VDDD.n640 9.3005
R3387 VDDD.n642 VDDD.n133 9.3005
R3388 VDDD.n645 VDDD.n644 9.3005
R3389 VDDD.n646 VDDD.n132 9.3005
R3390 VDDD.n648 VDDD.n647 9.3005
R3391 VDDD.n649 VDDD.n130 9.3005
R3392 VDDD.n651 VDDD.n650 9.3005
R3393 VDDD.n652 VDDD.n129 9.3005
R3394 VDDD.n654 VDDD.n653 9.3005
R3395 VDDD.n655 VDDD.n128 9.3005
R3396 VDDD.n659 VDDD.n658 9.3005
R3397 VDDD.n660 VDDD.n127 9.3005
R3398 VDDD.n662 VDDD.n661 9.3005
R3399 VDDD.n663 VDDD.n126 9.3005
R3400 VDDD.n665 VDDD.n664 9.3005
R3401 VDDD.n666 VDDD.n125 9.3005
R3402 VDDD.n668 VDDD.n667 9.3005
R3403 VDDD.n670 VDDD.n124 9.3005
R3404 VDDD.n672 VDDD.n671 9.3005
R3405 VDDD.n673 VDDD.n123 9.3005
R3406 VDDD.n675 VDDD.n674 9.3005
R3407 VDDD.n676 VDDD.n122 9.3005
R3408 VDDD.n679 VDDD.n678 9.3005
R3409 VDDD.n680 VDDD.n120 9.3005
R3410 VDDD.n682 VDDD.n681 9.3005
R3411 VDDD.n683 VDDD.n119 9.3005
R3412 VDDD.n685 VDDD.n684 9.3005
R3413 VDDD.n686 VDDD.n118 9.3005
R3414 VDDD.n688 VDDD.n687 9.3005
R3415 VDDD.n689 VDDD.n117 9.3005
R3416 VDDD.n691 VDDD.n690 9.3005
R3417 VDDD.n693 VDDD.n692 9.3005
R3418 VDDD.n694 VDDD.n114 9.3005
R3419 VDDD.n696 VDDD.n695 9.3005
R3420 VDDD.n697 VDDD.n113 9.3005
R3421 VDDD.n699 VDDD.n698 9.3005
R3422 VDDD.n700 VDDD.n112 9.3005
R3423 VDDD.n702 VDDD.n701 9.3005
R3424 VDDD.n703 VDDD.n111 9.3005
R3425 VDDD.n705 VDDD.n704 9.3005
R3426 VDDD.n707 VDDD.n706 9.3005
R3427 VDDD.n708 VDDD.n109 9.3005
R3428 VDDD.n710 VDDD.n709 9.3005
R3429 VDDD.n711 VDDD.n108 9.3005
R3430 VDDD.n714 VDDD.n713 9.3005
R3431 VDDD.n715 VDDD.n107 9.3005
R3432 VDDD.n717 VDDD.n716 9.3005
R3433 VDDD.n718 VDDD.n105 9.3005
R3434 VDDD.n720 VDDD.n719 9.3005
R3435 VDDD.n721 VDDD.n104 9.3005
R3436 VDDD.n723 VDDD.n722 9.3005
R3437 VDDD.n724 VDDD.n103 9.3005
R3438 VDDD.n728 VDDD.n727 9.3005
R3439 VDDD.n729 VDDD.n102 9.3005
R3440 VDDD.n731 VDDD.n730 9.3005
R3441 VDDD.n732 VDDD.n101 9.3005
R3442 VDDD.n734 VDDD.n733 9.3005
R3443 VDDD.n735 VDDD.n100 9.3005
R3444 VDDD.n737 VDDD.n736 9.3005
R3445 VDDD.n739 VDDD.n99 9.3005
R3446 VDDD.n741 VDDD.n740 9.3005
R3447 VDDD.n742 VDDD.n98 9.3005
R3448 VDDD.n744 VDDD.n743 9.3005
R3449 VDDD.n745 VDDD.n97 9.3005
R3450 VDDD.n748 VDDD.n747 9.3005
R3451 VDDD.n749 VDDD.n95 9.3005
R3452 VDDD.n751 VDDD.n750 9.3005
R3453 VDDD.n752 VDDD.n94 9.3005
R3454 VDDD.n754 VDDD.n753 9.3005
R3455 VDDD.n755 VDDD.n93 9.3005
R3456 VDDD.n757 VDDD.n756 9.3005
R3457 VDDD.n758 VDDD.n92 9.3005
R3458 VDDD.n760 VDDD.n759 9.3005
R3459 VDDD.n762 VDDD.n761 9.3005
R3460 VDDD.n763 VDDD.n89 9.3005
R3461 VDDD.n765 VDDD.n764 9.3005
R3462 VDDD.n766 VDDD.n88 9.3005
R3463 VDDD.n768 VDDD.n767 9.3005
R3464 VDDD.n769 VDDD.n87 9.3005
R3465 VDDD.n771 VDDD.n770 9.3005
R3466 VDDD.n772 VDDD.n86 9.3005
R3467 VDDD.n774 VDDD.n773 9.3005
R3468 VDDD.n776 VDDD.n775 9.3005
R3469 VDDD.n777 VDDD.n84 9.3005
R3470 VDDD.n779 VDDD.n778 9.3005
R3471 VDDD.n780 VDDD.n83 9.3005
R3472 VDDD.n783 VDDD.n782 9.3005
R3473 VDDD.n784 VDDD.n82 9.3005
R3474 VDDD.n786 VDDD.n785 9.3005
R3475 VDDD.n787 VDDD.n80 9.3005
R3476 VDDD.n789 VDDD.n788 9.3005
R3477 VDDD.n790 VDDD.n79 9.3005
R3478 VDDD.n792 VDDD.n791 9.3005
R3479 VDDD.n793 VDDD.n78 9.3005
R3480 VDDD.n797 VDDD.n796 9.3005
R3481 VDDD.n798 VDDD.n77 9.3005
R3482 VDDD.n800 VDDD.n799 9.3005
R3483 VDDD.n801 VDDD.n76 9.3005
R3484 VDDD.n803 VDDD.n802 9.3005
R3485 VDDD.n804 VDDD.n75 9.3005
R3486 VDDD.n806 VDDD.n805 9.3005
R3487 VDDD.n808 VDDD.n74 9.3005
R3488 VDDD.n810 VDDD.n809 9.3005
R3489 VDDD.n811 VDDD.n73 9.3005
R3490 VDDD.n813 VDDD.n812 9.3005
R3491 VDDD.n814 VDDD.n72 9.3005
R3492 VDDD.n817 VDDD.n816 9.3005
R3493 VDDD.n818 VDDD.n70 9.3005
R3494 VDDD.n820 VDDD.n819 9.3005
R3495 VDDD.n821 VDDD.n69 9.3005
R3496 VDDD.n823 VDDD.n822 9.3005
R3497 VDDD.n824 VDDD.n68 9.3005
R3498 VDDD.n826 VDDD.n825 9.3005
R3499 VDDD.n827 VDDD.n67 9.3005
R3500 VDDD.n829 VDDD.n828 9.3005
R3501 VDDD.n831 VDDD.n830 9.3005
R3502 VDDD.n832 VDDD.n64 9.3005
R3503 VDDD.n834 VDDD.n833 9.3005
R3504 VDDD.n835 VDDD.n63 9.3005
R3505 VDDD.n837 VDDD.n836 9.3005
R3506 VDDD.n838 VDDD.n62 9.3005
R3507 VDDD.n840 VDDD.n839 9.3005
R3508 VDDD.n841 VDDD.n61 9.3005
R3509 VDDD.n843 VDDD.n842 9.3005
R3510 VDDD.n845 VDDD.n844 9.3005
R3511 VDDD.n846 VDDD.n59 9.3005
R3512 VDDD.n848 VDDD.n847 9.3005
R3513 VDDD.n849 VDDD.n58 9.3005
R3514 VDDD.n852 VDDD.n851 9.3005
R3515 VDDD.n853 VDDD.n57 9.3005
R3516 VDDD.n855 VDDD.n854 9.3005
R3517 VDDD.n856 VDDD.n55 9.3005
R3518 VDDD.n858 VDDD.n857 9.3005
R3519 VDDD.n859 VDDD.n54 9.3005
R3520 VDDD.n861 VDDD.n860 9.3005
R3521 VDDD.n862 VDDD.n53 9.3005
R3522 VDDD.n866 VDDD.n865 9.3005
R3523 VDDD.n867 VDDD.n52 9.3005
R3524 VDDD.n869 VDDD.n868 9.3005
R3525 VDDD.n870 VDDD.n51 9.3005
R3526 VDDD.n872 VDDD.n871 9.3005
R3527 VDDD.n873 VDDD.n50 9.3005
R3528 VDDD.n875 VDDD.n874 9.3005
R3529 VDDD.n877 VDDD.n49 9.3005
R3530 VDDD.n879 VDDD.n878 9.3005
R3531 VDDD.n880 VDDD.n48 9.3005
R3532 VDDD.n882 VDDD.n881 9.3005
R3533 VDDD.n883 VDDD.n47 9.3005
R3534 VDDD.n886 VDDD.n885 9.3005
R3535 VDDD.n887 VDDD.n45 9.3005
R3536 VDDD.n889 VDDD.n888 9.3005
R3537 VDDD.n890 VDDD.n44 9.3005
R3538 VDDD.n892 VDDD.n891 9.3005
R3539 VDDD.n893 VDDD.n43 9.3005
R3540 VDDD.n895 VDDD.n894 9.3005
R3541 VDDD.n896 VDDD.n42 9.3005
R3542 VDDD.n898 VDDD.n897 9.3005
R3543 VDDD.n900 VDDD.n899 9.3005
R3544 VDDD.n901 VDDD.n39 9.3005
R3545 VDDD.n903 VDDD.n902 9.3005
R3546 VDDD.n904 VDDD.n38 9.3005
R3547 VDDD.n906 VDDD.n905 9.3005
R3548 VDDD.n907 VDDD.n37 9.3005
R3549 VDDD.n909 VDDD.n908 9.3005
R3550 VDDD.n910 VDDD.n36 9.3005
R3551 VDDD.n912 VDDD.n911 9.3005
R3552 VDDD.n914 VDDD.n913 9.3005
R3553 VDDD.n915 VDDD.n34 9.3005
R3554 VDDD.n917 VDDD.n916 9.3005
R3555 VDDD.n918 VDDD.n33 9.3005
R3556 VDDD.n921 VDDD.n920 9.3005
R3557 VDDD.n922 VDDD.n32 9.3005
R3558 VDDD.n924 VDDD.n923 9.3005
R3559 VDDD.n925 VDDD.n30 9.3005
R3560 VDDD.n927 VDDD.n926 9.3005
R3561 VDDD.n928 VDDD.n29 9.3005
R3562 VDDD.n930 VDDD.n929 9.3005
R3563 VDDD.n931 VDDD.n28 9.3005
R3564 VDDD.n935 VDDD.n934 9.3005
R3565 VDDD.n936 VDDD.n27 9.3005
R3566 VDDD.n938 VDDD.n937 9.3005
R3567 VDDD.n939 VDDD.n26 9.3005
R3568 VDDD.n941 VDDD.n940 9.3005
R3569 VDDD.n942 VDDD.n25 9.3005
R3570 VDDD.n944 VDDD.n943 9.3005
R3571 VDDD.n946 VDDD.n24 9.3005
R3572 VDDD.n948 VDDD.n947 9.3005
R3573 VDDD.n949 VDDD.n23 9.3005
R3574 VDDD.n951 VDDD.n950 9.3005
R3575 VDDD.n952 VDDD.n22 9.3005
R3576 VDDD.n955 VDDD.n954 9.3005
R3577 VDDD.n956 VDDD.n20 9.3005
R3578 VDDD.n958 VDDD.n957 9.3005
R3579 VDDD.n959 VDDD.n19 9.3005
R3580 VDDD.n961 VDDD.n960 9.3005
R3581 VDDD.n962 VDDD.n18 9.3005
R3582 VDDD.n964 VDDD.n963 9.3005
R3583 VDDD.n965 VDDD.n17 9.3005
R3584 VDDD.n967 VDDD.n966 9.3005
R3585 VDDD.n969 VDDD.n968 9.3005
R3586 VDDD.n970 VDDD.n14 9.3005
R3587 VDDD.n972 VDDD.n971 9.3005
R3588 VDDD.n973 VDDD.n13 9.3005
R3589 VDDD.n975 VDDD.n974 9.3005
R3590 VDDD.n976 VDDD.n12 9.3005
R3591 VDDD.n978 VDDD.n977 9.3005
R3592 VDDD.n979 VDDD.n11 9.3005
R3593 VDDD.n981 VDDD.n980 9.3005
R3594 VDDD.n983 VDDD.n982 9.3005
R3595 VDDD.n636 VDDD.n635 9.3005
R3596 VDDD.n634 VDDD.n135 9.3005
R3597 VDDD.n633 VDDD.n632 9.3005
R3598 VDDD.n631 VDDD.n136 9.3005
R3599 VDDD.n630 VDDD.n629 9.3005
R3600 VDDD.n628 VDDD.n137 9.3005
R3601 VDDD.n626 VDDD.n625 9.3005
R3602 VDDD.n624 VDDD.n139 9.3005
R3603 VDDD.n623 VDDD.n622 9.3005
R3604 VDDD.n621 VDDD.n140 9.3005
R3605 VDDD.n620 VDDD.n619 9.3005
R3606 VDDD.n618 VDDD.n141 9.3005
R3607 VDDD.n617 VDDD.n616 9.3005
R3608 VDDD.n615 VDDD.n142 9.3005
R3609 VDDD.n614 VDDD.n613 9.3005
R3610 VDDD.n612 VDDD.n145 9.3005
R3611 VDDD.n611 VDDD.n610 9.3005
R3612 VDDD.n609 VDDD.n146 9.3005
R3613 VDDD.n608 VDDD.n607 9.3005
R3614 VDDD.n606 VDDD.n148 9.3005
R3615 VDDD.n605 VDDD.n604 9.3005
R3616 VDDD.n603 VDDD.n602 9.3005
R3617 VDDD.n601 VDDD.n149 9.3005
R3618 VDDD.n600 VDDD.n599 9.3005
R3619 VDDD.n598 VDDD.n150 9.3005
R3620 VDDD.n596 VDDD.n595 9.3005
R3621 VDDD.n594 VDDD.n152 9.3005
R3622 VDDD.n593 VDDD.n592 9.3005
R3623 VDDD.n591 VDDD.n153 9.3005
R3624 VDDD.n590 VDDD.n589 9.3005
R3625 VDDD.n588 VDDD.n154 9.3005
R3626 VDDD.n587 VDDD.n586 9.3005
R3627 VDDD.n585 VDDD.n155 9.3005
R3628 VDDD.n582 VDDD.n581 9.3005
R3629 VDDD.n580 VDDD.n156 9.3005
R3630 VDDD.n579 VDDD.n578 9.3005
R3631 VDDD.n577 VDDD.n157 9.3005
R3632 VDDD.n576 VDDD.n575 9.3005
R3633 VDDD.n574 VDDD.n158 9.3005
R3634 VDDD.n573 VDDD.n572 9.3005
R3635 VDDD.n571 VDDD.n159 9.3005
R3636 VDDD.n569 VDDD.n568 9.3005
R3637 VDDD.n567 VDDD.n160 9.3005
R3638 VDDD.n566 VDDD.n565 9.3005
R3639 VDDD.n564 VDDD.n161 9.3005
R3640 VDDD.n563 VDDD.n562 9.3005
R3641 VDDD.n561 VDDD.n560 9.3005
R3642 VDDD.n559 VDDD.n163 9.3005
R3643 VDDD.n557 VDDD.n556 9.3005
R3644 VDDD.n555 VDDD.n164 9.3005
R3645 VDDD.n554 VDDD.n553 9.3005
R3646 VDDD.n552 VDDD.n165 9.3005
R3647 VDDD.n551 VDDD.n550 9.3005
R3648 VDDD.n549 VDDD.n166 9.3005
R3649 VDDD.n548 VDDD.n547 9.3005
R3650 VDDD.n546 VDDD.n167 9.3005
R3651 VDDD.n545 VDDD.n544 9.3005
R3652 VDDD.n543 VDDD.n170 9.3005
R3653 VDDD.n542 VDDD.n541 9.3005
R3654 VDDD.n540 VDDD.n171 9.3005
R3655 VDDD.n539 VDDD.n538 9.3005
R3656 VDDD.n537 VDDD.n173 9.3005
R3657 VDDD.n536 VDDD.n535 9.3005
R3658 VDDD.n534 VDDD.n533 9.3005
R3659 VDDD.n532 VDDD.n174 9.3005
R3660 VDDD.n531 VDDD.n530 9.3005
R3661 VDDD.n529 VDDD.n175 9.3005
R3662 VDDD.n527 VDDD.n526 9.3005
R3663 VDDD.n525 VDDD.n177 9.3005
R3664 VDDD.n524 VDDD.n523 9.3005
R3665 VDDD.n522 VDDD.n178 9.3005
R3666 VDDD.n521 VDDD.n520 9.3005
R3667 VDDD.n519 VDDD.n179 9.3005
R3668 VDDD.n518 VDDD.n517 9.3005
R3669 VDDD.n516 VDDD.n180 9.3005
R3670 VDDD.n513 VDDD.n512 9.3005
R3671 VDDD.n511 VDDD.n181 9.3005
R3672 VDDD.n510 VDDD.n509 9.3005
R3673 VDDD.n508 VDDD.n182 9.3005
R3674 VDDD.n507 VDDD.n506 9.3005
R3675 VDDD.n505 VDDD.n183 9.3005
R3676 VDDD.n504 VDDD.n503 9.3005
R3677 VDDD.n502 VDDD.n184 9.3005
R3678 VDDD.n500 VDDD.n499 9.3005
R3679 VDDD.n498 VDDD.n185 9.3005
R3680 VDDD.n497 VDDD.n496 9.3005
R3681 VDDD.n495 VDDD.n186 9.3005
R3682 VDDD.n494 VDDD.n493 9.3005
R3683 VDDD.n492 VDDD.n491 9.3005
R3684 VDDD.n490 VDDD.n188 9.3005
R3685 VDDD.n488 VDDD.n487 9.3005
R3686 VDDD.n486 VDDD.n189 9.3005
R3687 VDDD.n485 VDDD.n484 9.3005
R3688 VDDD.n483 VDDD.n190 9.3005
R3689 VDDD.n482 VDDD.n481 9.3005
R3690 VDDD.n480 VDDD.n191 9.3005
R3691 VDDD.n479 VDDD.n478 9.3005
R3692 VDDD.n477 VDDD.n192 9.3005
R3693 VDDD.n476 VDDD.n475 9.3005
R3694 VDDD.n474 VDDD.n195 9.3005
R3695 VDDD.n473 VDDD.n472 9.3005
R3696 VDDD.n471 VDDD.n196 9.3005
R3697 VDDD.n470 VDDD.n469 9.3005
R3698 VDDD.n468 VDDD.n198 9.3005
R3699 VDDD.n467 VDDD.n466 9.3005
R3700 VDDD.n465 VDDD.n464 9.3005
R3701 VDDD.n463 VDDD.n199 9.3005
R3702 VDDD.n462 VDDD.n461 9.3005
R3703 VDDD.n460 VDDD.n200 9.3005
R3704 VDDD.n458 VDDD.n457 9.3005
R3705 VDDD.n456 VDDD.n202 9.3005
R3706 VDDD.n455 VDDD.n454 9.3005
R3707 VDDD.n453 VDDD.n203 9.3005
R3708 VDDD.n452 VDDD.n451 9.3005
R3709 VDDD.n450 VDDD.n204 9.3005
R3710 VDDD.n449 VDDD.n448 9.3005
R3711 VDDD.n447 VDDD.n205 9.3005
R3712 VDDD.n444 VDDD.n443 9.3005
R3713 VDDD.n442 VDDD.n206 9.3005
R3714 VDDD.n441 VDDD.n440 9.3005
R3715 VDDD.n439 VDDD.n207 9.3005
R3716 VDDD.n438 VDDD.n437 9.3005
R3717 VDDD.n436 VDDD.n208 9.3005
R3718 VDDD.n435 VDDD.n434 9.3005
R3719 VDDD.n433 VDDD.n209 9.3005
R3720 VDDD.n431 VDDD.n430 9.3005
R3721 VDDD.n429 VDDD.n210 9.3005
R3722 VDDD.n428 VDDD.n427 9.3005
R3723 VDDD.n426 VDDD.n211 9.3005
R3724 VDDD.n425 VDDD.n424 9.3005
R3725 VDDD.n423 VDDD.n422 9.3005
R3726 VDDD.n421 VDDD.n213 9.3005
R3727 VDDD.n419 VDDD.n418 9.3005
R3728 VDDD.n417 VDDD.n214 9.3005
R3729 VDDD.n416 VDDD.n415 9.3005
R3730 VDDD.n414 VDDD.n215 9.3005
R3731 VDDD.n413 VDDD.n412 9.3005
R3732 VDDD.n411 VDDD.n216 9.3005
R3733 VDDD.n410 VDDD.n409 9.3005
R3734 VDDD.n408 VDDD.n217 9.3005
R3735 VDDD.n407 VDDD.n406 9.3005
R3736 VDDD.n405 VDDD.n220 9.3005
R3737 VDDD.n404 VDDD.n403 9.3005
R3738 VDDD.n402 VDDD.n221 9.3005
R3739 VDDD.n401 VDDD.n400 9.3005
R3740 VDDD.n399 VDDD.n223 9.3005
R3741 VDDD.n398 VDDD.n397 9.3005
R3742 VDDD.n396 VDDD.n395 9.3005
R3743 VDDD.n394 VDDD.n224 9.3005
R3744 VDDD.n393 VDDD.n392 9.3005
R3745 VDDD.n391 VDDD.n225 9.3005
R3746 VDDD.n389 VDDD.n388 9.3005
R3747 VDDD.n387 VDDD.n227 9.3005
R3748 VDDD.n386 VDDD.n385 9.3005
R3749 VDDD.n384 VDDD.n228 9.3005
R3750 VDDD.n383 VDDD.n382 9.3005
R3751 VDDD.n381 VDDD.n229 9.3005
R3752 VDDD.n380 VDDD.n379 9.3005
R3753 VDDD.n378 VDDD.n230 9.3005
R3754 VDDD.n375 VDDD.n374 9.3005
R3755 VDDD.n373 VDDD.n231 9.3005
R3756 VDDD.n372 VDDD.n371 9.3005
R3757 VDDD.n370 VDDD.n232 9.3005
R3758 VDDD.n369 VDDD.n368 9.3005
R3759 VDDD.n367 VDDD.n233 9.3005
R3760 VDDD.n366 VDDD.n365 9.3005
R3761 VDDD.n364 VDDD.n234 9.3005
R3762 VDDD.n362 VDDD.n361 9.3005
R3763 VDDD.n360 VDDD.n235 9.3005
R3764 VDDD.n359 VDDD.n358 9.3005
R3765 VDDD.n357 VDDD.n236 9.3005
R3766 VDDD.n356 VDDD.n355 9.3005
R3767 VDDD.n354 VDDD.n353 9.3005
R3768 VDDD.n352 VDDD.n238 9.3005
R3769 VDDD.n350 VDDD.n349 9.3005
R3770 VDDD.n348 VDDD.n239 9.3005
R3771 VDDD.n347 VDDD.n346 9.3005
R3772 VDDD.n345 VDDD.n240 9.3005
R3773 VDDD.n344 VDDD.n343 9.3005
R3774 VDDD.n342 VDDD.n241 9.3005
R3775 VDDD.n341 VDDD.n340 9.3005
R3776 VDDD.n339 VDDD.n242 9.3005
R3777 VDDD.n338 VDDD.n337 9.3005
R3778 VDDD.n336 VDDD.n245 9.3005
R3779 VDDD.n335 VDDD.n334 9.3005
R3780 VDDD.n333 VDDD.n246 9.3005
R3781 VDDD.n332 VDDD.n331 9.3005
R3782 VDDD.n330 VDDD.n248 9.3005
R3783 VDDD.n329 VDDD.n328 9.3005
R3784 VDDD.n327 VDDD.n326 9.3005
R3785 VDDD.n325 VDDD.n249 9.3005
R3786 VDDD.n324 VDDD.n323 9.3005
R3787 VDDD.n322 VDDD.n250 9.3005
R3788 VDDD.n320 VDDD.n319 9.3005
R3789 VDDD.n318 VDDD.n252 9.3005
R3790 VDDD.n317 VDDD.n316 9.3005
R3791 VDDD.n315 VDDD.n253 9.3005
R3792 VDDD.n314 VDDD.n313 9.3005
R3793 VDDD.n312 VDDD.n254 9.3005
R3794 VDDD.n311 VDDD.n310 9.3005
R3795 VDDD.n309 VDDD.n255 9.3005
R3796 VDDD.n306 VDDD.n305 9.3005
R3797 VDDD.n304 VDDD.n256 9.3005
R3798 VDDD.n303 VDDD.n302 9.3005
R3799 VDDD.n301 VDDD.n257 9.3005
R3800 VDDD.n300 VDDD.n299 9.3005
R3801 VDDD.n298 VDDD.n258 9.3005
R3802 VDDD.n297 VDDD.n296 9.3005
R3803 VDDD.n295 VDDD.n259 9.3005
R3804 VDDD.n293 VDDD.n292 9.3005
R3805 VDDD.n291 VDDD.n260 9.3005
R3806 VDDD.n290 VDDD.n289 9.3005
R3807 VDDD.n288 VDDD.n261 9.3005
R3808 VDDD.n287 VDDD.n285 9.3005
R3809 VDDD.n284 VDDD.n262 9.3005
R3810 VDDD.n283 VDDD.n282 9.3005
R3811 VDDD.n281 VDDD.n263 9.3005
R3812 VDDD.n278 VDDD.n277 9.3005
R3813 VDDD.n276 VDDD.n266 9.3005
R3814 VDDD.n275 VDDD.n274 9.3005
R3815 VDDD.n273 VDDD.n267 9.3005
R3816 VDDD.n321 VDDD.n320 9.03579
R3817 VDDD.n353 VDDD.n237 9.03579
R3818 VDDD.n390 VDDD.n389 9.03579
R3819 VDDD.n422 VDDD.n212 9.03579
R3820 VDDD.n459 VDDD.n458 9.03579
R3821 VDDD.n491 VDDD.n187 9.03579
R3822 VDDD.n528 VDDD.n527 9.03579
R3823 VDDD.n560 VDDD.n162 9.03579
R3824 VDDD.n597 VDDD.n596 9.03579
R3825 VDDD.n629 VDDD.n138 9.03579
R3826 VDDD.n644 VDDD.n643 9.03579
R3827 VDDD.n677 VDDD.n120 9.03579
R3828 VDDD.n713 VDDD.n712 9.03579
R3829 VDDD.n746 VDDD.n95 9.03579
R3830 VDDD.n782 VDDD.n781 9.03579
R3831 VDDD.n815 VDDD.n70 9.03579
R3832 VDDD.n851 VDDD.n850 9.03579
R3833 VDDD.n884 VDDD.n45 9.03579
R3834 VDDD.n920 VDDD.n919 9.03579
R3835 VDDD.n953 VDDD.n20 9.03579
R3836 VDDD.n2448 VDDD.n2188 9.03579
R3837 VDDD.n2414 VDDD.n2413 9.03579
R3838 VDDD.n2381 VDDD.n2380 9.03579
R3839 VDDD.n2348 VDDD.n2347 9.03579
R3840 VDDD.n2315 VDDD.n2314 9.03579
R3841 VDDD.n2282 VDDD.n2281 9.03579
R3842 VDDD.n2152 VDDD.n1896 9.03579
R3843 VDDD.n2118 VDDD.n2117 9.03579
R3844 VDDD.n2085 VDDD.n2084 9.03579
R3845 VDDD.n2052 VDDD.n2051 9.03579
R3846 VDDD.n2019 VDDD.n2018 9.03579
R3847 VDDD.n1986 VDDD.n1985 9.03579
R3848 VDDD.n1615 VDDD.n1614 9.03579
R3849 VDDD.n1582 VDDD.n1581 9.03579
R3850 VDDD.n1549 VDDD.n1548 9.03579
R3851 VDDD.n1516 VDDD.n1515 9.03579
R3852 VDDD.n1483 VDDD.n1482 9.03579
R3853 VDDD.n1806 VDDD.n1317 9.03579
R3854 VDDD.n1772 VDDD.n1771 9.03579
R3855 VDDD.n1739 VDDD.n1738 9.03579
R3856 VDDD.n1706 VDDD.n1705 9.03579
R3857 VDDD.n1673 VDDD.n1672 9.03579
R3858 VDDD.n1869 VDDD.n1868 8.65932
R3859 VDDD.n2274 VDDD.n2273 8.28285
R3860 VDDD.n2489 VDDD.n1006 8.19295
R3861 VDDD.n1123 VDDD.n1122 7.15344
R3862 VDDD.n1144 VDDD.n1143 7.15344
R3863 VDDD.n1160 VDDD.n1159 7.15344
R3864 VDDD.n1181 VDDD.n1180 7.15344
R3865 VDDD.n1197 VDDD.n1196 7.15344
R3866 VDDD.n1218 VDDD.n1217 7.15344
R3867 VDDD.n1234 VDDD.n1233 7.15344
R3868 VDDD.n1255 VDDD.n1254 7.15344
R3869 VDDD.n1271 VDDD.n1270 7.15344
R3870 VDDD.n1296 VDDD.n1295 7.15344
R3871 VDDD.n2472 VDDD.n2471 7.12063
R3872 VDDD.n2176 VDDD.n2175 7.12063
R3873 VDDD.n1830 VDDD.n1829 7.12063
R3874 VDDD.n1458 VDDD.n1457 6.94395
R3875 VDDD.n269 VDDD.n266 6.77697
R3876 VDDD.n999 VDDD.n5 6.77697
R3877 VDDD.n1469 VDDD.n1450 6.77697
R3878 VDDD.n2488 VDDD.n1007 6.50081
R3879 VDDD.n265 VDDD.n262 6.4005
R3880 VDDD.n991 VDDD.n990 6.4005
R3881 VDDD.n1462 VDDD.n1455 6.4005
R3882 VDDD.n1110 VDDD.n1109 6.4005
R3883 VDDD.n308 VDDD.n306 6.02403
R3884 VDDD.n340 VDDD.n244 6.02403
R3885 VDDD.n377 VDDD.n375 6.02403
R3886 VDDD.n409 VDDD.n219 6.02403
R3887 VDDD.n446 VDDD.n444 6.02403
R3888 VDDD.n478 VDDD.n194 6.02403
R3889 VDDD.n515 VDDD.n513 6.02403
R3890 VDDD.n547 VDDD.n169 6.02403
R3891 VDDD.n584 VDDD.n582 6.02403
R3892 VDDD.n616 VDDD.n144 6.02403
R3893 VDDD.n658 VDDD.n657 6.02403
R3894 VDDD.n693 VDDD.n116 6.02403
R3895 VDDD.n727 VDDD.n726 6.02403
R3896 VDDD.n762 VDDD.n91 6.02403
R3897 VDDD.n796 VDDD.n795 6.02403
R3898 VDDD.n831 VDDD.n66 6.02403
R3899 VDDD.n865 VDDD.n864 6.02403
R3900 VDDD.n900 VDDD.n41 6.02403
R3901 VDDD.n934 VDDD.n933 6.02403
R3902 VDDD.n969 VDDD.n16 6.02403
R3903 VDDD.n2458 VDDD.n2182 6.02403
R3904 VDDD.n2427 VDDD.n2426 6.02403
R3905 VDDD.n2394 VDDD.n2393 6.02403
R3906 VDDD.n2361 VDDD.n2360 6.02403
R3907 VDDD.n2328 VDDD.n2327 6.02403
R3908 VDDD.n2295 VDDD.n2294 6.02403
R3909 VDDD.n2162 VDDD.n1890 6.02403
R3910 VDDD.n2131 VDDD.n2130 6.02403
R3911 VDDD.n2098 VDDD.n2097 6.02403
R3912 VDDD.n2065 VDDD.n2064 6.02403
R3913 VDDD.n2032 VDDD.n2031 6.02403
R3914 VDDD.n1999 VDDD.n1998 6.02403
R3915 VDDD.n1628 VDDD.n1627 6.02403
R3916 VDDD.n1595 VDDD.n1594 6.02403
R3917 VDDD.n1562 VDDD.n1561 6.02403
R3918 VDDD.n1529 VDDD.n1528 6.02403
R3919 VDDD.n1496 VDDD.n1495 6.02403
R3920 VDDD.n1816 VDDD.n1311 6.02403
R3921 VDDD.n1785 VDDD.n1784 6.02403
R3922 VDDD.n1752 VDDD.n1751 6.02403
R3923 VDDD.n1719 VDDD.n1718 6.02403
R3924 VDDD.n1686 VDDD.n1685 6.02403
R3925 VDDD.n1129 VDDD.n1083 6.02403
R3926 VDDD.n1137 VDDD.n1080 6.02403
R3927 VDDD.n1166 VDDD.n1066 6.02403
R3928 VDDD.n1174 VDDD.n1063 6.02403
R3929 VDDD.n1203 VDDD.n1049 6.02403
R3930 VDDD.n1211 VDDD.n1046 6.02403
R3931 VDDD.n1240 VDDD.n1032 6.02403
R3932 VDDD.n1248 VDDD.n1029 6.02403
R3933 VDDD.n1279 VDDD.n1278 6.02403
R3934 VDDD.n1287 VDDD.n1286 6.02403
R3935 VDDD.n2488 VDDD.n2487 5.8805
R3936 VDDD.n2490 VDDD.n2489 5.8805
R3937 VDDD.n2479 VDDD.n1306 5.71175
R3938 VDDD.n2477 VDDD.n1305 5.31607
R3939 VDDD.n2483 VDDD.n2482 5.02133
R3940 VDDD.n2485 VDDD.n2484 5.02003
R3941 VDDD.n2487 VDDD.n2486 4.8155
R3942 VDDD.n2484 VDDD.n1007 4.8155
R3943 VDDD.n2490 VDDD.n1 4.8155
R3944 VDDD VDDD.n1855 4.7712
R3945 VDDD.n2486 VDDD.n2485 4.5005
R3946 VDDD.n2482 VDDD.n1008 4.5005
R3947 VDDD.n2477 VDDD.n2476 4.5005
R3948 VDDD.n1304 VDDD.n1 4.5005
R3949 VDDD.n2481 VDDD.n2480 4.5005
R3950 VDDD.n2479 VDDD.n2478 4.5005
R3951 VDDD.n2474 VDDD.n1306 4.5005
R3952 VDDD.n2486 VDDD.n1008 4.38425
R3953 VDDD.n2484 VDDD.n2483 4.38425
R3954 VDDD.n2480 VDDD.n1 4.38425
R3955 VDDD.n2177 VDDD.n1885 4.29868
R3956 VDDD.n309 VDDD.n308 3.76521
R3957 VDDD.n244 VDDD.n241 3.76521
R3958 VDDD.n378 VDDD.n377 3.76521
R3959 VDDD.n219 VDDD.n216 3.76521
R3960 VDDD.n447 VDDD.n446 3.76521
R3961 VDDD.n194 VDDD.n191 3.76521
R3962 VDDD.n516 VDDD.n515 3.76521
R3963 VDDD.n169 VDDD.n166 3.76521
R3964 VDDD.n585 VDDD.n584 3.76521
R3965 VDDD.n144 VDDD.n141 3.76521
R3966 VDDD.n657 VDDD.n655 3.76521
R3967 VDDD.n690 VDDD.n116 3.76521
R3968 VDDD.n726 VDDD.n724 3.76521
R3969 VDDD.n759 VDDD.n91 3.76521
R3970 VDDD.n795 VDDD.n793 3.76521
R3971 VDDD.n828 VDDD.n66 3.76521
R3972 VDDD.n864 VDDD.n862 3.76521
R3973 VDDD.n897 VDDD.n41 3.76521
R3974 VDDD.n933 VDDD.n931 3.76521
R3975 VDDD.n966 VDDD.n16 3.76521
R3976 VDDD.n2459 VDDD.n2458 3.76521
R3977 VDDD.n2426 VDDD.n2425 3.76521
R3978 VDDD.n2393 VDDD.n2392 3.76521
R3979 VDDD.n2360 VDDD.n2359 3.76521
R3980 VDDD.n2327 VDDD.n2326 3.76521
R3981 VDDD.n2294 VDDD.n2293 3.76521
R3982 VDDD.n2163 VDDD.n2162 3.76521
R3983 VDDD.n2130 VDDD.n2129 3.76521
R3984 VDDD.n2097 VDDD.n2096 3.76521
R3985 VDDD.n2064 VDDD.n2063 3.76521
R3986 VDDD.n2031 VDDD.n2030 3.76521
R3987 VDDD.n1998 VDDD.n1997 3.76521
R3988 VDDD.n1627 VDDD.n1626 3.76521
R3989 VDDD.n1594 VDDD.n1593 3.76521
R3990 VDDD.n1561 VDDD.n1560 3.76521
R3991 VDDD.n1528 VDDD.n1527 3.76521
R3992 VDDD.n1495 VDDD.n1494 3.76521
R3993 VDDD.n1817 VDDD.n1816 3.76521
R3994 VDDD.n1784 VDDD.n1783 3.76521
R3995 VDDD.n1751 VDDD.n1750 3.76521
R3996 VDDD.n1718 VDDD.n1717 3.76521
R3997 VDDD.n1685 VDDD.n1684 3.76521
R3998 VDDD.n1007 VDDD.n0 3.63545
R3999 VDDD.n2487 VDDD.n0 3.4105
R4000 VDDD.n2491 VDDD.n2490 3.4105
R4001 VDDD.n282 VDDD.n265 3.38874
R4002 VDDD.n990 VDDD.n7 3.38874
R4003 VDDD.n1860 VDDD.n1859 3.38874
R4004 VDDD.n1455 VDDD.n1452 3.38874
R4005 VDDD.n1109 VDDD.n1090 3.38874
R4006 VDDD.n1862 VDDD.n1851 2.63579
R4007 VDDD.n1873 VDDD.n1848 1.88285
R4008 VDDD.n638 VDDD.n636 1.68279
R4009 VDDD.n2476 VDDD.n1008 1.38175
R4010 VDDD.n2483 VDDD.n1305 1.38175
R4011 VDDD.n2480 VDDD.n2479 1.38175
R4012 VDDD.n1132 VDDD.n1083 1.12991
R4013 VDDD.n1134 VDDD.n1080 1.12991
R4014 VDDD.n1169 VDDD.n1066 1.12991
R4015 VDDD.n1171 VDDD.n1063 1.12991
R4016 VDDD.n1206 VDDD.n1049 1.12991
R4017 VDDD.n1208 VDDD.n1046 1.12991
R4018 VDDD.n1243 VDDD.n1032 1.12991
R4019 VDDD.n1245 VDDD.n1029 1.12991
R4020 VDDD.n1278 VDDD.n1015 1.12991
R4021 VDDD.n1286 VDDD.n1284 1.12991
R4022 VDDD.n1654 VDDD.n1653 1.01388
R4023 VDDD.n2473 VDDD.n2177 0.96925
R4024 VDDD.n2478 VDDD.n2477 0.807877
R4025 VDDD.n273 VDDD.n272 0.753441
R4026 VDDD.n322 VDDD.n321 0.753441
R4027 VDDD.n356 VDDD.n237 0.753441
R4028 VDDD.n391 VDDD.n390 0.753441
R4029 VDDD.n425 VDDD.n212 0.753441
R4030 VDDD.n460 VDDD.n459 0.753441
R4031 VDDD.n494 VDDD.n187 0.753441
R4032 VDDD.n529 VDDD.n528 0.753441
R4033 VDDD.n563 VDDD.n162 0.753441
R4034 VDDD.n598 VDDD.n597 0.753441
R4035 VDDD.n138 VDDD.n136 0.753441
R4036 VDDD.n643 VDDD.n642 0.753441
R4037 VDDD.n678 VDDD.n677 0.753441
R4038 VDDD.n712 VDDD.n711 0.753441
R4039 VDDD.n747 VDDD.n746 0.753441
R4040 VDDD.n781 VDDD.n780 0.753441
R4041 VDDD.n816 VDDD.n815 0.753441
R4042 VDDD.n850 VDDD.n849 0.753441
R4043 VDDD.n885 VDDD.n884 0.753441
R4044 VDDD.n919 VDDD.n918 0.753441
R4045 VDDD.n954 VDDD.n953 0.753441
R4046 VDDD.n1004 VDDD.n1003 0.753441
R4047 VDDD.n2445 VDDD.n2188 0.753441
R4048 VDDD.n2413 VDDD.n2412 0.753441
R4049 VDDD.n2380 VDDD.n2379 0.753441
R4050 VDDD.n2347 VDDD.n2346 0.753441
R4051 VDDD.n2314 VDDD.n2313 0.753441
R4052 VDDD.n2281 VDDD.n2280 0.753441
R4053 VDDD.n2149 VDDD.n1896 0.753441
R4054 VDDD.n2117 VDDD.n2116 0.753441
R4055 VDDD.n2084 VDDD.n2083 0.753441
R4056 VDDD.n2051 VDDD.n2050 0.753441
R4057 VDDD.n2018 VDDD.n2017 0.753441
R4058 VDDD.n1985 VDDD.n1984 0.753441
R4059 VDDD.n1614 VDDD.n1613 0.753441
R4060 VDDD.n1581 VDDD.n1580 0.753441
R4061 VDDD.n1548 VDDD.n1547 0.753441
R4062 VDDD.n1515 VDDD.n1514 0.753441
R4063 VDDD.n1482 VDDD.n1481 0.753441
R4064 VDDD.n1474 VDDD.n1473 0.753441
R4065 VDDD.n1803 VDDD.n1317 0.753441
R4066 VDDD.n1771 VDDD.n1770 0.753441
R4067 VDDD.n1738 VDDD.n1737 0.753441
R4068 VDDD.n1705 VDDD.n1704 0.753441
R4069 VDDD.n1672 VDDD.n1671 0.753441
R4070 VDDD.n2489 VDDD.n2488 0.620813
R4071 VDDD.n2485 VDDD.n1304 0.523938
R4072 VDDD.n2475 VDDD.n2474 0.522635
R4073 VDDD.n2482 VDDD.n2481 0.520031
R4074 VDDD.n1306 VDDD 0.4705
R4075 VDDD.n2473 VDDD 0.40024
R4076 VDDD.n2177 VDDD 0.398938
R4077 VDDD.n281 VDDD.n280 0.376971
R4078 VDDD.n997 VDDD.n995 0.376971
R4079 VDDD.n1467 VDDD.n1466 0.376971
R4080 VDDD.n2491 VDDD.n0 0.227797
R4081 VDDD.n1885 VDDD 0.184094
R4082 VDDD.n1641 VDDD.n1640 0.166812
R4083 VDDD.n1667 VDDD.n1666 0.164863
R4084 VDDD.n1459 VDDD.n1458 0.150766
R4085 VDDD.n1458 VDDD 0.150327
R4086 VDDD.n2176 VDDD.n1886 0.148519
R4087 VDDD.n2472 VDDD.n2178 0.148519
R4088 VDDD.n1830 VDDD.n1307 0.148519
R4089 VDDD.n2275 VDDD.n2272 0.141672
R4090 VDDD.n1104 VDDD.n1103 0.130708
R4091 VDDD.n1857 VDDD.n1856 0.120292
R4092 VDDD.n1857 VDDD.n1852 0.120292
R4093 VDDD.n1864 VDDD.n1852 0.120292
R4094 VDDD.n1865 VDDD.n1864 0.120292
R4095 VDDD.n1866 VDDD.n1865 0.120292
R4096 VDDD.n1866 VDDD.n1849 0.120292
R4097 VDDD.n1871 VDDD.n1849 0.120292
R4098 VDDD.n1872 VDDD.n1871 0.120292
R4099 VDDD.n1876 VDDD.n1847 0.120292
R4100 VDDD.n1877 VDDD.n1876 0.120292
R4101 VDDD.n1878 VDDD.n1877 0.120292
R4102 VDDD.n1878 VDDD.n1844 0.120292
R4103 VDDD.n1843 VDDD.n1842 0.120292
R4104 VDDD.n1884 VDDD.n1842 0.120292
R4105 VDDD.n1981 VDDD.n1980 0.120292
R4106 VDDD.n1981 VDDD.n1967 0.120292
R4107 VDDD.n1967 VDDD.n1966 0.120292
R4108 VDDD.n1987 VDDD.n1966 0.120292
R4109 VDDD.n1988 VDDD.n1987 0.120292
R4110 VDDD.n1989 VDDD.n1988 0.120292
R4111 VDDD.n1989 VDDD.n1963 0.120292
R4112 VDDD.n1993 VDDD.n1963 0.120292
R4113 VDDD.n1994 VDDD.n1993 0.120292
R4114 VDDD.n1995 VDDD.n1994 0.120292
R4115 VDDD.n1995 VDDD.n1960 0.120292
R4116 VDDD.n2000 VDDD.n1960 0.120292
R4117 VDDD.n2001 VDDD.n2000 0.120292
R4118 VDDD.n2002 VDDD.n2001 0.120292
R4119 VDDD.n2002 VDDD.n1958 0.120292
R4120 VDDD.n2006 VDDD.n1958 0.120292
R4121 VDDD.n2007 VDDD.n2006 0.120292
R4122 VDDD.n2008 VDDD.n2007 0.120292
R4123 VDDD.n2008 VDDD.n1955 0.120292
R4124 VDDD.n2012 VDDD.n1955 0.120292
R4125 VDDD.n2014 VDDD.n2013 0.120292
R4126 VDDD.n2014 VDDD.n1953 0.120292
R4127 VDDD.n1953 VDDD.n1952 0.120292
R4128 VDDD.n2020 VDDD.n1952 0.120292
R4129 VDDD.n2021 VDDD.n2020 0.120292
R4130 VDDD.n2022 VDDD.n2021 0.120292
R4131 VDDD.n2022 VDDD.n1949 0.120292
R4132 VDDD.n2026 VDDD.n1949 0.120292
R4133 VDDD.n2027 VDDD.n2026 0.120292
R4134 VDDD.n2028 VDDD.n2027 0.120292
R4135 VDDD.n2028 VDDD.n1946 0.120292
R4136 VDDD.n2033 VDDD.n1946 0.120292
R4137 VDDD.n2034 VDDD.n2033 0.120292
R4138 VDDD.n2035 VDDD.n2034 0.120292
R4139 VDDD.n2035 VDDD.n1944 0.120292
R4140 VDDD.n2039 VDDD.n1944 0.120292
R4141 VDDD.n2040 VDDD.n2039 0.120292
R4142 VDDD.n2041 VDDD.n2040 0.120292
R4143 VDDD.n2041 VDDD.n1941 0.120292
R4144 VDDD.n2045 VDDD.n1941 0.120292
R4145 VDDD.n2047 VDDD.n2046 0.120292
R4146 VDDD.n2047 VDDD.n1939 0.120292
R4147 VDDD.n1939 VDDD.n1938 0.120292
R4148 VDDD.n2053 VDDD.n1938 0.120292
R4149 VDDD.n2054 VDDD.n2053 0.120292
R4150 VDDD.n2055 VDDD.n2054 0.120292
R4151 VDDD.n2055 VDDD.n1935 0.120292
R4152 VDDD.n2059 VDDD.n1935 0.120292
R4153 VDDD.n2060 VDDD.n2059 0.120292
R4154 VDDD.n2061 VDDD.n2060 0.120292
R4155 VDDD.n2061 VDDD.n1932 0.120292
R4156 VDDD.n2066 VDDD.n1932 0.120292
R4157 VDDD.n2067 VDDD.n2066 0.120292
R4158 VDDD.n2068 VDDD.n2067 0.120292
R4159 VDDD.n2068 VDDD.n1930 0.120292
R4160 VDDD.n2072 VDDD.n1930 0.120292
R4161 VDDD.n2073 VDDD.n2072 0.120292
R4162 VDDD.n2074 VDDD.n2073 0.120292
R4163 VDDD.n2074 VDDD.n1927 0.120292
R4164 VDDD.n2078 VDDD.n1927 0.120292
R4165 VDDD.n2080 VDDD.n2079 0.120292
R4166 VDDD.n2080 VDDD.n1925 0.120292
R4167 VDDD.n1925 VDDD.n1924 0.120292
R4168 VDDD.n2086 VDDD.n1924 0.120292
R4169 VDDD.n2087 VDDD.n2086 0.120292
R4170 VDDD.n2088 VDDD.n2087 0.120292
R4171 VDDD.n2088 VDDD.n1921 0.120292
R4172 VDDD.n2092 VDDD.n1921 0.120292
R4173 VDDD.n2093 VDDD.n2092 0.120292
R4174 VDDD.n2094 VDDD.n2093 0.120292
R4175 VDDD.n2094 VDDD.n1918 0.120292
R4176 VDDD.n2099 VDDD.n1918 0.120292
R4177 VDDD.n2100 VDDD.n2099 0.120292
R4178 VDDD.n2101 VDDD.n2100 0.120292
R4179 VDDD.n2101 VDDD.n1916 0.120292
R4180 VDDD.n2105 VDDD.n1916 0.120292
R4181 VDDD.n2106 VDDD.n2105 0.120292
R4182 VDDD.n2107 VDDD.n2106 0.120292
R4183 VDDD.n2107 VDDD.n1913 0.120292
R4184 VDDD.n2111 VDDD.n1913 0.120292
R4185 VDDD.n2113 VDDD.n2112 0.120292
R4186 VDDD.n2113 VDDD.n1911 0.120292
R4187 VDDD.n1911 VDDD.n1910 0.120292
R4188 VDDD.n2119 VDDD.n1910 0.120292
R4189 VDDD.n2120 VDDD.n2119 0.120292
R4190 VDDD.n2121 VDDD.n2120 0.120292
R4191 VDDD.n2121 VDDD.n1907 0.120292
R4192 VDDD.n2125 VDDD.n1907 0.120292
R4193 VDDD.n2126 VDDD.n2125 0.120292
R4194 VDDD.n2127 VDDD.n2126 0.120292
R4195 VDDD.n2127 VDDD.n1904 0.120292
R4196 VDDD.n2132 VDDD.n1904 0.120292
R4197 VDDD.n2133 VDDD.n2132 0.120292
R4198 VDDD.n2134 VDDD.n2133 0.120292
R4199 VDDD.n2134 VDDD.n1902 0.120292
R4200 VDDD.n2138 VDDD.n1902 0.120292
R4201 VDDD.n2139 VDDD.n2138 0.120292
R4202 VDDD.n2140 VDDD.n2139 0.120292
R4203 VDDD.n2140 VDDD.n1899 0.120292
R4204 VDDD.n2144 VDDD.n1899 0.120292
R4205 VDDD.n2146 VDDD.n2145 0.120292
R4206 VDDD.n2146 VDDD.n1897 0.120292
R4207 VDDD.n2150 VDDD.n1897 0.120292
R4208 VDDD.n2151 VDDD.n2150 0.120292
R4209 VDDD.n2151 VDDD.n1894 0.120292
R4210 VDDD.n2155 VDDD.n1894 0.120292
R4211 VDDD.n2156 VDDD.n2155 0.120292
R4212 VDDD.n2157 VDDD.n2156 0.120292
R4213 VDDD.n2157 VDDD.n1892 0.120292
R4214 VDDD.n1892 VDDD.n1891 0.120292
R4215 VDDD.n2164 VDDD.n1891 0.120292
R4216 VDDD.n2165 VDDD.n2164 0.120292
R4217 VDDD.n2166 VDDD.n2165 0.120292
R4218 VDDD.n2166 VDDD.n1889 0.120292
R4219 VDDD.n2170 VDDD.n1889 0.120292
R4220 VDDD.n2171 VDDD.n2170 0.120292
R4221 VDDD.n2172 VDDD.n2171 0.120292
R4222 VDDD.n2172 VDDD.n1886 0.120292
R4223 VDDD.n2277 VDDD.n2276 0.120292
R4224 VDDD.n2277 VDDD.n2259 0.120292
R4225 VDDD.n2259 VDDD.n2258 0.120292
R4226 VDDD.n2283 VDDD.n2258 0.120292
R4227 VDDD.n2284 VDDD.n2283 0.120292
R4228 VDDD.n2285 VDDD.n2284 0.120292
R4229 VDDD.n2285 VDDD.n2255 0.120292
R4230 VDDD.n2289 VDDD.n2255 0.120292
R4231 VDDD.n2290 VDDD.n2289 0.120292
R4232 VDDD.n2291 VDDD.n2290 0.120292
R4233 VDDD.n2291 VDDD.n2252 0.120292
R4234 VDDD.n2296 VDDD.n2252 0.120292
R4235 VDDD.n2297 VDDD.n2296 0.120292
R4236 VDDD.n2298 VDDD.n2297 0.120292
R4237 VDDD.n2298 VDDD.n2250 0.120292
R4238 VDDD.n2302 VDDD.n2250 0.120292
R4239 VDDD.n2303 VDDD.n2302 0.120292
R4240 VDDD.n2304 VDDD.n2303 0.120292
R4241 VDDD.n2304 VDDD.n2247 0.120292
R4242 VDDD.n2308 VDDD.n2247 0.120292
R4243 VDDD.n2310 VDDD.n2309 0.120292
R4244 VDDD.n2310 VDDD.n2245 0.120292
R4245 VDDD.n2245 VDDD.n2244 0.120292
R4246 VDDD.n2316 VDDD.n2244 0.120292
R4247 VDDD.n2317 VDDD.n2316 0.120292
R4248 VDDD.n2318 VDDD.n2317 0.120292
R4249 VDDD.n2318 VDDD.n2241 0.120292
R4250 VDDD.n2322 VDDD.n2241 0.120292
R4251 VDDD.n2323 VDDD.n2322 0.120292
R4252 VDDD.n2324 VDDD.n2323 0.120292
R4253 VDDD.n2324 VDDD.n2238 0.120292
R4254 VDDD.n2329 VDDD.n2238 0.120292
R4255 VDDD.n2330 VDDD.n2329 0.120292
R4256 VDDD.n2331 VDDD.n2330 0.120292
R4257 VDDD.n2331 VDDD.n2236 0.120292
R4258 VDDD.n2335 VDDD.n2236 0.120292
R4259 VDDD.n2336 VDDD.n2335 0.120292
R4260 VDDD.n2337 VDDD.n2336 0.120292
R4261 VDDD.n2337 VDDD.n2233 0.120292
R4262 VDDD.n2341 VDDD.n2233 0.120292
R4263 VDDD.n2343 VDDD.n2342 0.120292
R4264 VDDD.n2343 VDDD.n2231 0.120292
R4265 VDDD.n2231 VDDD.n2230 0.120292
R4266 VDDD.n2349 VDDD.n2230 0.120292
R4267 VDDD.n2350 VDDD.n2349 0.120292
R4268 VDDD.n2351 VDDD.n2350 0.120292
R4269 VDDD.n2351 VDDD.n2227 0.120292
R4270 VDDD.n2355 VDDD.n2227 0.120292
R4271 VDDD.n2356 VDDD.n2355 0.120292
R4272 VDDD.n2357 VDDD.n2356 0.120292
R4273 VDDD.n2357 VDDD.n2224 0.120292
R4274 VDDD.n2362 VDDD.n2224 0.120292
R4275 VDDD.n2363 VDDD.n2362 0.120292
R4276 VDDD.n2364 VDDD.n2363 0.120292
R4277 VDDD.n2364 VDDD.n2222 0.120292
R4278 VDDD.n2368 VDDD.n2222 0.120292
R4279 VDDD.n2369 VDDD.n2368 0.120292
R4280 VDDD.n2370 VDDD.n2369 0.120292
R4281 VDDD.n2370 VDDD.n2219 0.120292
R4282 VDDD.n2374 VDDD.n2219 0.120292
R4283 VDDD.n2376 VDDD.n2375 0.120292
R4284 VDDD.n2376 VDDD.n2217 0.120292
R4285 VDDD.n2217 VDDD.n2216 0.120292
R4286 VDDD.n2382 VDDD.n2216 0.120292
R4287 VDDD.n2383 VDDD.n2382 0.120292
R4288 VDDD.n2384 VDDD.n2383 0.120292
R4289 VDDD.n2384 VDDD.n2213 0.120292
R4290 VDDD.n2388 VDDD.n2213 0.120292
R4291 VDDD.n2389 VDDD.n2388 0.120292
R4292 VDDD.n2390 VDDD.n2389 0.120292
R4293 VDDD.n2390 VDDD.n2210 0.120292
R4294 VDDD.n2395 VDDD.n2210 0.120292
R4295 VDDD.n2396 VDDD.n2395 0.120292
R4296 VDDD.n2397 VDDD.n2396 0.120292
R4297 VDDD.n2397 VDDD.n2208 0.120292
R4298 VDDD.n2401 VDDD.n2208 0.120292
R4299 VDDD.n2402 VDDD.n2401 0.120292
R4300 VDDD.n2403 VDDD.n2402 0.120292
R4301 VDDD.n2403 VDDD.n2205 0.120292
R4302 VDDD.n2407 VDDD.n2205 0.120292
R4303 VDDD.n2409 VDDD.n2408 0.120292
R4304 VDDD.n2409 VDDD.n2203 0.120292
R4305 VDDD.n2203 VDDD.n2202 0.120292
R4306 VDDD.n2415 VDDD.n2202 0.120292
R4307 VDDD.n2416 VDDD.n2415 0.120292
R4308 VDDD.n2417 VDDD.n2416 0.120292
R4309 VDDD.n2417 VDDD.n2199 0.120292
R4310 VDDD.n2421 VDDD.n2199 0.120292
R4311 VDDD.n2422 VDDD.n2421 0.120292
R4312 VDDD.n2423 VDDD.n2422 0.120292
R4313 VDDD.n2423 VDDD.n2196 0.120292
R4314 VDDD.n2428 VDDD.n2196 0.120292
R4315 VDDD.n2429 VDDD.n2428 0.120292
R4316 VDDD.n2430 VDDD.n2429 0.120292
R4317 VDDD.n2430 VDDD.n2194 0.120292
R4318 VDDD.n2434 VDDD.n2194 0.120292
R4319 VDDD.n2435 VDDD.n2434 0.120292
R4320 VDDD.n2436 VDDD.n2435 0.120292
R4321 VDDD.n2436 VDDD.n2191 0.120292
R4322 VDDD.n2440 VDDD.n2191 0.120292
R4323 VDDD.n2442 VDDD.n2441 0.120292
R4324 VDDD.n2442 VDDD.n2189 0.120292
R4325 VDDD.n2446 VDDD.n2189 0.120292
R4326 VDDD.n2447 VDDD.n2446 0.120292
R4327 VDDD.n2447 VDDD.n2186 0.120292
R4328 VDDD.n2451 VDDD.n2186 0.120292
R4329 VDDD.n2452 VDDD.n2451 0.120292
R4330 VDDD.n2453 VDDD.n2452 0.120292
R4331 VDDD.n2453 VDDD.n2184 0.120292
R4332 VDDD.n2184 VDDD.n2183 0.120292
R4333 VDDD.n2460 VDDD.n2183 0.120292
R4334 VDDD.n2461 VDDD.n2460 0.120292
R4335 VDDD.n2462 VDDD.n2461 0.120292
R4336 VDDD.n2462 VDDD.n2181 0.120292
R4337 VDDD.n2466 VDDD.n2181 0.120292
R4338 VDDD.n2467 VDDD.n2466 0.120292
R4339 VDDD.n2468 VDDD.n2467 0.120292
R4340 VDDD.n2468 VDDD.n2178 0.120292
R4341 VDDD.n1668 VDDD.n1667 0.120292
R4342 VDDD.n1668 VDDD.n1374 0.120292
R4343 VDDD.n1374 VDDD.n1373 0.120292
R4344 VDDD.n1674 VDDD.n1373 0.120292
R4345 VDDD.n1675 VDDD.n1674 0.120292
R4346 VDDD.n1676 VDDD.n1675 0.120292
R4347 VDDD.n1676 VDDD.n1370 0.120292
R4348 VDDD.n1680 VDDD.n1370 0.120292
R4349 VDDD.n1681 VDDD.n1680 0.120292
R4350 VDDD.n1682 VDDD.n1681 0.120292
R4351 VDDD.n1682 VDDD.n1367 0.120292
R4352 VDDD.n1687 VDDD.n1367 0.120292
R4353 VDDD.n1688 VDDD.n1687 0.120292
R4354 VDDD.n1689 VDDD.n1688 0.120292
R4355 VDDD.n1689 VDDD.n1365 0.120292
R4356 VDDD.n1693 VDDD.n1365 0.120292
R4357 VDDD.n1694 VDDD.n1693 0.120292
R4358 VDDD.n1695 VDDD.n1694 0.120292
R4359 VDDD.n1695 VDDD.n1362 0.120292
R4360 VDDD.n1699 VDDD.n1362 0.120292
R4361 VDDD.n1701 VDDD.n1700 0.120292
R4362 VDDD.n1701 VDDD.n1360 0.120292
R4363 VDDD.n1360 VDDD.n1359 0.120292
R4364 VDDD.n1707 VDDD.n1359 0.120292
R4365 VDDD.n1708 VDDD.n1707 0.120292
R4366 VDDD.n1709 VDDD.n1708 0.120292
R4367 VDDD.n1709 VDDD.n1356 0.120292
R4368 VDDD.n1713 VDDD.n1356 0.120292
R4369 VDDD.n1714 VDDD.n1713 0.120292
R4370 VDDD.n1715 VDDD.n1714 0.120292
R4371 VDDD.n1715 VDDD.n1353 0.120292
R4372 VDDD.n1720 VDDD.n1353 0.120292
R4373 VDDD.n1721 VDDD.n1720 0.120292
R4374 VDDD.n1722 VDDD.n1721 0.120292
R4375 VDDD.n1722 VDDD.n1351 0.120292
R4376 VDDD.n1726 VDDD.n1351 0.120292
R4377 VDDD.n1727 VDDD.n1726 0.120292
R4378 VDDD.n1728 VDDD.n1727 0.120292
R4379 VDDD.n1728 VDDD.n1348 0.120292
R4380 VDDD.n1732 VDDD.n1348 0.120292
R4381 VDDD.n1734 VDDD.n1733 0.120292
R4382 VDDD.n1734 VDDD.n1346 0.120292
R4383 VDDD.n1346 VDDD.n1345 0.120292
R4384 VDDD.n1740 VDDD.n1345 0.120292
R4385 VDDD.n1741 VDDD.n1740 0.120292
R4386 VDDD.n1742 VDDD.n1741 0.120292
R4387 VDDD.n1742 VDDD.n1342 0.120292
R4388 VDDD.n1746 VDDD.n1342 0.120292
R4389 VDDD.n1747 VDDD.n1746 0.120292
R4390 VDDD.n1748 VDDD.n1747 0.120292
R4391 VDDD.n1748 VDDD.n1339 0.120292
R4392 VDDD.n1753 VDDD.n1339 0.120292
R4393 VDDD.n1754 VDDD.n1753 0.120292
R4394 VDDD.n1755 VDDD.n1754 0.120292
R4395 VDDD.n1755 VDDD.n1337 0.120292
R4396 VDDD.n1759 VDDD.n1337 0.120292
R4397 VDDD.n1760 VDDD.n1759 0.120292
R4398 VDDD.n1761 VDDD.n1760 0.120292
R4399 VDDD.n1761 VDDD.n1334 0.120292
R4400 VDDD.n1765 VDDD.n1334 0.120292
R4401 VDDD.n1767 VDDD.n1766 0.120292
R4402 VDDD.n1767 VDDD.n1332 0.120292
R4403 VDDD.n1332 VDDD.n1331 0.120292
R4404 VDDD.n1773 VDDD.n1331 0.120292
R4405 VDDD.n1774 VDDD.n1773 0.120292
R4406 VDDD.n1775 VDDD.n1774 0.120292
R4407 VDDD.n1775 VDDD.n1328 0.120292
R4408 VDDD.n1779 VDDD.n1328 0.120292
R4409 VDDD.n1780 VDDD.n1779 0.120292
R4410 VDDD.n1781 VDDD.n1780 0.120292
R4411 VDDD.n1781 VDDD.n1325 0.120292
R4412 VDDD.n1786 VDDD.n1325 0.120292
R4413 VDDD.n1787 VDDD.n1786 0.120292
R4414 VDDD.n1788 VDDD.n1787 0.120292
R4415 VDDD.n1788 VDDD.n1323 0.120292
R4416 VDDD.n1792 VDDD.n1323 0.120292
R4417 VDDD.n1793 VDDD.n1792 0.120292
R4418 VDDD.n1794 VDDD.n1793 0.120292
R4419 VDDD.n1794 VDDD.n1320 0.120292
R4420 VDDD.n1798 VDDD.n1320 0.120292
R4421 VDDD.n1800 VDDD.n1799 0.120292
R4422 VDDD.n1800 VDDD.n1318 0.120292
R4423 VDDD.n1804 VDDD.n1318 0.120292
R4424 VDDD.n1805 VDDD.n1804 0.120292
R4425 VDDD.n1805 VDDD.n1315 0.120292
R4426 VDDD.n1809 VDDD.n1315 0.120292
R4427 VDDD.n1810 VDDD.n1809 0.120292
R4428 VDDD.n1811 VDDD.n1810 0.120292
R4429 VDDD.n1811 VDDD.n1313 0.120292
R4430 VDDD.n1313 VDDD.n1312 0.120292
R4431 VDDD.n1818 VDDD.n1312 0.120292
R4432 VDDD.n1819 VDDD.n1818 0.120292
R4433 VDDD.n1820 VDDD.n1819 0.120292
R4434 VDDD.n1820 VDDD.n1310 0.120292
R4435 VDDD.n1824 VDDD.n1310 0.120292
R4436 VDDD.n1825 VDDD.n1824 0.120292
R4437 VDDD.n1826 VDDD.n1825 0.120292
R4438 VDDD.n1826 VDDD.n1307 0.120292
R4439 VDDD.n1637 VDDD.n1377 0.120292
R4440 VDDD.n1637 VDDD.n1636 0.120292
R4441 VDDD.n1636 VDDD.n1635 0.120292
R4442 VDDD.n1635 VDDD.n1379 0.120292
R4443 VDDD.n1631 VDDD.n1379 0.120292
R4444 VDDD.n1631 VDDD.n1630 0.120292
R4445 VDDD.n1630 VDDD.n1629 0.120292
R4446 VDDD.n1629 VDDD.n1381 0.120292
R4447 VDDD.n1624 VDDD.n1381 0.120292
R4448 VDDD.n1624 VDDD.n1623 0.120292
R4449 VDDD.n1623 VDDD.n1622 0.120292
R4450 VDDD.n1622 VDDD.n1384 0.120292
R4451 VDDD.n1618 VDDD.n1384 0.120292
R4452 VDDD.n1618 VDDD.n1617 0.120292
R4453 VDDD.n1617 VDDD.n1616 0.120292
R4454 VDDD.n1616 VDDD.n1387 0.120292
R4455 VDDD.n1388 VDDD.n1387 0.120292
R4456 VDDD.n1610 VDDD.n1388 0.120292
R4457 VDDD.n1610 VDDD.n1609 0.120292
R4458 VDDD.n1604 VDDD.n1391 0.120292
R4459 VDDD.n1604 VDDD.n1603 0.120292
R4460 VDDD.n1603 VDDD.n1602 0.120292
R4461 VDDD.n1602 VDDD.n1393 0.120292
R4462 VDDD.n1598 VDDD.n1393 0.120292
R4463 VDDD.n1598 VDDD.n1597 0.120292
R4464 VDDD.n1597 VDDD.n1596 0.120292
R4465 VDDD.n1596 VDDD.n1395 0.120292
R4466 VDDD.n1591 VDDD.n1395 0.120292
R4467 VDDD.n1591 VDDD.n1590 0.120292
R4468 VDDD.n1590 VDDD.n1589 0.120292
R4469 VDDD.n1589 VDDD.n1398 0.120292
R4470 VDDD.n1585 VDDD.n1398 0.120292
R4471 VDDD.n1585 VDDD.n1584 0.120292
R4472 VDDD.n1584 VDDD.n1583 0.120292
R4473 VDDD.n1583 VDDD.n1401 0.120292
R4474 VDDD.n1402 VDDD.n1401 0.120292
R4475 VDDD.n1577 VDDD.n1402 0.120292
R4476 VDDD.n1577 VDDD.n1576 0.120292
R4477 VDDD.n1571 VDDD.n1405 0.120292
R4478 VDDD.n1571 VDDD.n1570 0.120292
R4479 VDDD.n1570 VDDD.n1569 0.120292
R4480 VDDD.n1569 VDDD.n1407 0.120292
R4481 VDDD.n1565 VDDD.n1407 0.120292
R4482 VDDD.n1565 VDDD.n1564 0.120292
R4483 VDDD.n1564 VDDD.n1563 0.120292
R4484 VDDD.n1563 VDDD.n1409 0.120292
R4485 VDDD.n1558 VDDD.n1409 0.120292
R4486 VDDD.n1558 VDDD.n1557 0.120292
R4487 VDDD.n1557 VDDD.n1556 0.120292
R4488 VDDD.n1556 VDDD.n1412 0.120292
R4489 VDDD.n1552 VDDD.n1412 0.120292
R4490 VDDD.n1552 VDDD.n1551 0.120292
R4491 VDDD.n1551 VDDD.n1550 0.120292
R4492 VDDD.n1550 VDDD.n1415 0.120292
R4493 VDDD.n1416 VDDD.n1415 0.120292
R4494 VDDD.n1544 VDDD.n1416 0.120292
R4495 VDDD.n1544 VDDD.n1543 0.120292
R4496 VDDD.n1538 VDDD.n1419 0.120292
R4497 VDDD.n1538 VDDD.n1537 0.120292
R4498 VDDD.n1537 VDDD.n1536 0.120292
R4499 VDDD.n1536 VDDD.n1421 0.120292
R4500 VDDD.n1532 VDDD.n1421 0.120292
R4501 VDDD.n1532 VDDD.n1531 0.120292
R4502 VDDD.n1531 VDDD.n1530 0.120292
R4503 VDDD.n1530 VDDD.n1423 0.120292
R4504 VDDD.n1525 VDDD.n1423 0.120292
R4505 VDDD.n1525 VDDD.n1524 0.120292
R4506 VDDD.n1524 VDDD.n1523 0.120292
R4507 VDDD.n1523 VDDD.n1426 0.120292
R4508 VDDD.n1519 VDDD.n1426 0.120292
R4509 VDDD.n1519 VDDD.n1518 0.120292
R4510 VDDD.n1518 VDDD.n1517 0.120292
R4511 VDDD.n1517 VDDD.n1429 0.120292
R4512 VDDD.n1430 VDDD.n1429 0.120292
R4513 VDDD.n1511 VDDD.n1430 0.120292
R4514 VDDD.n1511 VDDD.n1510 0.120292
R4515 VDDD.n1505 VDDD.n1433 0.120292
R4516 VDDD.n1505 VDDD.n1504 0.120292
R4517 VDDD.n1504 VDDD.n1503 0.120292
R4518 VDDD.n1503 VDDD.n1435 0.120292
R4519 VDDD.n1499 VDDD.n1435 0.120292
R4520 VDDD.n1499 VDDD.n1498 0.120292
R4521 VDDD.n1498 VDDD.n1497 0.120292
R4522 VDDD.n1497 VDDD.n1437 0.120292
R4523 VDDD.n1492 VDDD.n1437 0.120292
R4524 VDDD.n1492 VDDD.n1491 0.120292
R4525 VDDD.n1491 VDDD.n1490 0.120292
R4526 VDDD.n1490 VDDD.n1440 0.120292
R4527 VDDD.n1486 VDDD.n1440 0.120292
R4528 VDDD.n1486 VDDD.n1485 0.120292
R4529 VDDD.n1485 VDDD.n1484 0.120292
R4530 VDDD.n1484 VDDD.n1443 0.120292
R4531 VDDD.n1444 VDDD.n1443 0.120292
R4532 VDDD.n1478 VDDD.n1444 0.120292
R4533 VDDD.n1478 VDDD.n1477 0.120292
R4534 VDDD.n1472 VDDD.n1471 0.120292
R4535 VDDD.n1471 VDDD.n1470 0.120292
R4536 VDDD.n1470 VDDD.n1448 0.120292
R4537 VDDD.n1465 VDDD.n1448 0.120292
R4538 VDDD.n1465 VDDD.n1464 0.120292
R4539 VDDD.n1464 VDDD.n1463 0.120292
R4540 VDDD.n1463 VDDD.n1453 0.120292
R4541 VDDD.n1459 VDDD.n1453 0.120292
R4542 VDDD.n1111 VDDD.n1091 0.120292
R4543 VDDD.n1112 VDDD.n1111 0.120292
R4544 VDDD.n1113 VDDD.n1112 0.120292
R4545 VDDD.n1118 VDDD.n1117 0.120292
R4546 VDDD.n1118 VDDD.n1087 0.120292
R4547 VDDD.n1124 VDDD.n1087 0.120292
R4548 VDDD.n1125 VDDD.n1124 0.120292
R4549 VDDD.n1126 VDDD.n1125 0.120292
R4550 VDDD.n1126 VDDD.n1084 0.120292
R4551 VDDD.n1130 VDDD.n1084 0.120292
R4552 VDDD.n1131 VDDD.n1130 0.120292
R4553 VDDD.n1131 VDDD.n1081 0.120292
R4554 VDDD.n1135 VDDD.n1081 0.120292
R4555 VDDD.n1136 VDDD.n1135 0.120292
R4556 VDDD.n1136 VDDD.n1078 0.120292
R4557 VDDD.n1140 VDDD.n1078 0.120292
R4558 VDDD.n1141 VDDD.n1140 0.120292
R4559 VDDD.n1142 VDDD.n1141 0.120292
R4560 VDDD.n1142 VDDD.n1075 0.120292
R4561 VDDD.n1148 VDDD.n1075 0.120292
R4562 VDDD.n1149 VDDD.n1148 0.120292
R4563 VDDD.n1150 VDDD.n1149 0.120292
R4564 VDDD.n1155 VDDD.n1154 0.120292
R4565 VDDD.n1155 VDDD.n1070 0.120292
R4566 VDDD.n1161 VDDD.n1070 0.120292
R4567 VDDD.n1162 VDDD.n1161 0.120292
R4568 VDDD.n1163 VDDD.n1162 0.120292
R4569 VDDD.n1163 VDDD.n1067 0.120292
R4570 VDDD.n1167 VDDD.n1067 0.120292
R4571 VDDD.n1168 VDDD.n1167 0.120292
R4572 VDDD.n1168 VDDD.n1064 0.120292
R4573 VDDD.n1172 VDDD.n1064 0.120292
R4574 VDDD.n1173 VDDD.n1172 0.120292
R4575 VDDD.n1173 VDDD.n1061 0.120292
R4576 VDDD.n1177 VDDD.n1061 0.120292
R4577 VDDD.n1178 VDDD.n1177 0.120292
R4578 VDDD.n1179 VDDD.n1178 0.120292
R4579 VDDD.n1179 VDDD.n1058 0.120292
R4580 VDDD.n1185 VDDD.n1058 0.120292
R4581 VDDD.n1186 VDDD.n1185 0.120292
R4582 VDDD.n1187 VDDD.n1186 0.120292
R4583 VDDD.n1192 VDDD.n1191 0.120292
R4584 VDDD.n1192 VDDD.n1053 0.120292
R4585 VDDD.n1198 VDDD.n1053 0.120292
R4586 VDDD.n1199 VDDD.n1198 0.120292
R4587 VDDD.n1200 VDDD.n1199 0.120292
R4588 VDDD.n1200 VDDD.n1050 0.120292
R4589 VDDD.n1204 VDDD.n1050 0.120292
R4590 VDDD.n1205 VDDD.n1204 0.120292
R4591 VDDD.n1205 VDDD.n1047 0.120292
R4592 VDDD.n1209 VDDD.n1047 0.120292
R4593 VDDD.n1210 VDDD.n1209 0.120292
R4594 VDDD.n1210 VDDD.n1044 0.120292
R4595 VDDD.n1214 VDDD.n1044 0.120292
R4596 VDDD.n1215 VDDD.n1214 0.120292
R4597 VDDD.n1216 VDDD.n1215 0.120292
R4598 VDDD.n1216 VDDD.n1041 0.120292
R4599 VDDD.n1222 VDDD.n1041 0.120292
R4600 VDDD.n1223 VDDD.n1222 0.120292
R4601 VDDD.n1224 VDDD.n1223 0.120292
R4602 VDDD.n1229 VDDD.n1228 0.120292
R4603 VDDD.n1229 VDDD.n1036 0.120292
R4604 VDDD.n1235 VDDD.n1036 0.120292
R4605 VDDD.n1236 VDDD.n1235 0.120292
R4606 VDDD.n1237 VDDD.n1236 0.120292
R4607 VDDD.n1237 VDDD.n1033 0.120292
R4608 VDDD.n1241 VDDD.n1033 0.120292
R4609 VDDD.n1242 VDDD.n1241 0.120292
R4610 VDDD.n1242 VDDD.n1030 0.120292
R4611 VDDD.n1246 VDDD.n1030 0.120292
R4612 VDDD.n1247 VDDD.n1246 0.120292
R4613 VDDD.n1247 VDDD.n1027 0.120292
R4614 VDDD.n1251 VDDD.n1027 0.120292
R4615 VDDD.n1252 VDDD.n1251 0.120292
R4616 VDDD.n1253 VDDD.n1252 0.120292
R4617 VDDD.n1253 VDDD.n1024 0.120292
R4618 VDDD.n1259 VDDD.n1024 0.120292
R4619 VDDD.n1260 VDDD.n1259 0.120292
R4620 VDDD.n1261 VDDD.n1260 0.120292
R4621 VDDD.n1266 VDDD.n1265 0.120292
R4622 VDDD.n1266 VDDD.n1019 0.120292
R4623 VDDD.n1272 VDDD.n1019 0.120292
R4624 VDDD.n1273 VDDD.n1272 0.120292
R4625 VDDD.n1274 VDDD.n1273 0.120292
R4626 VDDD.n1274 VDDD.n1016 0.120292
R4627 VDDD.n1280 VDDD.n1016 0.120292
R4628 VDDD.n1281 VDDD.n1280 0.120292
R4629 VDDD.n1282 VDDD.n1281 0.120292
R4630 VDDD.n1282 VDDD.n1014 0.120292
R4631 VDDD.n1288 VDDD.n1014 0.120292
R4632 VDDD.n1289 VDDD.n1288 0.120292
R4633 VDDD.n1290 VDDD.n1289 0.120292
R4634 VDDD.n1290 VDDD.n1012 0.120292
R4635 VDDD.n1297 VDDD.n1012 0.120292
R4636 VDDD.n1298 VDDD.n1297 0.120292
R4637 VDDD.n1299 VDDD.n1298 0.120292
R4638 VDDD.n1299 VDDD.n1009 0.120292
R4639 VDDD.n1303 VDDD.n1009 0.120292
R4640 VDDD.n639 VDDD.n638 0.120292
R4641 VDDD.n640 VDDD.n639 0.120292
R4642 VDDD.n640 VDDD.n133 0.120292
R4643 VDDD.n645 VDDD.n133 0.120292
R4644 VDDD.n646 VDDD.n645 0.120292
R4645 VDDD.n647 VDDD.n646 0.120292
R4646 VDDD.n647 VDDD.n130 0.120292
R4647 VDDD.n651 VDDD.n130 0.120292
R4648 VDDD.n652 VDDD.n651 0.120292
R4649 VDDD.n653 VDDD.n652 0.120292
R4650 VDDD.n653 VDDD.n128 0.120292
R4651 VDDD.n659 VDDD.n128 0.120292
R4652 VDDD.n660 VDDD.n659 0.120292
R4653 VDDD.n661 VDDD.n660 0.120292
R4654 VDDD.n661 VDDD.n126 0.120292
R4655 VDDD.n665 VDDD.n126 0.120292
R4656 VDDD.n666 VDDD.n665 0.120292
R4657 VDDD.n667 VDDD.n666 0.120292
R4658 VDDD.n667 VDDD.n124 0.120292
R4659 VDDD.n672 VDDD.n124 0.120292
R4660 VDDD.n674 VDDD.n673 0.120292
R4661 VDDD.n674 VDDD.n122 0.120292
R4662 VDDD.n679 VDDD.n122 0.120292
R4663 VDDD.n680 VDDD.n679 0.120292
R4664 VDDD.n681 VDDD.n680 0.120292
R4665 VDDD.n681 VDDD.n119 0.120292
R4666 VDDD.n685 VDDD.n119 0.120292
R4667 VDDD.n686 VDDD.n685 0.120292
R4668 VDDD.n687 VDDD.n686 0.120292
R4669 VDDD.n687 VDDD.n117 0.120292
R4670 VDDD.n691 VDDD.n117 0.120292
R4671 VDDD.n692 VDDD.n691 0.120292
R4672 VDDD.n692 VDDD.n114 0.120292
R4673 VDDD.n696 VDDD.n114 0.120292
R4674 VDDD.n697 VDDD.n696 0.120292
R4675 VDDD.n698 VDDD.n697 0.120292
R4676 VDDD.n698 VDDD.n112 0.120292
R4677 VDDD.n702 VDDD.n112 0.120292
R4678 VDDD.n703 VDDD.n702 0.120292
R4679 VDDD.n704 VDDD.n703 0.120292
R4680 VDDD.n708 VDDD.n707 0.120292
R4681 VDDD.n709 VDDD.n708 0.120292
R4682 VDDD.n709 VDDD.n108 0.120292
R4683 VDDD.n714 VDDD.n108 0.120292
R4684 VDDD.n715 VDDD.n714 0.120292
R4685 VDDD.n716 VDDD.n715 0.120292
R4686 VDDD.n716 VDDD.n105 0.120292
R4687 VDDD.n720 VDDD.n105 0.120292
R4688 VDDD.n721 VDDD.n720 0.120292
R4689 VDDD.n722 VDDD.n721 0.120292
R4690 VDDD.n722 VDDD.n103 0.120292
R4691 VDDD.n728 VDDD.n103 0.120292
R4692 VDDD.n729 VDDD.n728 0.120292
R4693 VDDD.n730 VDDD.n729 0.120292
R4694 VDDD.n730 VDDD.n101 0.120292
R4695 VDDD.n734 VDDD.n101 0.120292
R4696 VDDD.n735 VDDD.n734 0.120292
R4697 VDDD.n736 VDDD.n735 0.120292
R4698 VDDD.n736 VDDD.n99 0.120292
R4699 VDDD.n741 VDDD.n99 0.120292
R4700 VDDD.n743 VDDD.n742 0.120292
R4701 VDDD.n743 VDDD.n97 0.120292
R4702 VDDD.n748 VDDD.n97 0.120292
R4703 VDDD.n749 VDDD.n748 0.120292
R4704 VDDD.n750 VDDD.n749 0.120292
R4705 VDDD.n750 VDDD.n94 0.120292
R4706 VDDD.n754 VDDD.n94 0.120292
R4707 VDDD.n755 VDDD.n754 0.120292
R4708 VDDD.n756 VDDD.n755 0.120292
R4709 VDDD.n756 VDDD.n92 0.120292
R4710 VDDD.n760 VDDD.n92 0.120292
R4711 VDDD.n761 VDDD.n760 0.120292
R4712 VDDD.n761 VDDD.n89 0.120292
R4713 VDDD.n765 VDDD.n89 0.120292
R4714 VDDD.n766 VDDD.n765 0.120292
R4715 VDDD.n767 VDDD.n766 0.120292
R4716 VDDD.n767 VDDD.n87 0.120292
R4717 VDDD.n771 VDDD.n87 0.120292
R4718 VDDD.n772 VDDD.n771 0.120292
R4719 VDDD.n773 VDDD.n772 0.120292
R4720 VDDD.n777 VDDD.n776 0.120292
R4721 VDDD.n778 VDDD.n777 0.120292
R4722 VDDD.n778 VDDD.n83 0.120292
R4723 VDDD.n783 VDDD.n83 0.120292
R4724 VDDD.n784 VDDD.n783 0.120292
R4725 VDDD.n785 VDDD.n784 0.120292
R4726 VDDD.n785 VDDD.n80 0.120292
R4727 VDDD.n789 VDDD.n80 0.120292
R4728 VDDD.n790 VDDD.n789 0.120292
R4729 VDDD.n791 VDDD.n790 0.120292
R4730 VDDD.n791 VDDD.n78 0.120292
R4731 VDDD.n797 VDDD.n78 0.120292
R4732 VDDD.n798 VDDD.n797 0.120292
R4733 VDDD.n799 VDDD.n798 0.120292
R4734 VDDD.n799 VDDD.n76 0.120292
R4735 VDDD.n803 VDDD.n76 0.120292
R4736 VDDD.n804 VDDD.n803 0.120292
R4737 VDDD.n805 VDDD.n804 0.120292
R4738 VDDD.n805 VDDD.n74 0.120292
R4739 VDDD.n810 VDDD.n74 0.120292
R4740 VDDD.n812 VDDD.n811 0.120292
R4741 VDDD.n812 VDDD.n72 0.120292
R4742 VDDD.n817 VDDD.n72 0.120292
R4743 VDDD.n818 VDDD.n817 0.120292
R4744 VDDD.n819 VDDD.n818 0.120292
R4745 VDDD.n819 VDDD.n69 0.120292
R4746 VDDD.n823 VDDD.n69 0.120292
R4747 VDDD.n824 VDDD.n823 0.120292
R4748 VDDD.n825 VDDD.n824 0.120292
R4749 VDDD.n825 VDDD.n67 0.120292
R4750 VDDD.n829 VDDD.n67 0.120292
R4751 VDDD.n830 VDDD.n829 0.120292
R4752 VDDD.n830 VDDD.n64 0.120292
R4753 VDDD.n834 VDDD.n64 0.120292
R4754 VDDD.n835 VDDD.n834 0.120292
R4755 VDDD.n836 VDDD.n835 0.120292
R4756 VDDD.n836 VDDD.n62 0.120292
R4757 VDDD.n840 VDDD.n62 0.120292
R4758 VDDD.n841 VDDD.n840 0.120292
R4759 VDDD.n842 VDDD.n841 0.120292
R4760 VDDD.n846 VDDD.n845 0.120292
R4761 VDDD.n847 VDDD.n846 0.120292
R4762 VDDD.n847 VDDD.n58 0.120292
R4763 VDDD.n852 VDDD.n58 0.120292
R4764 VDDD.n853 VDDD.n852 0.120292
R4765 VDDD.n854 VDDD.n853 0.120292
R4766 VDDD.n854 VDDD.n55 0.120292
R4767 VDDD.n858 VDDD.n55 0.120292
R4768 VDDD.n859 VDDD.n858 0.120292
R4769 VDDD.n860 VDDD.n859 0.120292
R4770 VDDD.n860 VDDD.n53 0.120292
R4771 VDDD.n866 VDDD.n53 0.120292
R4772 VDDD.n867 VDDD.n866 0.120292
R4773 VDDD.n868 VDDD.n867 0.120292
R4774 VDDD.n868 VDDD.n51 0.120292
R4775 VDDD.n872 VDDD.n51 0.120292
R4776 VDDD.n873 VDDD.n872 0.120292
R4777 VDDD.n874 VDDD.n873 0.120292
R4778 VDDD.n874 VDDD.n49 0.120292
R4779 VDDD.n879 VDDD.n49 0.120292
R4780 VDDD.n881 VDDD.n880 0.120292
R4781 VDDD.n881 VDDD.n47 0.120292
R4782 VDDD.n886 VDDD.n47 0.120292
R4783 VDDD.n887 VDDD.n886 0.120292
R4784 VDDD.n888 VDDD.n887 0.120292
R4785 VDDD.n888 VDDD.n44 0.120292
R4786 VDDD.n892 VDDD.n44 0.120292
R4787 VDDD.n893 VDDD.n892 0.120292
R4788 VDDD.n894 VDDD.n893 0.120292
R4789 VDDD.n894 VDDD.n42 0.120292
R4790 VDDD.n898 VDDD.n42 0.120292
R4791 VDDD.n899 VDDD.n898 0.120292
R4792 VDDD.n899 VDDD.n39 0.120292
R4793 VDDD.n903 VDDD.n39 0.120292
R4794 VDDD.n904 VDDD.n903 0.120292
R4795 VDDD.n905 VDDD.n904 0.120292
R4796 VDDD.n905 VDDD.n37 0.120292
R4797 VDDD.n909 VDDD.n37 0.120292
R4798 VDDD.n910 VDDD.n909 0.120292
R4799 VDDD.n911 VDDD.n910 0.120292
R4800 VDDD.n915 VDDD.n914 0.120292
R4801 VDDD.n916 VDDD.n915 0.120292
R4802 VDDD.n916 VDDD.n33 0.120292
R4803 VDDD.n921 VDDD.n33 0.120292
R4804 VDDD.n922 VDDD.n921 0.120292
R4805 VDDD.n923 VDDD.n922 0.120292
R4806 VDDD.n923 VDDD.n30 0.120292
R4807 VDDD.n927 VDDD.n30 0.120292
R4808 VDDD.n928 VDDD.n927 0.120292
R4809 VDDD.n929 VDDD.n928 0.120292
R4810 VDDD.n929 VDDD.n28 0.120292
R4811 VDDD.n935 VDDD.n28 0.120292
R4812 VDDD.n936 VDDD.n935 0.120292
R4813 VDDD.n937 VDDD.n936 0.120292
R4814 VDDD.n937 VDDD.n26 0.120292
R4815 VDDD.n941 VDDD.n26 0.120292
R4816 VDDD.n942 VDDD.n941 0.120292
R4817 VDDD.n943 VDDD.n942 0.120292
R4818 VDDD.n943 VDDD.n24 0.120292
R4819 VDDD.n948 VDDD.n24 0.120292
R4820 VDDD.n950 VDDD.n949 0.120292
R4821 VDDD.n950 VDDD.n22 0.120292
R4822 VDDD.n955 VDDD.n22 0.120292
R4823 VDDD.n956 VDDD.n955 0.120292
R4824 VDDD.n957 VDDD.n956 0.120292
R4825 VDDD.n957 VDDD.n19 0.120292
R4826 VDDD.n961 VDDD.n19 0.120292
R4827 VDDD.n962 VDDD.n961 0.120292
R4828 VDDD.n963 VDDD.n962 0.120292
R4829 VDDD.n963 VDDD.n17 0.120292
R4830 VDDD.n967 VDDD.n17 0.120292
R4831 VDDD.n968 VDDD.n967 0.120292
R4832 VDDD.n968 VDDD.n14 0.120292
R4833 VDDD.n972 VDDD.n14 0.120292
R4834 VDDD.n973 VDDD.n972 0.120292
R4835 VDDD.n974 VDDD.n973 0.120292
R4836 VDDD.n974 VDDD.n12 0.120292
R4837 VDDD.n978 VDDD.n12 0.120292
R4838 VDDD.n979 VDDD.n978 0.120292
R4839 VDDD.n980 VDDD.n979 0.120292
R4840 VDDD.n984 VDDD.n983 0.120292
R4841 VDDD.n985 VDDD.n984 0.120292
R4842 VDDD.n985 VDDD.n8 0.120292
R4843 VDDD.n992 VDDD.n8 0.120292
R4844 VDDD.n993 VDDD.n992 0.120292
R4845 VDDD.n994 VDDD.n993 0.120292
R4846 VDDD.n994 VDDD.n6 0.120292
R4847 VDDD.n1000 VDDD.n6 0.120292
R4848 VDDD.n1001 VDDD.n1000 0.120292
R4849 VDDD.n1001 VDDD.n2 0.120292
R4850 VDDD.n1005 VDDD.n2 0.120292
R4851 VDDD.n636 VDDD.n135 0.120292
R4852 VDDD.n632 VDDD.n135 0.120292
R4853 VDDD.n632 VDDD.n631 0.120292
R4854 VDDD.n631 VDDD.n630 0.120292
R4855 VDDD.n630 VDDD.n137 0.120292
R4856 VDDD.n625 VDDD.n137 0.120292
R4857 VDDD.n625 VDDD.n624 0.120292
R4858 VDDD.n624 VDDD.n623 0.120292
R4859 VDDD.n623 VDDD.n140 0.120292
R4860 VDDD.n619 VDDD.n140 0.120292
R4861 VDDD.n619 VDDD.n618 0.120292
R4862 VDDD.n618 VDDD.n617 0.120292
R4863 VDDD.n617 VDDD.n142 0.120292
R4864 VDDD.n613 VDDD.n142 0.120292
R4865 VDDD.n613 VDDD.n612 0.120292
R4866 VDDD.n612 VDDD.n611 0.120292
R4867 VDDD.n611 VDDD.n146 0.120292
R4868 VDDD.n607 VDDD.n146 0.120292
R4869 VDDD.n607 VDDD.n606 0.120292
R4870 VDDD.n606 VDDD.n605 0.120292
R4871 VDDD.n602 VDDD.n601 0.120292
R4872 VDDD.n601 VDDD.n600 0.120292
R4873 VDDD.n600 VDDD.n150 0.120292
R4874 VDDD.n595 VDDD.n150 0.120292
R4875 VDDD.n595 VDDD.n594 0.120292
R4876 VDDD.n594 VDDD.n593 0.120292
R4877 VDDD.n593 VDDD.n153 0.120292
R4878 VDDD.n589 VDDD.n153 0.120292
R4879 VDDD.n589 VDDD.n588 0.120292
R4880 VDDD.n588 VDDD.n587 0.120292
R4881 VDDD.n587 VDDD.n155 0.120292
R4882 VDDD.n581 VDDD.n155 0.120292
R4883 VDDD.n581 VDDD.n580 0.120292
R4884 VDDD.n580 VDDD.n579 0.120292
R4885 VDDD.n579 VDDD.n157 0.120292
R4886 VDDD.n575 VDDD.n157 0.120292
R4887 VDDD.n575 VDDD.n574 0.120292
R4888 VDDD.n574 VDDD.n573 0.120292
R4889 VDDD.n573 VDDD.n159 0.120292
R4890 VDDD.n568 VDDD.n159 0.120292
R4891 VDDD.n567 VDDD.n566 0.120292
R4892 VDDD.n566 VDDD.n161 0.120292
R4893 VDDD.n562 VDDD.n161 0.120292
R4894 VDDD.n562 VDDD.n561 0.120292
R4895 VDDD.n561 VDDD.n163 0.120292
R4896 VDDD.n556 VDDD.n163 0.120292
R4897 VDDD.n556 VDDD.n555 0.120292
R4898 VDDD.n555 VDDD.n554 0.120292
R4899 VDDD.n554 VDDD.n165 0.120292
R4900 VDDD.n550 VDDD.n165 0.120292
R4901 VDDD.n550 VDDD.n549 0.120292
R4902 VDDD.n549 VDDD.n548 0.120292
R4903 VDDD.n548 VDDD.n167 0.120292
R4904 VDDD.n544 VDDD.n167 0.120292
R4905 VDDD.n544 VDDD.n543 0.120292
R4906 VDDD.n543 VDDD.n542 0.120292
R4907 VDDD.n542 VDDD.n171 0.120292
R4908 VDDD.n538 VDDD.n171 0.120292
R4909 VDDD.n538 VDDD.n537 0.120292
R4910 VDDD.n537 VDDD.n536 0.120292
R4911 VDDD.n533 VDDD.n532 0.120292
R4912 VDDD.n532 VDDD.n531 0.120292
R4913 VDDD.n531 VDDD.n175 0.120292
R4914 VDDD.n526 VDDD.n175 0.120292
R4915 VDDD.n526 VDDD.n525 0.120292
R4916 VDDD.n525 VDDD.n524 0.120292
R4917 VDDD.n524 VDDD.n178 0.120292
R4918 VDDD.n520 VDDD.n178 0.120292
R4919 VDDD.n520 VDDD.n519 0.120292
R4920 VDDD.n519 VDDD.n518 0.120292
R4921 VDDD.n518 VDDD.n180 0.120292
R4922 VDDD.n512 VDDD.n180 0.120292
R4923 VDDD.n512 VDDD.n511 0.120292
R4924 VDDD.n511 VDDD.n510 0.120292
R4925 VDDD.n510 VDDD.n182 0.120292
R4926 VDDD.n506 VDDD.n182 0.120292
R4927 VDDD.n506 VDDD.n505 0.120292
R4928 VDDD.n505 VDDD.n504 0.120292
R4929 VDDD.n504 VDDD.n184 0.120292
R4930 VDDD.n499 VDDD.n184 0.120292
R4931 VDDD.n498 VDDD.n497 0.120292
R4932 VDDD.n497 VDDD.n186 0.120292
R4933 VDDD.n493 VDDD.n186 0.120292
R4934 VDDD.n493 VDDD.n492 0.120292
R4935 VDDD.n492 VDDD.n188 0.120292
R4936 VDDD.n487 VDDD.n188 0.120292
R4937 VDDD.n487 VDDD.n486 0.120292
R4938 VDDD.n486 VDDD.n485 0.120292
R4939 VDDD.n485 VDDD.n190 0.120292
R4940 VDDD.n481 VDDD.n190 0.120292
R4941 VDDD.n481 VDDD.n480 0.120292
R4942 VDDD.n480 VDDD.n479 0.120292
R4943 VDDD.n479 VDDD.n192 0.120292
R4944 VDDD.n475 VDDD.n192 0.120292
R4945 VDDD.n475 VDDD.n474 0.120292
R4946 VDDD.n474 VDDD.n473 0.120292
R4947 VDDD.n473 VDDD.n196 0.120292
R4948 VDDD.n469 VDDD.n196 0.120292
R4949 VDDD.n469 VDDD.n468 0.120292
R4950 VDDD.n468 VDDD.n467 0.120292
R4951 VDDD.n464 VDDD.n463 0.120292
R4952 VDDD.n463 VDDD.n462 0.120292
R4953 VDDD.n462 VDDD.n200 0.120292
R4954 VDDD.n457 VDDD.n200 0.120292
R4955 VDDD.n457 VDDD.n456 0.120292
R4956 VDDD.n456 VDDD.n455 0.120292
R4957 VDDD.n455 VDDD.n203 0.120292
R4958 VDDD.n451 VDDD.n203 0.120292
R4959 VDDD.n451 VDDD.n450 0.120292
R4960 VDDD.n450 VDDD.n449 0.120292
R4961 VDDD.n449 VDDD.n205 0.120292
R4962 VDDD.n443 VDDD.n205 0.120292
R4963 VDDD.n443 VDDD.n442 0.120292
R4964 VDDD.n442 VDDD.n441 0.120292
R4965 VDDD.n441 VDDD.n207 0.120292
R4966 VDDD.n437 VDDD.n207 0.120292
R4967 VDDD.n437 VDDD.n436 0.120292
R4968 VDDD.n436 VDDD.n435 0.120292
R4969 VDDD.n435 VDDD.n209 0.120292
R4970 VDDD.n430 VDDD.n209 0.120292
R4971 VDDD.n429 VDDD.n428 0.120292
R4972 VDDD.n428 VDDD.n211 0.120292
R4973 VDDD.n424 VDDD.n211 0.120292
R4974 VDDD.n424 VDDD.n423 0.120292
R4975 VDDD.n423 VDDD.n213 0.120292
R4976 VDDD.n418 VDDD.n213 0.120292
R4977 VDDD.n418 VDDD.n417 0.120292
R4978 VDDD.n417 VDDD.n416 0.120292
R4979 VDDD.n416 VDDD.n215 0.120292
R4980 VDDD.n412 VDDD.n215 0.120292
R4981 VDDD.n412 VDDD.n411 0.120292
R4982 VDDD.n411 VDDD.n410 0.120292
R4983 VDDD.n410 VDDD.n217 0.120292
R4984 VDDD.n406 VDDD.n217 0.120292
R4985 VDDD.n406 VDDD.n405 0.120292
R4986 VDDD.n405 VDDD.n404 0.120292
R4987 VDDD.n404 VDDD.n221 0.120292
R4988 VDDD.n400 VDDD.n221 0.120292
R4989 VDDD.n400 VDDD.n399 0.120292
R4990 VDDD.n399 VDDD.n398 0.120292
R4991 VDDD.n395 VDDD.n394 0.120292
R4992 VDDD.n394 VDDD.n393 0.120292
R4993 VDDD.n393 VDDD.n225 0.120292
R4994 VDDD.n388 VDDD.n225 0.120292
R4995 VDDD.n388 VDDD.n387 0.120292
R4996 VDDD.n387 VDDD.n386 0.120292
R4997 VDDD.n386 VDDD.n228 0.120292
R4998 VDDD.n382 VDDD.n228 0.120292
R4999 VDDD.n382 VDDD.n381 0.120292
R5000 VDDD.n381 VDDD.n380 0.120292
R5001 VDDD.n380 VDDD.n230 0.120292
R5002 VDDD.n374 VDDD.n230 0.120292
R5003 VDDD.n374 VDDD.n373 0.120292
R5004 VDDD.n373 VDDD.n372 0.120292
R5005 VDDD.n372 VDDD.n232 0.120292
R5006 VDDD.n368 VDDD.n232 0.120292
R5007 VDDD.n368 VDDD.n367 0.120292
R5008 VDDD.n367 VDDD.n366 0.120292
R5009 VDDD.n366 VDDD.n234 0.120292
R5010 VDDD.n361 VDDD.n234 0.120292
R5011 VDDD.n360 VDDD.n359 0.120292
R5012 VDDD.n359 VDDD.n236 0.120292
R5013 VDDD.n355 VDDD.n236 0.120292
R5014 VDDD.n355 VDDD.n354 0.120292
R5015 VDDD.n354 VDDD.n238 0.120292
R5016 VDDD.n349 VDDD.n238 0.120292
R5017 VDDD.n349 VDDD.n348 0.120292
R5018 VDDD.n348 VDDD.n347 0.120292
R5019 VDDD.n347 VDDD.n240 0.120292
R5020 VDDD.n343 VDDD.n240 0.120292
R5021 VDDD.n343 VDDD.n342 0.120292
R5022 VDDD.n342 VDDD.n341 0.120292
R5023 VDDD.n341 VDDD.n242 0.120292
R5024 VDDD.n337 VDDD.n242 0.120292
R5025 VDDD.n337 VDDD.n336 0.120292
R5026 VDDD.n336 VDDD.n335 0.120292
R5027 VDDD.n335 VDDD.n246 0.120292
R5028 VDDD.n331 VDDD.n246 0.120292
R5029 VDDD.n331 VDDD.n330 0.120292
R5030 VDDD.n330 VDDD.n329 0.120292
R5031 VDDD.n326 VDDD.n325 0.120292
R5032 VDDD.n325 VDDD.n324 0.120292
R5033 VDDD.n324 VDDD.n250 0.120292
R5034 VDDD.n319 VDDD.n250 0.120292
R5035 VDDD.n319 VDDD.n318 0.120292
R5036 VDDD.n318 VDDD.n317 0.120292
R5037 VDDD.n317 VDDD.n253 0.120292
R5038 VDDD.n313 VDDD.n253 0.120292
R5039 VDDD.n313 VDDD.n312 0.120292
R5040 VDDD.n312 VDDD.n311 0.120292
R5041 VDDD.n311 VDDD.n255 0.120292
R5042 VDDD.n305 VDDD.n255 0.120292
R5043 VDDD.n305 VDDD.n304 0.120292
R5044 VDDD.n304 VDDD.n303 0.120292
R5045 VDDD.n303 VDDD.n257 0.120292
R5046 VDDD.n299 VDDD.n257 0.120292
R5047 VDDD.n299 VDDD.n298 0.120292
R5048 VDDD.n298 VDDD.n297 0.120292
R5049 VDDD.n297 VDDD.n259 0.120292
R5050 VDDD.n292 VDDD.n259 0.120292
R5051 VDDD.n291 VDDD.n290 0.120292
R5052 VDDD.n290 VDDD.n261 0.120292
R5053 VDDD.n285 VDDD.n261 0.120292
R5054 VDDD.n285 VDDD.n284 0.120292
R5055 VDDD.n284 VDDD.n283 0.120292
R5056 VDDD.n283 VDDD.n263 0.120292
R5057 VDDD.n277 VDDD.n263 0.120292
R5058 VDDD.n277 VDDD.n276 0.120292
R5059 VDDD.n276 VDDD.n275 0.120292
R5060 VDDD.n275 VDDD.n267 0.120292
R5061 VDDD.n271 VDDD.n267 0.120292
R5062 VDDD VDDD.n2176 0.114842
R5063 VDDD VDDD.n2472 0.114842
R5064 VDDD VDDD.n1830 0.114842
R5065 VDDD.n1377 VDDD 0.0981562
R5066 VDDD.n1391 VDDD 0.0981562
R5067 VDDD.n1405 VDDD 0.0981562
R5068 VDDD.n1419 VDDD 0.0981562
R5069 VDDD.n1433 VDDD 0.0981562
R5070 VDDD VDDD.n1091 0.0981562
R5071 VDDD.n1117 VDDD 0.0981562
R5072 VDDD.n1154 VDDD 0.0981562
R5073 VDDD.n1191 VDDD 0.0981562
R5074 VDDD.n1228 VDDD 0.0981562
R5075 VDDD.n1265 VDDD 0.0981562
R5076 VDDD.n1653 VDDD.n1641 0.0979026
R5077 VDDD.n1472 VDDD 0.0968542
R5078 VDDD.n1666 VDDD.n1654 0.0966538
R5079 VDDD.n1856 VDDD 0.0603958
R5080 VDDD VDDD.n1847 0.0603958
R5081 VDDD VDDD.n1843 0.0603958
R5082 VDDD.n2013 VDDD 0.0603958
R5083 VDDD.n2046 VDDD 0.0603958
R5084 VDDD.n2079 VDDD 0.0603958
R5085 VDDD.n2112 VDDD 0.0603958
R5086 VDDD.n2145 VDDD 0.0603958
R5087 VDDD.n2276 VDDD 0.0603958
R5088 VDDD.n2309 VDDD 0.0603958
R5089 VDDD.n2342 VDDD 0.0603958
R5090 VDDD.n2375 VDDD 0.0603958
R5091 VDDD.n2408 VDDD 0.0603958
R5092 VDDD.n2441 VDDD 0.0603958
R5093 VDDD.n1700 VDDD 0.0603958
R5094 VDDD.n1733 VDDD 0.0603958
R5095 VDDD.n1766 VDDD 0.0603958
R5096 VDDD.n1799 VDDD 0.0603958
R5097 VDDD.n1609 VDDD 0.0603958
R5098 VDDD VDDD.n1608 0.0603958
R5099 VDDD.n1576 VDDD 0.0603958
R5100 VDDD VDDD.n1575 0.0603958
R5101 VDDD.n1543 VDDD 0.0603958
R5102 VDDD VDDD.n1542 0.0603958
R5103 VDDD.n1510 VDDD 0.0603958
R5104 VDDD VDDD.n1509 0.0603958
R5105 VDDD.n1477 VDDD 0.0603958
R5106 VDDD.n1113 VDDD 0.0603958
R5107 VDDD.n1153 VDDD 0.0603958
R5108 VDDD.n1190 VDDD 0.0603958
R5109 VDDD.n1227 VDDD 0.0603958
R5110 VDDD.n1264 VDDD 0.0603958
R5111 VDDD.n673 VDDD 0.0603958
R5112 VDDD.n707 VDDD 0.0603958
R5113 VDDD.n742 VDDD 0.0603958
R5114 VDDD.n776 VDDD 0.0603958
R5115 VDDD.n811 VDDD 0.0603958
R5116 VDDD.n845 VDDD 0.0603958
R5117 VDDD.n880 VDDD 0.0603958
R5118 VDDD.n914 VDDD 0.0603958
R5119 VDDD.n949 VDDD 0.0603958
R5120 VDDD.n983 VDDD 0.0603958
R5121 VDDD.n602 VDDD 0.0603958
R5122 VDDD VDDD.n567 0.0603958
R5123 VDDD.n533 VDDD 0.0603958
R5124 VDDD VDDD.n498 0.0603958
R5125 VDDD.n464 VDDD 0.0603958
R5126 VDDD VDDD.n429 0.0603958
R5127 VDDD.n395 VDDD 0.0603958
R5128 VDDD VDDD.n360 0.0603958
R5129 VDDD.n326 VDDD 0.0603958
R5130 VDDD VDDD.n291 0.0603958
R5131 VDDD VDDD.n1476 0.0590938
R5132 VDDD.n1116 VDDD 0.0590938
R5133 VDDD.n1006 VDDD 0.0577917
R5134 VDDD.n2492 VDDD 0.0343542
R5135 VDDD.n1476 VDDD 0.0239375
R5136 VDDD.n1872 VDDD 0.0226354
R5137 VDDD.n1844 VDDD 0.0226354
R5138 VDDD VDDD.n1884 0.0226354
R5139 VDDD VDDD.n2012 0.0226354
R5140 VDDD VDDD.n2045 0.0226354
R5141 VDDD VDDD.n2078 0.0226354
R5142 VDDD VDDD.n2111 0.0226354
R5143 VDDD VDDD.n2144 0.0226354
R5144 VDDD VDDD.n2275 0.0226354
R5145 VDDD VDDD.n2308 0.0226354
R5146 VDDD VDDD.n2341 0.0226354
R5147 VDDD VDDD.n2374 0.0226354
R5148 VDDD VDDD.n2407 0.0226354
R5149 VDDD VDDD.n2440 0.0226354
R5150 VDDD VDDD.n1699 0.0226354
R5151 VDDD VDDD.n1732 0.0226354
R5152 VDDD VDDD.n1765 0.0226354
R5153 VDDD VDDD.n1798 0.0226354
R5154 VDDD.n1640 VDDD 0.0226354
R5155 VDDD.n1608 VDDD 0.0226354
R5156 VDDD.n1575 VDDD 0.0226354
R5157 VDDD.n1542 VDDD 0.0226354
R5158 VDDD.n1509 VDDD 0.0226354
R5159 VDDD.n1104 VDDD 0.0226354
R5160 VDDD VDDD.n1116 0.0226354
R5161 VDDD.n1150 VDDD 0.0226354
R5162 VDDD VDDD.n1153 0.0226354
R5163 VDDD.n1187 VDDD 0.0226354
R5164 VDDD VDDD.n1190 0.0226354
R5165 VDDD.n1224 VDDD 0.0226354
R5166 VDDD VDDD.n1227 0.0226354
R5167 VDDD.n1261 VDDD 0.0226354
R5168 VDDD VDDD.n1264 0.0226354
R5169 VDDD VDDD.n1303 0.0226354
R5170 VDDD VDDD.n672 0.0226354
R5171 VDDD.n704 VDDD 0.0226354
R5172 VDDD VDDD.n741 0.0226354
R5173 VDDD.n773 VDDD 0.0226354
R5174 VDDD VDDD.n810 0.0226354
R5175 VDDD.n842 VDDD 0.0226354
R5176 VDDD VDDD.n879 0.0226354
R5177 VDDD.n911 VDDD 0.0226354
R5178 VDDD VDDD.n948 0.0226354
R5179 VDDD.n980 VDDD 0.0226354
R5180 VDDD.n605 VDDD 0.0226354
R5181 VDDD.n568 VDDD 0.0226354
R5182 VDDD.n536 VDDD 0.0226354
R5183 VDDD.n499 VDDD 0.0226354
R5184 VDDD.n467 VDDD 0.0226354
R5185 VDDD.n430 VDDD 0.0226354
R5186 VDDD.n398 VDDD 0.0226354
R5187 VDDD.n361 VDDD 0.0226354
R5188 VDDD.n329 VDDD 0.0226354
R5189 VDDD.n292 VDDD 0.0226354
R5190 VDDD VDDD.n1005 0.0213333
R5191 VDDD.n271 VDDD 0.0213333
R5192 VDDD VDDD.n2492 0.0213333
R5193 VDDD VDDD.n2473 0.016125
R5194 a_n1709_3557.n1 a_n1709_3557.t2 530.01
R5195 a_n1709_3557.t1 a_n1709_3557.n5 421.021
R5196 a_n1709_3557.n0 a_n1709_3557.t3 337.142
R5197 a_n1709_3557.n3 a_n1709_3557.t0 280.223
R5198 a_n1709_3557.n4 a_n1709_3557.t5 263.173
R5199 a_n1709_3557.n4 a_n1709_3557.t6 227.826
R5200 a_n1709_3557.n0 a_n1709_3557.t4 199.762
R5201 a_n1709_3557.n2 a_n1709_3557.n1 170.81
R5202 a_n1709_3557.n2 a_n1709_3557.n0 167.321
R5203 a_n1709_3557.n5 a_n1709_3557.n4 152
R5204 a_n1709_3557.n1 a_n1709_3557.t7 141.923
R5205 a_n1709_3557.n3 a_n1709_3557.n2 10.8376
R5206 a_n1709_3557.n5 a_n1709_3557.n3 2.50485
R5207 a_n1193_3557.n3 a_n1193_3557.n2 674.338
R5208 a_n1193_3557.n1 a_n1193_3557.t5 332.58
R5209 a_n1193_3557.n2 a_n1193_3557.n0 284.012
R5210 a_n1193_3557.n2 a_n1193_3557.n1 253.648
R5211 a_n1193_3557.n1 a_n1193_3557.t4 168.701
R5212 a_n1193_3557.n3 a_n1193_3557.t2 96.1553
R5213 a_n1193_3557.t0 a_n1193_3557.n3 65.6672
R5214 a_n1193_3557.n0 a_n1193_3557.t3 65.0005
R5215 a_n1193_3557.n0 a_n1193_3557.t1 45.0005
R5216 a_n1085_3923.t0 a_n1085_3923.n0 1327.82
R5217 a_n1085_3923.n0 a_n1085_3923.t2 194.655
R5218 a_n1085_3923.n0 a_n1085_3923.t1 63.3219
R5219 a_n4909_n9650.n3 a_n4909_n9650.n2 674.338
R5220 a_n4909_n9650.n1 a_n4909_n9650.t4 332.58
R5221 a_n4909_n9650.n2 a_n4909_n9650.n0 284.012
R5222 a_n4909_n9650.n2 a_n4909_n9650.n1 253.648
R5223 a_n4909_n9650.n1 a_n4909_n9650.t5 168.701
R5224 a_n4909_n9650.t0 a_n4909_n9650.n3 96.1553
R5225 a_n4909_n9650.n3 a_n4909_n9650.t2 65.6672
R5226 a_n4909_n9650.n0 a_n4909_n9650.t1 65.0005
R5227 a_n4909_n9650.n0 a_n4909_n9650.t3 45.0005
R5228 a_n4691_n10054.n3 a_n4691_n10054.n2 647.119
R5229 a_n4691_n10054.n1 a_n4691_n10054.t5 350.253
R5230 a_n4691_n10054.n2 a_n4691_n10054.n0 260.339
R5231 a_n4691_n10054.n2 a_n4691_n10054.n1 246.119
R5232 a_n4691_n10054.n1 a_n4691_n10054.t4 189.588
R5233 a_n4691_n10054.n3 a_n4691_n10054.t0 89.1195
R5234 a_n4691_n10054.n0 a_n4691_n10054.t1 63.3338
R5235 a_n4691_n10054.t2 a_n4691_n10054.n3 41.0422
R5236 a_n4691_n10054.n0 a_n4691_n10054.t3 31.9797
R5237 CLKS.n334 CLKS.t23 408.63
R5238 CLKS.n323 CLKS.t59 408.63
R5239 CLKS.n312 CLKS.t17 408.63
R5240 CLKS.n301 CLKS.t61 408.63
R5241 CLKS.n291 CLKS.t53 408.63
R5242 CLKS.n282 CLKS.t87 408.63
R5243 CLKS.n274 CLKS.t30 408.63
R5244 CLKS.n266 CLKS.t113 408.63
R5245 CLKS.n258 CLKS.t125 408.63
R5246 CLKS.n250 CLKS.t98 408.63
R5247 CLKS.n211 CLKS.t19 408.63
R5248 CLKS.n222 CLKS.t135 408.63
R5249 CLKS.n188 CLKS.t51 408.63
R5250 CLKS.n199 CLKS.t47 408.63
R5251 CLKS.n165 CLKS.t46 408.63
R5252 CLKS.n176 CLKS.t97 408.63
R5253 CLKS.n142 CLKS.t78 408.63
R5254 CLKS.n153 CLKS.t18 408.63
R5255 CLKS.n119 CLKS.t136 408.63
R5256 CLKS.n130 CLKS.t22 408.63
R5257 CLKS.n96 CLKS.t132 408.63
R5258 CLKS.n107 CLKS.t117 408.63
R5259 CLKS.n73 CLKS.t88 408.63
R5260 CLKS.n84 CLKS.t74 408.63
R5261 CLKS.n50 CLKS.t57 408.63
R5262 CLKS.n61 CLKS.t39 408.63
R5263 CLKS.n27 CLKS.t40 408.63
R5264 CLKS.n38 CLKS.t62 408.63
R5265 CLKS.n5 CLKS.t138 408.63
R5266 CLKS.n16 CLKS.t52 408.63
R5267 CLKS.n337 CLKS.t99 347.577
R5268 CLKS.n326 CLKS.t32 347.577
R5269 CLKS.n315 CLKS.t21 347.577
R5270 CLKS.n304 CLKS.t92 347.577
R5271 CLKS.n294 CLKS.t27 347.577
R5272 CLKS.n285 CLKS.t116 347.577
R5273 CLKS.n277 CLKS.t70 347.577
R5274 CLKS.n269 CLKS.t42 347.577
R5275 CLKS.n261 CLKS.t140 347.577
R5276 CLKS.n253 CLKS.t100 347.577
R5277 CLKS.n207 CLKS.t37 347.577
R5278 CLKS.n218 CLKS.t56 347.577
R5279 CLKS.n184 CLKS.t64 347.577
R5280 CLKS.n195 CLKS.t90 347.577
R5281 CLKS.n161 CLKS.t119 347.577
R5282 CLKS.n172 CLKS.t26 347.577
R5283 CLKS.n138 CLKS.t108 347.577
R5284 CLKS.n149 CLKS.t76 347.577
R5285 CLKS.n115 CLKS.t137 347.577
R5286 CLKS.n126 CLKS.t123 347.577
R5287 CLKS.n92 CLKS.t81 347.577
R5288 CLKS.n103 CLKS.t33 347.577
R5289 CLKS.n69 CLKS.t86 347.577
R5290 CLKS.n80 CLKS.t93 347.577
R5291 CLKS.n46 CLKS.t29 347.577
R5292 CLKS.n57 CLKS.t94 347.577
R5293 CLKS.n23 CLKS.t110 347.577
R5294 CLKS.n34 CLKS.t58 347.577
R5295 CLKS.n1 CLKS.t122 347.577
R5296 CLKS.n12 CLKS.t131 347.577
R5297 CLKS.n346 CLKS.t106 261.887
R5298 CLKS.n348 CLKS.t139 261.887
R5299 CLKS.n229 CLKS.t63 230.576
R5300 CLKS.n242 CLKS.n237 205.28
R5301 CLKS.n241 CLKS.n238 205.28
R5302 CLKS.n240 CLKS.n239 205.28
R5303 CLKS.n232 CLKS.n231 205.28
R5304 CLKS.n337 CLKS.t20 193.337
R5305 CLKS.n326 CLKS.t28 193.337
R5306 CLKS.n315 CLKS.t79 193.337
R5307 CLKS.n304 CLKS.t48 193.337
R5308 CLKS.n294 CLKS.t54 193.337
R5309 CLKS.n285 CLKS.t60 193.337
R5310 CLKS.n277 CLKS.t24 193.337
R5311 CLKS.n269 CLKS.t105 193.337
R5312 CLKS.n261 CLKS.t83 193.337
R5313 CLKS.n253 CLKS.t50 193.337
R5314 CLKS.n207 CLKS.t121 193.337
R5315 CLKS.n218 CLKS.t38 193.337
R5316 CLKS.n184 CLKS.t35 193.337
R5317 CLKS.n195 CLKS.t67 193.337
R5318 CLKS.n161 CLKS.t80 193.337
R5319 CLKS.n172 CLKS.t124 193.337
R5320 CLKS.n138 CLKS.t72 193.337
R5321 CLKS.n149 CLKS.t112 193.337
R5322 CLKS.n115 CLKS.t95 193.337
R5323 CLKS.n126 CLKS.t141 193.337
R5324 CLKS.n92 CLKS.t49 193.337
R5325 CLKS.n103 CLKS.t84 193.337
R5326 CLKS.n69 CLKS.t55 193.337
R5327 CLKS.n80 CLKS.t89 193.337
R5328 CLKS.n46 CLKS.t109 193.337
R5329 CLKS.n57 CLKS.t31 193.337
R5330 CLKS.n23 CLKS.t75 193.337
R5331 CLKS.n34 CLKS.t115 193.337
R5332 CLKS.n1 CLKS.t82 193.337
R5333 CLKS.n12 CLKS.t128 193.337
R5334 CLKS CLKS.n282 165.201
R5335 CLKS CLKS.n274 165.201
R5336 CLKS CLKS.n266 165.201
R5337 CLKS CLKS.n258 165.201
R5338 CLKS CLKS.n250 165.201
R5339 CLKS.n335 CLKS.n334 165.072
R5340 CLKS.n324 CLKS.n323 165.072
R5341 CLKS.n313 CLKS.n312 165.072
R5342 CLKS.n302 CLKS.n301 165.072
R5343 CLKS.n292 CLKS.n291 165.072
R5344 CLKS.n212 CLKS.n211 165.072
R5345 CLKS.n223 CLKS.n222 165.072
R5346 CLKS.n189 CLKS.n188 165.072
R5347 CLKS.n200 CLKS.n199 165.072
R5348 CLKS.n166 CLKS.n165 165.072
R5349 CLKS.n177 CLKS.n176 165.072
R5350 CLKS.n143 CLKS.n142 165.072
R5351 CLKS.n154 CLKS.n153 165.072
R5352 CLKS.n120 CLKS.n119 165.072
R5353 CLKS.n131 CLKS.n130 165.072
R5354 CLKS.n97 CLKS.n96 165.072
R5355 CLKS.n108 CLKS.n107 165.072
R5356 CLKS.n74 CLKS.n73 165.072
R5357 CLKS.n85 CLKS.n84 165.072
R5358 CLKS.n51 CLKS.n50 165.072
R5359 CLKS.n62 CLKS.n61 165.072
R5360 CLKS.n28 CLKS.n27 165.072
R5361 CLKS.n39 CLKS.n38 165.072
R5362 CLKS.n6 CLKS.n5 165.072
R5363 CLKS.n17 CLKS.n16 165.072
R5364 CLKS.n229 CLKS.t130 158.275
R5365 CLKS.n346 CLKS.t66 155.847
R5366 CLKS.n348 CLKS.t120 155.847
R5367 CLKS.n230 CLKS.n229 154.133
R5368 CLKS.n347 CLKS.n346 153.13
R5369 CLKS.n338 CLKS.n337 152
R5370 CLKS.n327 CLKS.n326 152
R5371 CLKS.n316 CLKS.n315 152
R5372 CLKS.n305 CLKS.n304 152
R5373 CLKS.n295 CLKS.n294 152
R5374 CLKS.n286 CLKS.n285 152
R5375 CLKS.n278 CLKS.n277 152
R5376 CLKS.n270 CLKS.n269 152
R5377 CLKS.n262 CLKS.n261 152
R5378 CLKS.n254 CLKS.n253 152
R5379 CLKS.n349 CLKS.n348 152
R5380 CLKS.n208 CLKS.n207 152
R5381 CLKS.n219 CLKS.n218 152
R5382 CLKS.n185 CLKS.n184 152
R5383 CLKS.n196 CLKS.n195 152
R5384 CLKS.n162 CLKS.n161 152
R5385 CLKS.n173 CLKS.n172 152
R5386 CLKS.n139 CLKS.n138 152
R5387 CLKS.n150 CLKS.n149 152
R5388 CLKS.n116 CLKS.n115 152
R5389 CLKS.n127 CLKS.n126 152
R5390 CLKS.n93 CLKS.n92 152
R5391 CLKS.n104 CLKS.n103 152
R5392 CLKS.n70 CLKS.n69 152
R5393 CLKS.n81 CLKS.n80 152
R5394 CLKS.n47 CLKS.n46 152
R5395 CLKS.n58 CLKS.n57 152
R5396 CLKS.n24 CLKS.n23 152
R5397 CLKS.n35 CLKS.n34 152
R5398 CLKS.n2 CLKS.n1 152
R5399 CLKS.n13 CLKS.n12 152
R5400 CLKS.n334 CLKS.t133 132.282
R5401 CLKS.n323 CLKS.t102 132.282
R5402 CLKS.n312 CLKS.t68 132.282
R5403 CLKS.n301 CLKS.t77 132.282
R5404 CLKS.n291 CLKS.t45 132.282
R5405 CLKS.n282 CLKS.t91 132.282
R5406 CLKS.n274 CLKS.t34 132.282
R5407 CLKS.n266 CLKS.t118 132.282
R5408 CLKS.n258 CLKS.t129 132.282
R5409 CLKS.n250 CLKS.t101 132.282
R5410 CLKS.n211 CLKS.t41 132.282
R5411 CLKS.n222 CLKS.t73 132.282
R5412 CLKS.n188 CLKS.t69 132.282
R5413 CLKS.n199 CLKS.t107 132.282
R5414 CLKS.n165 CLKS.t103 132.282
R5415 CLKS.n176 CLKS.t25 132.282
R5416 CLKS.n142 CLKS.t96 132.282
R5417 CLKS.n153 CLKS.t16 132.282
R5418 CLKS.n119 CLKS.t127 132.282
R5419 CLKS.n130 CLKS.t44 132.282
R5420 CLKS.n96 CLKS.t114 132.282
R5421 CLKS.n107 CLKS.t36 132.282
R5422 CLKS.n73 CLKS.t126 132.282
R5423 CLKS.n84 CLKS.t43 132.282
R5424 CLKS.n50 CLKS.t85 132.282
R5425 CLKS.n61 CLKS.t134 132.282
R5426 CLKS.n27 CLKS.t65 132.282
R5427 CLKS.n38 CLKS.t104 132.282
R5428 CLKS.n5 CLKS.t71 132.282
R5429 CLKS.n16 CLKS.t111 132.282
R5430 CLKS.n246 CLKS.n233 99.1759
R5431 CLKS.n245 CLKS.n234 99.1759
R5432 CLKS.n244 CLKS.n235 99.1759
R5433 CLKS.n243 CLKS.n236 99.1759
R5434 CLKS.n351 CLKS 52.8283
R5435 CLKS.n249 CLKS 51.414
R5436 CLKS.n242 CLKS.n241 38.4005
R5437 CLKS.n241 CLKS.n240 38.4005
R5438 CLKS.n240 CLKS.n232 38.4005
R5439 CLKS.n345 CLKS 36.5456
R5440 CLKS CLKS.n242 36.4472
R5441 CLKS.n246 CLKS.n245 34.3584
R5442 CLKS.n245 CLKS.n244 34.3584
R5443 CLKS.n244 CLKS.n243 34.3584
R5444 CLKS.n247 CLKS.n232 31.0358
R5445 CLKS.n243 CLKS 27.7875
R5446 CLKS.n237 CLKS.t5 26.5955
R5447 CLKS.n237 CLKS.t7 26.5955
R5448 CLKS.n238 CLKS.t11 26.5955
R5449 CLKS.n238 CLKS.t10 26.5955
R5450 CLKS.n239 CLKS.t2 26.5955
R5451 CLKS.n239 CLKS.t12 26.5955
R5452 CLKS.n231 CLKS.t14 26.5955
R5453 CLKS.n231 CLKS.t9 26.5955
R5454 CLKS CLKS.n246 25.611
R5455 CLKS.n233 CLKS.t1 24.9236
R5456 CLKS.n233 CLKS.t4 24.9236
R5457 CLKS.n234 CLKS.t13 24.9236
R5458 CLKS.n234 CLKS.t0 24.9236
R5459 CLKS.n235 CLKS.t15 24.9236
R5460 CLKS.n235 CLKS.t6 24.9236
R5461 CLKS.n236 CLKS.t8 24.9236
R5462 CLKS.n236 CLKS.t3 24.9236
R5463 CLKS.n350 CLKS.n347 15.2668
R5464 CLKS.n350 CLKS.n349 14.8245
R5465 CLKS CLKS.n333 14.0185
R5466 CLKS CLKS.n322 14.0185
R5467 CLKS CLKS.n311 14.0185
R5468 CLKS CLKS.n300 14.0185
R5469 CLKS CLKS.n290 14.0185
R5470 CLKS.n209 CLKS 14.0185
R5471 CLKS.n186 CLKS 14.0185
R5472 CLKS.n163 CLKS 14.0185
R5473 CLKS.n140 CLKS 14.0185
R5474 CLKS.n117 CLKS 14.0185
R5475 CLKS.n94 CLKS 14.0185
R5476 CLKS.n71 CLKS 14.0185
R5477 CLKS.n48 CLKS 14.0185
R5478 CLKS.n25 CLKS 14.0185
R5479 CLKS.n3 CLKS 14.0185
R5480 CLKS.n220 CLKS 13.8909
R5481 CLKS.n197 CLKS 13.8909
R5482 CLKS.n174 CLKS 13.8909
R5483 CLKS.n151 CLKS 13.8909
R5484 CLKS.n128 CLKS 13.8909
R5485 CLKS.n105 CLKS 13.8909
R5486 CLKS.n82 CLKS 13.8909
R5487 CLKS.n59 CLKS 13.8909
R5488 CLKS.n36 CLKS 13.8909
R5489 CLKS.n14 CLKS 13.8909
R5490 CLKS.n287 CLKS 13.8338
R5491 CLKS.n279 CLKS 13.8338
R5492 CLKS.n271 CLKS 13.8338
R5493 CLKS.n263 CLKS 13.8338
R5494 CLKS.n255 CLKS 13.8338
R5495 CLKS.n286 CLKS.n284 12.0681
R5496 CLKS.n278 CLKS.n276 12.0681
R5497 CLKS.n270 CLKS.n268 12.0681
R5498 CLKS.n262 CLKS.n260 12.0681
R5499 CLKS.n254 CLKS.n252 12.0681
R5500 CLKS.n248 CLKS.n230 9.62563
R5501 CLKS CLKS.n351 9.49418
R5502 CLKS.n210 CLKS.n209 9.35757
R5503 CLKS.n187 CLKS.n186 9.35757
R5504 CLKS.n164 CLKS.n163 9.35757
R5505 CLKS.n141 CLKS.n140 9.35757
R5506 CLKS.n118 CLKS.n117 9.35757
R5507 CLKS.n95 CLKS.n94 9.35757
R5508 CLKS.n72 CLKS.n71 9.35757
R5509 CLKS.n49 CLKS.n48 9.35757
R5510 CLKS.n26 CLKS.n25 9.35757
R5511 CLKS.n4 CLKS.n3 9.35757
R5512 CLKS.n215 CLKS.n206 9.33714
R5513 CLKS.n192 CLKS.n183 9.33714
R5514 CLKS.n169 CLKS.n160 9.33714
R5515 CLKS.n146 CLKS.n137 9.33714
R5516 CLKS.n123 CLKS.n114 9.33714
R5517 CLKS.n100 CLKS.n91 9.33714
R5518 CLKS.n77 CLKS.n68 9.33714
R5519 CLKS.n54 CLKS.n45 9.33714
R5520 CLKS.n31 CLKS.n22 9.33714
R5521 CLKS.n9 CLKS.n0 9.33714
R5522 CLKS.n342 CLKS.n333 9.3029
R5523 CLKS.n331 CLKS.n322 9.3029
R5524 CLKS.n320 CLKS.n311 9.3029
R5525 CLKS.n309 CLKS.n300 9.3029
R5526 CLKS.n299 CLKS.n290 9.3029
R5527 CLKS.n248 CLKS.n247 9.3005
R5528 CLKS.n340 CLKS.n339 9.3005
R5529 CLKS.n329 CLKS.n328 9.3005
R5530 CLKS.n318 CLKS.n317 9.3005
R5531 CLKS.n307 CLKS.n306 9.3005
R5532 CLKS.n297 CLKS.n296 9.3005
R5533 CLKS.n217 CLKS.n216 9.3005
R5534 CLKS.n194 CLKS.n193 9.3005
R5535 CLKS.n171 CLKS.n170 9.3005
R5536 CLKS.n148 CLKS.n147 9.3005
R5537 CLKS.n125 CLKS.n124 9.3005
R5538 CLKS.n102 CLKS.n101 9.3005
R5539 CLKS.n79 CLKS.n78 9.3005
R5540 CLKS.n56 CLKS.n55 9.3005
R5541 CLKS.n33 CLKS.n32 9.3005
R5542 CLKS.n11 CLKS.n10 9.3005
R5543 CLKS.n310 CLKS.n299 9.14473
R5544 CLKS CLKS.n286 8.82212
R5545 CLKS CLKS.n278 8.82212
R5546 CLKS CLKS.n270 8.82212
R5547 CLKS CLKS.n262 8.82212
R5548 CLKS CLKS.n254 8.82212
R5549 CLKS.n351 CLKS.n345 6.733
R5550 CLKS CLKS.n248 5.90341
R5551 CLKS.n227 CLKS.n226 5.12373
R5552 CLKS.n204 CLKS.n203 5.12373
R5553 CLKS.n181 CLKS.n180 5.12373
R5554 CLKS.n158 CLKS.n157 5.12373
R5555 CLKS.n135 CLKS.n134 5.12373
R5556 CLKS.n112 CLKS.n111 5.12373
R5557 CLKS.n89 CLKS.n88 5.12373
R5558 CLKS.n66 CLKS.n65 5.12373
R5559 CLKS.n43 CLKS.n42 5.12173
R5560 CLKS.n21 CLKS.n20 5.12173
R5561 CLKS.n338 CLKS 4.67077
R5562 CLKS.n327 CLKS 4.67077
R5563 CLKS.n316 CLKS 4.67077
R5564 CLKS.n305 CLKS 4.67077
R5565 CLKS.n295 CLKS 4.67077
R5566 CLKS CLKS.n208 4.67077
R5567 CLKS CLKS.n219 4.67077
R5568 CLKS CLKS.n185 4.67077
R5569 CLKS CLKS.n196 4.67077
R5570 CLKS CLKS.n162 4.67077
R5571 CLKS CLKS.n173 4.67077
R5572 CLKS CLKS.n139 4.67077
R5573 CLKS CLKS.n150 4.67077
R5574 CLKS CLKS.n116 4.67077
R5575 CLKS CLKS.n127 4.67077
R5576 CLKS CLKS.n93 4.67077
R5577 CLKS CLKS.n104 4.67077
R5578 CLKS CLKS.n70 4.67077
R5579 CLKS CLKS.n81 4.67077
R5580 CLKS CLKS.n47 4.67077
R5581 CLKS CLKS.n58 4.67077
R5582 CLKS CLKS.n24 4.67077
R5583 CLKS CLKS.n35 4.67077
R5584 CLKS CLKS.n2 4.67077
R5585 CLKS CLKS.n13 4.67077
R5586 CLKS.n265 CLKS.n257 4.64473
R5587 CLKS.n273 CLKS.n265 4.64473
R5588 CLKS.n281 CLKS.n273 4.64473
R5589 CLKS.n321 CLKS.n310 4.64473
R5590 CLKS.n332 CLKS.n321 4.64473
R5591 CLKS.n343 CLKS.n332 4.64473
R5592 CLKS.n227 CLKS.n215 4.62373
R5593 CLKS.n204 CLKS.n192 4.62373
R5594 CLKS.n181 CLKS.n169 4.62373
R5595 CLKS.n158 CLKS.n146 4.62373
R5596 CLKS.n135 CLKS.n123 4.62373
R5597 CLKS.n112 CLKS.n100 4.62373
R5598 CLKS.n89 CLKS.n77 4.62373
R5599 CLKS.n66 CLKS.n54 4.62373
R5600 CLKS.n43 CLKS.n31 4.62173
R5601 CLKS.n21 CLKS.n9 4.62173
R5602 CLKS.n289 CLKS.n288 4.60534
R5603 CLKS.n44 CLKS.n21 4.53843
R5604 CLKS.n230 CLKS 4.53383
R5605 CLKS.n333 CLKS 4.53383
R5606 CLKS.n322 CLKS 4.53383
R5607 CLKS.n311 CLKS 4.53383
R5608 CLKS.n300 CLKS 4.53383
R5609 CLKS.n290 CLKS 4.53383
R5610 CLKS.n209 CLKS 4.53383
R5611 CLKS.n186 CLKS 4.53383
R5612 CLKS.n163 CLKS 4.53383
R5613 CLKS.n140 CLKS 4.53383
R5614 CLKS.n117 CLKS 4.53383
R5615 CLKS.n94 CLKS 4.53383
R5616 CLKS.n71 CLKS 4.53383
R5617 CLKS.n48 CLKS 4.53383
R5618 CLKS.n25 CLKS 4.53383
R5619 CLKS.n3 CLKS 4.53383
R5620 CLKS.n289 CLKS.n281 4.50965
R5621 CLKS.n257 CLKS.n256 4.5005
R5622 CLKS.n265 CLKS.n264 4.5005
R5623 CLKS.n273 CLKS.n272 4.5005
R5624 CLKS.n281 CLKS.n280 4.5005
R5625 CLKS.n310 CLKS.n309 4.5005
R5626 CLKS.n321 CLKS.n320 4.5005
R5627 CLKS.n332 CLKS.n331 4.5005
R5628 CLKS.n343 CLKS.n342 4.5005
R5629 CLKS.n257 CLKS 3.93319
R5630 CLKS.n349 CLKS 3.8405
R5631 CLKS.n249 CLKS 3.543
R5632 CLKS.n44 CLKS.n43 3.4105
R5633 CLKS.n67 CLKS.n66 3.4105
R5634 CLKS.n90 CLKS.n89 3.4105
R5635 CLKS.n113 CLKS.n112 3.4105
R5636 CLKS.n136 CLKS.n135 3.4105
R5637 CLKS.n159 CLKS.n158 3.4105
R5638 CLKS.n182 CLKS.n181 3.4105
R5639 CLKS.n205 CLKS.n204 3.4105
R5640 CLKS.n228 CLKS.n227 3.4105
R5641 CLKS.n247 CLKS 3.4005
R5642 CLKS.n347 CLKS 3.2005
R5643 CLKS.n345 CLKS.n249 3.12925
R5644 CLKS.n339 CLKS 2.94104
R5645 CLKS.n328 CLKS 2.94104
R5646 CLKS.n317 CLKS 2.94104
R5647 CLKS.n306 CLKS 2.94104
R5648 CLKS.n296 CLKS 2.94104
R5649 CLKS.n206 CLKS 2.94104
R5650 CLKS.n217 CLKS 2.94104
R5651 CLKS.n183 CLKS 2.94104
R5652 CLKS.n194 CLKS 2.94104
R5653 CLKS.n160 CLKS 2.94104
R5654 CLKS.n171 CLKS 2.94104
R5655 CLKS.n137 CLKS 2.94104
R5656 CLKS.n148 CLKS 2.94104
R5657 CLKS.n114 CLKS 2.94104
R5658 CLKS.n125 CLKS 2.94104
R5659 CLKS.n91 CLKS 2.94104
R5660 CLKS.n102 CLKS 2.94104
R5661 CLKS.n68 CLKS 2.94104
R5662 CLKS.n79 CLKS 2.94104
R5663 CLKS.n45 CLKS 2.94104
R5664 CLKS.n56 CLKS 2.94104
R5665 CLKS.n22 CLKS 2.94104
R5666 CLKS.n33 CLKS 2.94104
R5667 CLKS.n0 CLKS 2.94104
R5668 CLKS.n11 CLKS 2.94104
R5669 CLKS.n339 CLKS.n338 2.76807
R5670 CLKS.n328 CLKS.n327 2.76807
R5671 CLKS.n317 CLKS.n316 2.76807
R5672 CLKS.n306 CLKS.n305 2.76807
R5673 CLKS.n296 CLKS.n295 2.76807
R5674 CLKS.n208 CLKS.n206 2.76807
R5675 CLKS.n219 CLKS.n217 2.76807
R5676 CLKS.n185 CLKS.n183 2.76807
R5677 CLKS.n196 CLKS.n194 2.76807
R5678 CLKS.n162 CLKS.n160 2.76807
R5679 CLKS.n173 CLKS.n171 2.76807
R5680 CLKS.n139 CLKS.n137 2.76807
R5681 CLKS.n150 CLKS.n148 2.76807
R5682 CLKS.n116 CLKS.n114 2.76807
R5683 CLKS.n127 CLKS.n125 2.76807
R5684 CLKS.n93 CLKS.n91 2.76807
R5685 CLKS.n104 CLKS.n102 2.76807
R5686 CLKS.n70 CLKS.n68 2.76807
R5687 CLKS.n81 CLKS.n79 2.76807
R5688 CLKS.n47 CLKS.n45 2.76807
R5689 CLKS.n58 CLKS.n56 2.76807
R5690 CLKS.n24 CLKS.n22 2.76807
R5691 CLKS.n35 CLKS.n33 2.76807
R5692 CLKS.n2 CLKS.n0 2.76807
R5693 CLKS.n13 CLKS.n11 2.76807
R5694 CLKS.n344 CLKS.n343 2.42838
R5695 CLKS CLKS.n336 2.36657
R5696 CLKS CLKS.n325 2.36657
R5697 CLKS CLKS.n314 2.36657
R5698 CLKS CLKS.n303 2.36657
R5699 CLKS CLKS.n293 2.36657
R5700 CLKS.n283 CLKS 2.36657
R5701 CLKS.n275 CLKS 2.36657
R5702 CLKS.n267 CLKS 2.36657
R5703 CLKS.n259 CLKS 2.36657
R5704 CLKS.n251 CLKS 2.36657
R5705 CLKS.n214 CLKS.n213 2.32193
R5706 CLKS.n225 CLKS.n224 2.32193
R5707 CLKS.n191 CLKS.n190 2.32193
R5708 CLKS.n202 CLKS.n201 2.32193
R5709 CLKS.n168 CLKS.n167 2.32193
R5710 CLKS.n179 CLKS.n178 2.32193
R5711 CLKS.n145 CLKS.n144 2.32193
R5712 CLKS.n156 CLKS.n155 2.32193
R5713 CLKS.n122 CLKS.n121 2.32193
R5714 CLKS.n133 CLKS.n132 2.32193
R5715 CLKS.n99 CLKS.n98 2.32193
R5716 CLKS.n110 CLKS.n109 2.32193
R5717 CLKS.n76 CLKS.n75 2.32193
R5718 CLKS.n87 CLKS.n86 2.32193
R5719 CLKS.n53 CLKS.n52 2.32193
R5720 CLKS.n64 CLKS.n63 2.32193
R5721 CLKS.n30 CLKS.n29 2.32193
R5722 CLKS.n41 CLKS.n40 2.32193
R5723 CLKS.n8 CLKS.n7 2.32193
R5724 CLKS.n19 CLKS.n18 2.32193
R5725 CLKS CLKS.n228 1.68695
R5726 CLKS CLKS.n344 1.50531
R5727 CLKS.n214 CLKS 1.35467
R5728 CLKS.n225 CLKS 1.35467
R5729 CLKS.n191 CLKS 1.35467
R5730 CLKS.n202 CLKS 1.35467
R5731 CLKS.n168 CLKS 1.35467
R5732 CLKS.n179 CLKS 1.35467
R5733 CLKS.n145 CLKS 1.35467
R5734 CLKS.n156 CLKS 1.35467
R5735 CLKS.n122 CLKS 1.35467
R5736 CLKS.n133 CLKS 1.35467
R5737 CLKS.n99 CLKS 1.35467
R5738 CLKS.n110 CLKS 1.35467
R5739 CLKS.n76 CLKS 1.35467
R5740 CLKS.n87 CLKS 1.35467
R5741 CLKS.n53 CLKS 1.35467
R5742 CLKS.n64 CLKS 1.35467
R5743 CLKS.n30 CLKS 1.35467
R5744 CLKS.n41 CLKS 1.35467
R5745 CLKS.n8 CLKS 1.35467
R5746 CLKS.n19 CLKS 1.35467
R5747 CLKS CLKS.n350 1.19762
R5748 CLKS.n90 CLKS.n67 1.12915
R5749 CLKS.n113 CLKS.n90 1.12915
R5750 CLKS.n136 CLKS.n113 1.12915
R5751 CLKS.n159 CLKS.n136 1.12915
R5752 CLKS.n182 CLKS.n159 1.12915
R5753 CLKS.n205 CLKS.n182 1.12915
R5754 CLKS.n228 CLKS.n205 1.12915
R5755 CLKS.n67 CLKS.n44 1.12909
R5756 CLKS.n344 CLKS.n289 0.654346
R5757 CLKS.n336 CLKS 0.580857
R5758 CLKS.n325 CLKS 0.580857
R5759 CLKS.n314 CLKS 0.580857
R5760 CLKS.n303 CLKS 0.580857
R5761 CLKS.n293 CLKS 0.580857
R5762 CLKS.n213 CLKS 0.580857
R5763 CLKS.n224 CLKS 0.580857
R5764 CLKS.n190 CLKS 0.580857
R5765 CLKS.n201 CLKS 0.580857
R5766 CLKS.n167 CLKS 0.580857
R5767 CLKS.n178 CLKS 0.580857
R5768 CLKS.n144 CLKS 0.580857
R5769 CLKS.n155 CLKS 0.580857
R5770 CLKS.n121 CLKS 0.580857
R5771 CLKS.n132 CLKS 0.580857
R5772 CLKS.n98 CLKS 0.580857
R5773 CLKS.n109 CLKS 0.580857
R5774 CLKS.n75 CLKS 0.580857
R5775 CLKS.n86 CLKS 0.580857
R5776 CLKS.n52 CLKS 0.580857
R5777 CLKS.n63 CLKS 0.580857
R5778 CLKS.n29 CLKS 0.580857
R5779 CLKS.n40 CLKS 0.580857
R5780 CLKS.n7 CLKS 0.580857
R5781 CLKS.n18 CLKS 0.580857
R5782 CLKS.n283 CLKS 0.527286
R5783 CLKS.n275 CLKS 0.527286
R5784 CLKS.n267 CLKS 0.527286
R5785 CLKS.n259 CLKS 0.527286
R5786 CLKS.n251 CLKS 0.527286
R5787 CLKS.n335 CLKS 0.225552
R5788 CLKS.n324 CLKS 0.225552
R5789 CLKS.n313 CLKS 0.225552
R5790 CLKS.n302 CLKS 0.225552
R5791 CLKS.n292 CLKS 0.225552
R5792 CLKS.n212 CLKS 0.225552
R5793 CLKS.n223 CLKS 0.225552
R5794 CLKS.n189 CLKS 0.225552
R5795 CLKS.n200 CLKS 0.225552
R5796 CLKS.n166 CLKS 0.225552
R5797 CLKS.n177 CLKS 0.225552
R5798 CLKS.n143 CLKS 0.225552
R5799 CLKS.n154 CLKS 0.225552
R5800 CLKS.n120 CLKS 0.225552
R5801 CLKS.n131 CLKS 0.225552
R5802 CLKS.n97 CLKS 0.225552
R5803 CLKS.n108 CLKS 0.225552
R5804 CLKS.n74 CLKS 0.225552
R5805 CLKS.n85 CLKS 0.225552
R5806 CLKS.n51 CLKS 0.225552
R5807 CLKS.n62 CLKS 0.225552
R5808 CLKS.n28 CLKS 0.225552
R5809 CLKS.n39 CLKS 0.225552
R5810 CLKS.n6 CLKS 0.225552
R5811 CLKS.n17 CLKS 0.225552
R5812 CLKS.n341 CLKS 0.139923
R5813 CLKS.n330 CLKS 0.139923
R5814 CLKS.n319 CLKS 0.139923
R5815 CLKS.n308 CLKS 0.139923
R5816 CLKS.n298 CLKS 0.139923
R5817 CLKS.n336 CLKS.n335 0.128681
R5818 CLKS.n325 CLKS.n324 0.128681
R5819 CLKS.n314 CLKS.n313 0.128681
R5820 CLKS.n303 CLKS.n302 0.128681
R5821 CLKS.n293 CLKS.n292 0.128681
R5822 CLKS.n213 CLKS.n212 0.128681
R5823 CLKS.n224 CLKS.n223 0.128681
R5824 CLKS.n190 CLKS.n189 0.128681
R5825 CLKS.n201 CLKS.n200 0.128681
R5826 CLKS.n167 CLKS.n166 0.128681
R5827 CLKS.n178 CLKS.n177 0.128681
R5828 CLKS.n144 CLKS.n143 0.128681
R5829 CLKS.n155 CLKS.n154 0.128681
R5830 CLKS.n121 CLKS.n120 0.128681
R5831 CLKS.n132 CLKS.n131 0.128681
R5832 CLKS.n98 CLKS.n97 0.128681
R5833 CLKS.n109 CLKS.n108 0.128681
R5834 CLKS.n75 CLKS.n74 0.128681
R5835 CLKS.n86 CLKS.n85 0.128681
R5836 CLKS.n52 CLKS.n51 0.128681
R5837 CLKS.n63 CLKS.n62 0.128681
R5838 CLKS.n29 CLKS.n28 0.128681
R5839 CLKS.n40 CLKS.n39 0.128681
R5840 CLKS.n7 CLKS.n6 0.128681
R5841 CLKS.n18 CLKS.n17 0.128681
R5842 CLKS.n215 CLKS.n210 0.0809468
R5843 CLKS.n192 CLKS.n187 0.0809468
R5844 CLKS.n169 CLKS.n164 0.0809468
R5845 CLKS.n146 CLKS.n141 0.0809468
R5846 CLKS.n123 CLKS.n118 0.0809468
R5847 CLKS.n100 CLKS.n95 0.0809468
R5848 CLKS.n77 CLKS.n72 0.0809468
R5849 CLKS.n54 CLKS.n49 0.0809468
R5850 CLKS.n31 CLKS.n26 0.0809468
R5851 CLKS.n9 CLKS.n4 0.0809468
R5852 CLKS.n226 CLKS.n221 0.0734167
R5853 CLKS.n203 CLKS.n198 0.0734167
R5854 CLKS.n180 CLKS.n175 0.0734167
R5855 CLKS.n157 CLKS.n152 0.0734167
R5856 CLKS.n134 CLKS.n129 0.0734167
R5857 CLKS.n111 CLKS.n106 0.0734167
R5858 CLKS.n88 CLKS.n83 0.0734167
R5859 CLKS.n65 CLKS.n60 0.0734167
R5860 CLKS.n42 CLKS.n37 0.0734167
R5861 CLKS.n20 CLKS.n15 0.0734167
R5862 CLKS.n288 CLKS 0.0726154
R5863 CLKS.n280 CLKS 0.0726154
R5864 CLKS.n272 CLKS 0.0726154
R5865 CLKS.n264 CLKS 0.0726154
R5866 CLKS.n256 CLKS 0.0726154
R5867 CLKS.n287 CLKS 0.0702115
R5868 CLKS.n279 CLKS 0.0702115
R5869 CLKS.n271 CLKS 0.0702115
R5870 CLKS.n263 CLKS 0.0702115
R5871 CLKS.n255 CLKS 0.0702115
R5872 CLKS.n342 CLKS 0.0678077
R5873 CLKS.n331 CLKS 0.0678077
R5874 CLKS.n320 CLKS 0.0678077
R5875 CLKS.n309 CLKS 0.0678077
R5876 CLKS.n299 CLKS 0.0678077
R5877 CLKS.n210 CLKS 0.063
R5878 CLKS.n187 CLKS 0.063
R5879 CLKS.n164 CLKS 0.063
R5880 CLKS.n141 CLKS 0.063
R5881 CLKS.n118 CLKS 0.063
R5882 CLKS.n95 CLKS 0.063
R5883 CLKS.n72 CLKS 0.063
R5884 CLKS.n49 CLKS 0.063
R5885 CLKS.n26 CLKS 0.063
R5886 CLKS.n4 CLKS 0.063
R5887 CLKS.n215 CLKS 0.0609167
R5888 CLKS.n226 CLKS 0.0609167
R5889 CLKS.n192 CLKS 0.0609167
R5890 CLKS.n203 CLKS 0.0609167
R5891 CLKS.n169 CLKS 0.0609167
R5892 CLKS.n180 CLKS 0.0609167
R5893 CLKS.n146 CLKS 0.0609167
R5894 CLKS.n157 CLKS 0.0609167
R5895 CLKS.n123 CLKS 0.0609167
R5896 CLKS.n134 CLKS 0.0609167
R5897 CLKS.n100 CLKS 0.0609167
R5898 CLKS.n111 CLKS 0.0609167
R5899 CLKS.n77 CLKS 0.0609167
R5900 CLKS.n88 CLKS 0.0609167
R5901 CLKS.n54 CLKS 0.0609167
R5902 CLKS.n65 CLKS 0.0609167
R5903 CLKS.n31 CLKS 0.0609167
R5904 CLKS.n42 CLKS 0.0609167
R5905 CLKS.n9 CLKS 0.0609167
R5906 CLKS.n20 CLKS 0.0609167
R5907 CLKS.n221 CLKS 0.0560556
R5908 CLKS.n198 CLKS 0.0560556
R5909 CLKS.n175 CLKS 0.0560556
R5910 CLKS.n152 CLKS 0.0560556
R5911 CLKS.n129 CLKS 0.0560556
R5912 CLKS.n106 CLKS 0.0560556
R5913 CLKS.n83 CLKS 0.0560556
R5914 CLKS.n60 CLKS 0.0560556
R5915 CLKS.n37 CLKS 0.0560556
R5916 CLKS.n15 CLKS 0.0560556
R5917 CLKS.n215 CLKS 0.050069
R5918 CLKS.n216 CLKS 0.050069
R5919 CLKS.n192 CLKS 0.050069
R5920 CLKS.n193 CLKS 0.050069
R5921 CLKS.n169 CLKS 0.050069
R5922 CLKS.n170 CLKS 0.050069
R5923 CLKS.n146 CLKS 0.050069
R5924 CLKS.n147 CLKS 0.050069
R5925 CLKS.n123 CLKS 0.050069
R5926 CLKS.n124 CLKS 0.050069
R5927 CLKS.n100 CLKS 0.050069
R5928 CLKS.n101 CLKS 0.050069
R5929 CLKS.n77 CLKS 0.050069
R5930 CLKS.n78 CLKS 0.050069
R5931 CLKS.n54 CLKS 0.050069
R5932 CLKS.n55 CLKS 0.050069
R5933 CLKS.n31 CLKS 0.050069
R5934 CLKS.n32 CLKS 0.050069
R5935 CLKS.n9 CLKS 0.050069
R5936 CLKS.n10 CLKS 0.050069
R5937 CLKS.n226 CLKS.n216 0.0371379
R5938 CLKS.n203 CLKS.n193 0.0371379
R5939 CLKS.n180 CLKS.n170 0.0371379
R5940 CLKS.n157 CLKS.n147 0.0371379
R5941 CLKS.n134 CLKS.n124 0.0371379
R5942 CLKS.n111 CLKS.n101 0.0371379
R5943 CLKS.n88 CLKS.n78 0.0371379
R5944 CLKS.n65 CLKS.n55 0.0371379
R5945 CLKS.n42 CLKS.n32 0.0371379
R5946 CLKS.n20 CLKS.n10 0.0371379
R5947 CLKS.n340 CLKS 0.03675
R5948 CLKS.n329 CLKS 0.03675
R5949 CLKS.n318 CLKS 0.03675
R5950 CLKS.n307 CLKS 0.03675
R5951 CLKS.n297 CLKS 0.03675
R5952 CLKS.n284 CLKS.n283 0.03675
R5953 CLKS.n276 CLKS.n275 0.03675
R5954 CLKS.n268 CLKS.n267 0.03675
R5955 CLKS.n260 CLKS.n259 0.03675
R5956 CLKS.n252 CLKS.n251 0.03675
R5957 CLKS.n341 CLKS.n340 0.0366675
R5958 CLKS.n330 CLKS.n329 0.0366675
R5959 CLKS.n319 CLKS.n318 0.0366675
R5960 CLKS.n308 CLKS.n307 0.0366675
R5961 CLKS.n298 CLKS.n297 0.0366675
R5962 CLKS.n284 CLKS 0.036656
R5963 CLKS.n276 CLKS 0.036656
R5964 CLKS.n268 CLKS 0.036656
R5965 CLKS.n260 CLKS 0.036656
R5966 CLKS.n252 CLKS 0.036656
R5967 CLKS.n210 CLKS 0.0222391
R5968 CLKS.n220 CLKS 0.0222391
R5969 CLKS.n187 CLKS 0.0222391
R5970 CLKS.n197 CLKS 0.0222391
R5971 CLKS.n164 CLKS 0.0222391
R5972 CLKS.n174 CLKS 0.0222391
R5973 CLKS.n141 CLKS 0.0222391
R5974 CLKS.n151 CLKS 0.0222391
R5975 CLKS.n118 CLKS 0.0222391
R5976 CLKS.n128 CLKS 0.0222391
R5977 CLKS.n95 CLKS 0.0222391
R5978 CLKS.n105 CLKS 0.0222391
R5979 CLKS.n72 CLKS 0.0222391
R5980 CLKS.n82 CLKS 0.0222391
R5981 CLKS.n49 CLKS 0.0222391
R5982 CLKS.n59 CLKS 0.0222391
R5983 CLKS.n26 CLKS 0.0222391
R5984 CLKS.n36 CLKS 0.0222391
R5985 CLKS.n4 CLKS 0.0222391
R5986 CLKS.n14 CLKS 0.0222391
R5987 CLKS CLKS.n214 0.0213333
R5988 CLKS CLKS.n225 0.0213333
R5989 CLKS CLKS.n191 0.0213333
R5990 CLKS CLKS.n202 0.0213333
R5991 CLKS CLKS.n168 0.0213333
R5992 CLKS CLKS.n179 0.0213333
R5993 CLKS CLKS.n145 0.0213333
R5994 CLKS CLKS.n156 0.0213333
R5995 CLKS CLKS.n122 0.0213333
R5996 CLKS CLKS.n133 0.0213333
R5997 CLKS CLKS.n99 0.0213333
R5998 CLKS CLKS.n110 0.0213333
R5999 CLKS CLKS.n76 0.0213333
R6000 CLKS CLKS.n87 0.0213333
R6001 CLKS CLKS.n53 0.0213333
R6002 CLKS CLKS.n64 0.0213333
R6003 CLKS CLKS.n30 0.0213333
R6004 CLKS CLKS.n41 0.0213333
R6005 CLKS CLKS.n8 0.0213333
R6006 CLKS CLKS.n19 0.0213333
R6007 CLKS.n221 CLKS.n220 0.00774638
R6008 CLKS.n198 CLKS.n197 0.00774638
R6009 CLKS.n175 CLKS.n174 0.00774638
R6010 CLKS.n152 CLKS.n151 0.00774638
R6011 CLKS.n129 CLKS.n128 0.00774638
R6012 CLKS.n106 CLKS.n105 0.00774638
R6013 CLKS.n83 CLKS.n82 0.00774638
R6014 CLKS.n60 CLKS.n59 0.00774638
R6015 CLKS.n37 CLKS.n36 0.00774638
R6016 CLKS.n15 CLKS.n14 0.00774638
R6017 CLKS CLKS.n341 0.00530769
R6018 CLKS CLKS.n330 0.00530769
R6019 CLKS CLKS.n319 0.00530769
R6020 CLKS CLKS.n308 0.00530769
R6021 CLKS CLKS.n298 0.00530769
R6022 CLKS.n288 CLKS.n287 0.00290385
R6023 CLKS.n280 CLKS.n279 0.00290385
R6024 CLKS.n272 CLKS.n271 0.00290385
R6025 CLKS.n264 CLKS.n263 0.00290385
R6026 CLKS.n256 CLKS.n255 0.00290385
R6027 a_n2715_n9662.t0 a_n2715_n9662.t1 60.0005
R6028 VSSD.n2012 VSSD.n3 9.88368e+06
R6029 VSSD VSSD.n2 2.17857e+06
R6030 VSSD.n207 VSSD.n3 2.0636e+06
R6031 VSSD.n3 VSSD.n2 1.9578e+06
R6032 VSSD VSSD.n207 386458
R6033 VSSD.n207 VSSD.t722 84628.4
R6034 VSSD.n1632 VSSD.n1631 46983.9
R6035 VSSD.n1629 VSSD.n1628 31723.6
R6036 VSSD.n2016 VSSD.n1 28119.8
R6037 VSSD.n2014 VSSD 13376.6
R6038 VSSD.n2014 VSSD.t639 12312.9
R6039 VSSD.n2016 VSSD.n2015 4622.73
R6040 VSSD.n1630 VSSD.n1629 4525.33
R6041 VSSD.n208 VSSD.t294 2823.12
R6042 VSSD.n1631 VSSD 2722.79
R6043 VSSD.t946 VSSD.t331 2161.85
R6044 VSSD.t66 VSSD.t641 2161.85
R6045 VSSD.t676 VSSD.t587 2161.85
R6046 VSSD.t785 VSSD.t427 2161.85
R6047 VSSD.t582 VSSD.t773 2161.85
R6048 VSSD.t1186 VSSD.t830 2161.85
R6049 VSSD.t897 VSSD.t24 2149.43
R6050 VSSD.t227 VSSD.t202 2149.43
R6051 VSSD.t570 VSSD.t436 2149.43
R6052 VSSD.t97 VSSD.t790 2149.43
R6053 VSSD.t899 VSSD.t28 2149.43
R6054 VSSD.t363 VSSD.t870 2149.43
R6055 VSSD.t30 VSSD.t59 2149.43
R6056 VSSD.t536 VSSD.t424 2149.43
R6057 VSSD.t625 VSSD.t521 2149.43
R6058 VSSD.t365 VSSD.t631 2149.43
R6059 VSSD.n1629 VSSD 2118.34
R6060 VSSD.n2015 VSSD.n2 2115.99
R6061 VSSD.t396 VSSD.n764 1932.95
R6062 VSSD.t1132 VSSD.t50 1763.39
R6063 VSSD.t390 VSSD.t223 1763.39
R6064 VSSD.t99 VSSD.t102 1763.39
R6065 VSSD.t770 VSSD.t749 1763.39
R6066 VSSD.t781 VSSD.t457 1763.39
R6067 VSSD.t462 VSSD.t504 1763.39
R6068 VSSD.t893 VSSD.t1147 1763.39
R6069 VSSD.t1160 VSSD.t290 1753.26
R6070 VSSD.t382 VSSD.t1161 1753.26
R6071 VSSD.t833 VSSD.t847 1753.26
R6072 VSSD.t814 VSSD.t96 1753.26
R6073 VSSD.t872 VSSD.t180 1753.26
R6074 VSSD.t989 VSSD.t996 1753.26
R6075 VSSD.t901 VSSD.t1138 1753.26
R6076 VSSD.t788 VSSD.t199 1753.26
R6077 VSSD.t953 VSSD.t217 1753.26
R6078 VSSD.t914 VSSD.t415 1753.26
R6079 VSSD.t798 VSSD.t519 1753.26
R6080 VSSD.t733 VSSD.t584 1753.26
R6081 VSSD.t564 VSSD.t243 1753.26
R6082 VSSD.t41 VSSD.t465 1753.26
R6083 VSSD.t585 VSSD.t68 1753.26
R6084 VSSD.t139 VSSD.t273 1753.26
R6085 VSSD.t87 VSSD.t380 1753.26
R6086 VSSD.t502 VSSD.t560 1753.26
R6087 VSSD.t288 VSSD.t756 1753.26
R6088 VSSD.t32 VSSD.t531 1753.26
R6089 VSSD.n1630 VSSD.n3 1690.5
R6090 VSSD VSSD.t351 1677.39
R6091 VSSD.n1631 VSSD.n1 1446.09
R6092 VSSD.t707 VSSD.t672 1407.32
R6093 VSSD.t1135 VSSD.t126 1407.32
R6094 VSSD.t445 VSSD.t528 1407.32
R6095 VSSD.t500 VSSD.t700 1407.32
R6096 VSSD.t319 VSSD.t956 1407.32
R6097 VSSD.t573 VSSD.t20 1407.32
R6098 VSSD.t361 VSSD.t238 1407.32
R6099 VSSD.t452 VSSD.t69 1399.23
R6100 VSSD.t505 VSSD.t443 1399.23
R6101 VSSD.t926 VSSD.t935 1399.23
R6102 VSSD.t538 VSSD.t444 1399.23
R6103 VSSD.t133 VSSD.t591 1399.23
R6104 VSSD.t272 VSSD.t590 1399.23
R6105 VSSD.t142 VSSD.t335 1399.23
R6106 VSSD.t464 VSSD.t614 1399.23
R6107 VSSD.t151 VSSD.t890 1399.23
R6108 VSSD.t320 VSSD.t135 1399.23
R6109 VSSD.t46 VSSD.t282 1263.2
R6110 VSSD.t221 VSSD.t1169 1263.2
R6111 VSSD.t1133 VSSD.t730 1263.2
R6112 VSSD.t747 VSSD.t697 1263.2
R6113 VSSD.t724 VSSD.t951 1263.2
R6114 VSSD.t1175 VSSD.t341 1263.2
R6115 VSSD.t1171 VSSD.t1130 1263.2
R6116 VSSD.t1018 VSSD.t498 1255.94
R6117 VSSD.t1012 VSSD.t303 1255.94
R6118 VSSD.t1039 VSSD.t566 1255.94
R6119 VSSD.t1058 VSSD.t578 1255.94
R6120 VSSD.t1061 VSSD.t801 1255.94
R6121 VSSD.t1006 VSSD.t137 1255.94
R6122 VSSD.t1035 VSSD.t127 1255.94
R6123 VSSD.t1024 VSSD.t77 1255.94
R6124 VSSD.t1078 VSSD.t286 1255.94
R6125 VSSD.t1026 VSSD.t7 1255.94
R6126 VSSD.n1 VSSD.t106 1180.08
R6127 VSSD.n2012 VSSD.n2011 1179.43
R6128 VSSD.n2018 VSSD.n2017 1170
R6129 VSSD.t186 VSSD.t908 1119.08
R6130 VSSD.t515 VSSD.t368 1119.08
R6131 VSSD.t689 VSSD.t359 1119.08
R6132 VSSD.t276 VSSD.t705 1119.08
R6133 VSSD.t315 VSSD.t1120 1119.08
R6134 VSSD.t298 VSSD.t268 1119.08
R6135 VSSD.t843 VSSD.t621 1119.08
R6136 VSSD.t344 VSSD.t1037 1112.64
R6137 VSSD.t840 VSSD.t1045 1112.64
R6138 VSSD.t678 VSSD.t1008 1112.64
R6139 VSSD.t178 VSSD.t1022 1112.64
R6140 VSSD.t493 VSSD.t1030 1112.64
R6141 VSSD.t388 VSSD.t1020 1112.64
R6142 VSSD.t34 VSSD.t1053 1112.64
R6143 VSSD.t834 VSSD.t1047 1112.64
R6144 VSSD.t404 VSSD.t1041 1112.64
R6145 VSSD.t85 VSSD.t1071 1112.64
R6146 VSSD.t48 VSSD 1110.6
R6147 VSSD.t225 VSSD 1110.6
R6148 VSSD.t100 VSSD 1110.6
R6149 VSSD.t483 VSSD 1110.6
R6150 VSSD VSSD.t779 1110.6
R6151 VSSD VSSD.t460 1110.6
R6152 VSSD VSSD.t891 1110.6
R6153 VSSD VSSD.t917 1104.21
R6154 VSSD VSSD.t602 1104.21
R6155 VSSD VSSD.t79 1104.21
R6156 VSSD VSSD.t959 1104.21
R6157 VSSD VSSD.t168 1104.21
R6158 VSSD VSSD.t89 1104.21
R6159 VSSD VSSD.t75 1104.21
R6160 VSSD VSSD.t684 1104.21
R6161 VSSD VSSD.t26 1104.21
R6162 VSSD.n1631 VSSD.n1630 1101.19
R6163 VSSD VSSD.n2012 962.422
R6164 VSSD.t708 VSSD.t669 924.086
R6165 VSSD.t592 VSSD.t948 924.086
R6166 VSSD.t446 VSSD.t317 924.086
R6167 VSSD.t501 VSSD.t1128 924.086
R6168 VSSD.t429 VSSD.t399 924.086
R6169 VSSD.t1194 VSSD.t21 924.086
R6170 VSSD.t832 VSSD.t239 924.086
R6171 VSSD.t22 VSSD.t70 918.774
R6172 VSSD.t200 VSSD.t744 918.774
R6173 VSSD.t149 VSSD.t534 918.774
R6174 VSSD.t839 VSSD.t589 918.774
R6175 VSSD.t601 VSSD.t95 918.774
R6176 VSSD.t285 VSSD.t775 918.774
R6177 VSSD.t61 VSSD.t157 918.774
R6178 VSSD.t426 VSSD.t615 918.774
R6179 VSSD.t520 VSSD.t889 918.774
R6180 VSSD.t630 VSSD.t787 918.774
R6181 VSSD.t908 VSSD.t708 839.307
R6182 VSSD.t368 VSSD.t592 839.307
R6183 VSSD.t359 VSSD.t446 839.307
R6184 VSSD.t705 VSSD.t501 839.307
R6185 VSSD.t399 VSSD.t315 839.307
R6186 VSSD.t21 VSSD.t298 839.307
R6187 VSSD.t239 VSSD.t843 839.307
R6188 VSSD.t70 VSSD.t344 834.484
R6189 VSSD.t744 VSSD.t840 834.484
R6190 VSSD.t534 VSSD.t678 834.484
R6191 VSSD.t589 VSSD.t178 834.484
R6192 VSSD.t95 VSSD.t493 834.484
R6193 VSSD.t775 VSSD.t388 834.484
R6194 VSSD.t157 VSSD.t34 834.484
R6195 VSSD.t615 VSSD.t834 834.484
R6196 VSSD.t889 VSSD.t404 834.484
R6197 VSSD.t787 VSSD.t85 834.484
R6198 VSSD.t669 VSSD.t46 813.874
R6199 VSSD.t670 VSSD.t707 813.874
R6200 VSSD.t948 VSSD.t221 813.874
R6201 VSSD.t1005 VSSD.t1135 813.874
R6202 VSSD.t317 VSSD.t1133 813.874
R6203 VSSD.t318 VSSD.t445 813.874
R6204 VSSD.t1128 VSSD.t747 813.874
R6205 VSSD.t675 VSSD.t500 813.874
R6206 VSSD.t951 VSSD.t429 813.874
R6207 VSSD.t956 VSSD.t535 813.874
R6208 VSSD.t341 VSSD.t1194 813.874
R6209 VSSD.t20 VSSD.t643 813.874
R6210 VSSD.t1130 VSSD.t832 813.874
R6211 VSSD.t238 VSSD.t829 813.874
R6212 VSSD.t668 VSSD.t393 809.196
R6213 VSSD.t969 VSSD.t665 809.196
R6214 VSSD.t386 VSSD.t1004 809.196
R6215 VSSD.t508 VSSD.t949 809.196
R6216 VSSD.t740 VSSD.t1180 809.196
R6217 VSSD.t328 VSSD.t849 809.196
R6218 VSSD.t818 VSSD.t1181 809.196
R6219 VSSD.t329 VSSD.t62 809.196
R6220 VSSD.t778 VSSD.t234 809.196
R6221 VSSD.t478 VSSD.t551 809.196
R6222 VSSD.t965 VSSD.t972 809.196
R6223 VSSD.t109 VSSD.t757 809.196
R6224 VSSD.t660 VSSD.t797 809.196
R6225 VSSD.t38 VSSD.t333 809.196
R6226 VSSD.t970 VSSD.t794 809.196
R6227 VSSD.t629 VSSD.t556 809.196
R6228 VSSD.t867 VSSD.t497 809.196
R6229 VSSD.t325 VSSD.t215 809.196
R6230 VSSD.t912 VSSD.t924 809.196
R6231 VSSD.t324 VSSD.t865 809.196
R6232 VSSD.t498 VSSD.t22 809.196
R6233 VSSD.t69 VSSD.t23 809.196
R6234 VSSD.t303 VSSD.t200 809.196
R6235 VSSD.t443 VSSD.t201 809.196
R6236 VSSD.t566 VSSD.t149 809.196
R6237 VSSD.t935 VSSD.t150 809.196
R6238 VSSD.t578 VSSD.t839 809.196
R6239 VSSD.t444 VSSD.t190 809.196
R6240 VSSD.t801 VSSD.t601 809.196
R6241 VSSD.t591 VSSD.t112 809.196
R6242 VSSD.t137 VSSD.t285 809.196
R6243 VSSD.t590 VSSD.t284 809.196
R6244 VSSD.t127 VSSD.t61 809.196
R6245 VSSD.t335 VSSD.t58 809.196
R6246 VSSD.t77 VSSD.t426 809.196
R6247 VSSD.t614 VSSD.t711 809.196
R6248 VSSD.t286 VSSD.t520 809.196
R6249 VSSD.t890 VSSD.t4 809.196
R6250 VSSD.t7 VSSD.t630 809.196
R6251 VSSD.t135 VSSD.t116 809.196
R6252 VSSD.t618 VSSD.t670 805.395
R6253 VSSD.t331 VSSD.t1005 805.395
R6254 VSSD.t641 VSSD.t318 805.395
R6255 VSSD.t587 VSSD.t675 805.395
R6256 VSSD.t535 VSSD.t785 805.395
R6257 VSSD.t643 VSSD.t582 805.395
R6258 VSSD.t829 VSSD.t1186 805.395
R6259 VSSD.t23 VSSD.t897 800.766
R6260 VSSD.t201 VSSD.t227 800.766
R6261 VSSD.t150 VSSD.t570 800.766
R6262 VSSD.t190 VSSD.t97 800.766
R6263 VSSD.t112 VSSD.t899 800.766
R6264 VSSD.t284 VSSD.t363 800.766
R6265 VSSD.t58 VSSD.t30 800.766
R6266 VSSD.t711 VSSD.t536 800.766
R6267 VSSD.t4 VSSD.t625 800.766
R6268 VSSD.t116 VSSD.t365 800.766
R6269 VSSD.t282 VSSD.t1132 771.485
R6270 VSSD.t1169 VSSD.t390 771.485
R6271 VSSD.t730 VSSD.t99 771.485
R6272 VSSD.t697 VSSD.t770 771.485
R6273 VSSD.t457 VSSD.t724 771.485
R6274 VSSD.t504 VSSD.t1175 771.485
R6275 VSSD.t1147 VSSD.t1171 771.485
R6276 VSSD.t519 VSSD.t1018 767.051
R6277 VSSD.t584 VSSD.t1012 767.051
R6278 VSSD.t243 VSSD.t1039 767.051
R6279 VSSD.t465 VSSD.t1058 767.051
R6280 VSSD.t68 VSSD.t1061 767.051
R6281 VSSD.t273 VSSD.t1006 767.051
R6282 VSSD.t380 VSSD.t1035 767.051
R6283 VSSD.t560 VSSD.t1024 767.051
R6284 VSSD.t756 VSSD.t1078 767.051
R6285 VSSD.t531 VSSD.t1026 767.051
R6286 VSSD.t474 VSSD.t396 712.139
R6287 VSSD.t50 VSSD.t48 712.139
R6288 VSSD.t223 VSSD.t225 712.139
R6289 VSSD.t307 VSSD.t946 712.139
R6290 VSSD.t102 VSSD.t100 712.139
R6291 VSSD.t882 VSSD.t66 712.139
R6292 VSSD.t749 VSSD.t483 712.139
R6293 VSSD.t779 VSSD.t781 712.139
R6294 VSSD.t427 VSSD.t558 712.139
R6295 VSSD.t460 VSSD.t462 712.139
R6296 VSSD.t773 VSSD.t309 712.139
R6297 VSSD.t891 VSSD.t893 712.139
R6298 VSSD.t830 VSSD.t468 712.139
R6299 VSSD.t106 VSSD.t798 708.047
R6300 VSSD.t24 VSSD.t256 708.047
R6301 VSSD.t917 VSSD.t733 708.047
R6302 VSSD.t202 VSSD.t523 708.047
R6303 VSSD.t602 VSSD.t564 708.047
R6304 VSSD.t436 VSSD.t229 708.047
R6305 VSSD.t79 VSSD.t41 708.047
R6306 VSSD.t790 VSSD.t123 708.047
R6307 VSSD.t959 VSSD.t585 708.047
R6308 VSSD.t28 VSSD.t447 708.047
R6309 VSSD.t168 VSSD.t139 708.047
R6310 VSSD.t870 VSSD.t2 708.047
R6311 VSSD.t89 VSSD.t87 708.047
R6312 VSSD.t59 VSSD.t654 708.047
R6313 VSSD.t75 VSSD.t502 708.047
R6314 VSSD.t424 VSSD.t673 708.047
R6315 VSSD.t684 VSSD.t288 708.047
R6316 VSSD.t521 VSSD.t81 708.047
R6317 VSSD.t26 VSSD.t32 708.047
R6318 VSSD.t631 VSSD.t370 708.047
R6319 VSSD.t351 VSSD.t349 708.047
R6320 VSSD.t349 VSSD.t248 708.047
R6321 VSSD.t248 VSSD.t246 708.047
R6322 VSSD.t246 VSSD.t193 708.047
R6323 VSSD.t193 VSSD.t191 708.047
R6324 VSSD.t191 VSSD.t172 708.047
R6325 VSSD.t172 VSSD.t170 708.047
R6326 VSSD.t170 VSSD.t258 708.047
R6327 VSSD.t258 VSSD.t418 708.047
R6328 VSSD.t418 VSSD.t260 708.047
R6329 VSSD.t391 VSSD.t292 640.614
R6330 VSSD.t400 VSSD.t1051 640.614
R6331 VSSD.t1093 VSSD.t91 640.614
R6332 VSSD.t384 VSSD.t509 640.614
R6333 VSSD.t561 VSSD.t845 640.614
R6334 VSSD.t39 VSSD.t1016 640.614
R6335 VSSD.t1069 VSSD.t540 640.614
R6336 VSSD.t816 VSSD.t682 640.614
R6337 VSSD.t232 VSSD.t553 640.614
R6338 VSSD.t195 VSSD.t1032 640.614
R6339 VSSD.t1076 VSSD.t701 640.614
R6340 VSSD.t991 VSSD.t110 640.614
R6341 VSSD.t795 VSSD.t1136 640.614
R6342 VSSD.t717 VSSD.t1101 640.614
R6343 VSSD.t1049 VSSD.t411 640.614
R6344 VSSD.t973 VSSD.t36 640.614
R6345 VSSD.t495 VSSD.t219 640.614
R6346 VSSD.t402 VSSD.t1056 640.614
R6347 VSSD.t1010 VSSD.t1002 640.614
R6348 VSSD.t910 VSSD.t326 640.614
R6349 VSSD.t672 VSSD.t186 610.405
R6350 VSSD.t126 VSSD.t515 610.405
R6351 VSSD.t528 VSSD.t689 610.405
R6352 VSSD.t700 VSSD.t276 610.405
R6353 VSSD.t1120 VSSD.t319 610.405
R6354 VSSD.t268 VSSD.t573 610.405
R6355 VSSD.t621 VSSD.t361 610.405
R6356 VSSD.t1037 VSSD.t452 606.898
R6357 VSSD.t1045 VSSD.t505 606.898
R6358 VSSD.t1008 VSSD.t926 606.898
R6359 VSSD.t1022 VSSD.t538 606.898
R6360 VSSD.t1030 VSSD.t133 606.898
R6361 VSSD.t1020 VSSD.t272 606.898
R6362 VSSD.t1053 VSSD.t142 606.898
R6363 VSSD.t1047 VSSD.t464 606.898
R6364 VSSD.t1041 VSSD.t151 606.898
R6365 VSSD.t1071 VSSD.t320 606.898
R6366 VSSD.n2017 VSSD 606.898
R6367 VSSD.n2013 VSSD 564.751
R6368 VSSD VSSD.t474 551.061
R6369 VSSD VSSD.t307 551.061
R6370 VSSD VSSD.t882 551.061
R6371 VSSD.t803 VSSD 551.061
R6372 VSSD.t558 VSSD 551.061
R6373 VSSD.t309 VSSD 551.061
R6374 VSSD.t468 VSSD 551.061
R6375 VSSD VSSD.t876 547.894
R6376 VSSD VSSD.t472 547.894
R6377 VSSD VSSD.t648 547.894
R6378 VSSD VSSD.t644 547.894
R6379 VSSD VSSD.t878 547.894
R6380 VSSD.t256 VSSD 547.894
R6381 VSSD.t523 VSSD 547.894
R6382 VSSD.t229 VSSD 547.894
R6383 VSSD.t123 VSSD 547.894
R6384 VSSD.t447 VSSD 547.894
R6385 VSSD.t2 VSSD 547.894
R6386 VSSD.t654 VSSD 547.894
R6387 VSSD.t673 VSSD 547.894
R6388 VSSD.t81 VSSD 547.894
R6389 VSSD.t370 VSSD 547.894
R6390 VSSD.t260 VSSD 539.465
R6391 VSSD.n765 VSSD.t618 536.793
R6392 VSSD.t297 VSSD.t969 505.748
R6393 VSSD.t1004 VSSD.t1143 505.748
R6394 VSSD.t530 VSSD.t328 505.748
R6395 VSSD.t1181 VSSD.t1154 505.748
R6396 VSSD.t864 VSSD.t478 505.748
R6397 VSSD.t972 VSSD.t244 505.748
R6398 VSSD.t761 VSSD.t38 505.748
R6399 VSSD.t794 VSSD.t134 505.748
R6400 VSSD.t712 VSSD.t325 505.748
R6401 VSSD.t924 VSSD.t807 505.748
R6402 VSSD VSSD.n765 474.589
R6403 VSSD.t91 VSSD.t400 472.031
R6404 VSSD.t540 VSSD.t39 472.031
R6405 VSSD.t701 VSSD.t195 472.031
R6406 VSSD.t411 VSSD.t717 472.031
R6407 VSSD.t1002 VSSD.t402 472.031
R6408 VSSD.n208 VSSD 457.803
R6409 VSSD.n2017 VSSD.n2016 446.743
R6410 VSSD.t1086 VSSD.t182 438.315
R6411 VSSD.t574 VSSD.t1088 438.315
R6412 VSSD.t1091 VSSD.t0 438.315
R6413 VSSD.t776 VSSD.t1063 438.315
R6414 VSSD.t1067 VSSD.t656 438.315
R6415 VSSD.t525 VSSD.t1043 438.315
R6416 VSSD.t1104 VSSD.t544 438.315
R6417 VSSD.t254 VSSD.t1107 438.315
R6418 VSSD.t1109 VSSD.t83 438.315
R6419 VSSD.t11 VSSD.t1083 438.315
R6420 VSSD.t950 VSSD.t297 413.027
R6421 VSSD.t1143 VSSD.t667 413.027
R6422 VSSD.t539 VSSD.t530 413.027
R6423 VSSD.t1154 VSSD.t863 413.027
R6424 VSSD.t758 VSSD.t864 413.027
R6425 VSSD.t244 VSSD.t995 413.027
R6426 VSSD.t557 VSSD.t761 413.027
R6427 VSSD.t134 VSSD.t659 413.027
R6428 VSSD.t866 VSSD.t712 413.027
R6429 VSSD.t807 VSSD.t927 413.027
R6430 VSSD.n209 VSSD.t803 373.026
R6431 VSSD.t393 VSSD.t1086 362.452
R6432 VSSD.t1088 VSSD.t508 362.452
R6433 VSSD.t1180 VSSD.t1091 362.452
R6434 VSSD.t1063 VSSD.t329 362.452
R6435 VSSD.t234 VSSD.t1067 362.452
R6436 VSSD.t1043 VSSD.t109 362.452
R6437 VSSD.t797 VSSD.t1104 362.452
R6438 VSSD.t1107 VSSD.t629 362.452
R6439 VSSD.t497 VSSD.t1109 362.452
R6440 VSSD.t1083 VSSD.t324 362.452
R6441 VSSD.t768 VSSD.t409 352.166
R6442 VSSD.t979 VSSD.t491 352.166
R6443 VSSD.t633 VSSD.t931 352.166
R6444 VSSD.t44 VSSD.t438 352.166
R6445 VSSD.t886 VSSD.t64 352.166
R6446 VSSD.n209 VSSD.t676 339.115
R6447 VSSD.t874 VSSD.t751 330.07
R6448 VSSD.t182 VSSD.t1160 328.736
R6449 VSSD.t1161 VSSD.t574 328.736
R6450 VSSD.t0 VSSD.t833 328.736
R6451 VSSD.t96 VSSD.t776 328.736
R6452 VSSD.t656 VSSD.t872 328.736
R6453 VSSD.t996 VSSD.t525 328.736
R6454 VSSD.t544 VSSD.t901 328.736
R6455 VSSD.t199 VSSD.t254 328.736
R6456 VSSD.t83 VSSD.t953 328.736
R6457 VSSD.t415 VSSD.t11 328.736
R6458 VSSD.t117 VSSD.t235 327.591
R6459 VSSD.t1118 VSSD.t322 327.591
R6460 VSSD.t687 VSSD.t441 327.591
R6461 VSSD.t420 VSSD.t982 317.039
R6462 VSSD.t765 VSSD.t652 317.039
R6463 VSSD.t453 VSSD.t104 317.039
R6464 VSSD.t920 VSSD.t1152 317.039
R6465 VSSD.t933 VSSD.t975 317.039
R6466 VSSD.n1648 VSSD.t983 307.536
R6467 VSSD.n1681 VSSD.t653 307.536
R6468 VSSD.n1719 VSSD.t105 307.536
R6469 VSSD.n1752 VSSD.t1153 307.536
R6470 VSSD.n1790 VSSD.t976 307.536
R6471 VSSD.n1450 VSSD.t887 307.536
R6472 VSSD.n1434 VSSD.t45 307.536
R6473 VSSD.n1522 VSSD.t634 307.536
R6474 VSSD.n1556 VSSD.t980 307.536
R6475 VSSD.n1399 VSSD.t769 307.536
R6476 VSSD.n100 VSSD.t12 307.536
R6477 VSSD.n1881 VSSD.t84 307.536
R6478 VSSD.n2007 VSSD.t183 307.536
R6479 VSSD.n20 VSSD.t575 307.536
R6480 VSSD.n1976 VSSD.t1 307.536
R6481 VSSD.n41 VSSD.t777 307.536
R6482 VSSD.n1945 VSSD.t657 307.536
R6483 VSSD.n62 VSSD.t526 307.536
R6484 VSSD.n1914 VSSD.t545 307.536
R6485 VSSD.n83 VSSD.t255 307.536
R6486 VSSD.n438 VSSD.t332 307.536
R6487 VSSD.n403 VSSD.t642 307.536
R6488 VSSD.n368 VSSD.t588 307.536
R6489 VSSD.n333 VSSD.t786 307.536
R6490 VSSD.n298 VSSD.t583 307.536
R6491 VSSD.n263 VSSD.t1187 307.536
R6492 VSSD.n526 VSSD.t118 307.536
R6493 VSSD.n564 VSSD.t1119 307.536
R6494 VSSD.n604 VSSD.t688 307.536
R6495 VSSD.n731 VSSD.t968 307.536
R6496 VSSD.n696 VSSD.t619 307.536
R6497 VSSD.n661 VSSD.t613 307.536
R6498 VSSD.n1299 VSSD.t366 307.536
R6499 VSSD.n1299 VSSD.t568 307.536
R6500 VSSD.n1264 VSSD.t896 307.536
R6501 VSSD.n1264 VSSD.t626 307.536
R6502 VSSD.n1229 VSSD.t537 307.536
R6503 VSSD.n1229 VSSD.t812 307.536
R6504 VSSD.n1194 VSSD.t31 307.536
R6505 VSSD.n1194 VSSD.t813 307.536
R6506 VSSD.n1159 VSSD.t364 307.536
R6507 VSSD.n1159 VSSD.t885 307.536
R6508 VSSD.n1124 VSSD.t900 307.536
R6509 VSSD.n1124 VSSD.t937 307.536
R6510 VSSD.n1089 VSSD.t98 307.536
R6511 VSSD.n1089 VSSD.t569 307.536
R6512 VSSD.n1054 VSSD.t1192 307.536
R6513 VSSD.n1054 VSSD.t571 307.536
R6514 VSSD.n1019 VSSD.t228 307.536
R6515 VSSD.n1019 VSSD.t884 307.536
R6516 VSSD.n984 VSSD.t898 307.536
R6517 VSSD.n984 VSSD.t936 307.536
R6518 VSSD.n764 VSSD.t1014 304.682
R6519 VSSD.t481 VSSD.t242 287.257
R6520 VSSD.t264 VSSD.t343 287.257
R6521 VSSD.t434 VSSD.t837 287.257
R6522 VSSD.t598 VSSD.t988 287.257
R6523 VSSD.t313 VSSD.t764 287.257
R6524 VSSD.n119 VSSD.t163 282.885
R6525 VSSD.n777 VSSD.t120 282.327
R6526 VSSD.n118 VSSD.t175 281.13
R6527 VSSD.n473 VSSD.t161 280.457
R6528 VSSD.t357 VSSD.t555 267.212
R6529 VSSD.t55 VSSD.t627 267.212
R6530 VSSD.t152 VSSD.t296 267.212
R6531 VSSD.t529 VSSD.t808 267.212
R6532 VSSD.t650 VSSD 261.303
R6533 VSSD.t646 VSSD 261.303
R6534 VSSD.t822 VSSD 261.303
R6535 VSSD.t305 VSSD 261.303
R6536 VSSD.t470 VSSD 261.303
R6537 VSSD.t155 VSSD.t143 258.604
R6538 VSSD.t214 VSSD.t906 258.604
R6539 VSSD.t593 VSSD.t663 258.604
R6540 VSSD.t940 VSSD.t252 258.604
R6541 VSSD.t628 VSSD.t635 258.604
R6542 VSSD.t455 VSSD 248.659
R6543 VSSD VSSD.t160 241.702
R6544 VSSD.n1675 VSSD.t146 238.083
R6545 VSSD.n1360 VSSD.t903 238.083
R6546 VSSD.n1746 VSSD.t662 238.083
R6547 VSSD.n1337 VSSD.t714 238.083
R6548 VSSD.n1817 VSSD.t640 238.083
R6549 VSSD.n1436 VSSD.t312 238.083
R6550 VSSD.n1515 VSSD.t595 238.083
R6551 VSSD.n1549 VSSD.t433 238.083
R6552 VSSD.n1401 VSSD.t263 238.083
R6553 VSSD.n1621 VSSD.t752 238.083
R6554 VSSD.n1851 VSSD.t911 238.083
R6555 VSSD.n2010 VSSD.t293 238.083
R6556 VSSD.n1980 VSSD.t385 238.083
R6557 VSSD.n1979 VSSD.t846 238.083
R6558 VSSD.n1949 VSSD.t817 238.083
R6559 VSSD.n1948 VSSD.t554 238.083
R6560 VSSD.n1918 VSSD.t992 238.083
R6561 VSSD.n1917 VSSD.t1137 238.083
R6562 VSSD.n1887 VSSD.t974 238.083
R6563 VSSD.n1886 VSSD.t220 238.083
R6564 VSSD.n1270 VSSD.t154 238.083
R6565 VSSD.n1270 VSSD.t27 238.083
R6566 VSSD.n1235 VSSD.t685 238.083
R6567 VSSD.n1235 VSSD.t873 238.083
R6568 VSSD.n1200 VSSD.t1113 238.083
R6569 VSSD.n1200 VSSD.t76 238.083
R6570 VSSD.n1165 VSSD.t90 238.083
R6571 VSSD.n1165 VSSD.t130 238.083
R6572 VSSD.n1130 VSSD.t198 238.083
R6573 VSSD.n1130 VSSD.t169 238.083
R6574 VSSD.n1095 VSSD.t1179 238.083
R6575 VSSD.n1095 VSSD.t960 238.083
R6576 VSSD.n1060 VSSD.t1148 238.083
R6577 VSSD.n1060 VSSD.t80 238.083
R6578 VSSD.n1025 VSSD.t603 238.083
R6579 VSSD.n1025 VSSD.t754 238.083
R6580 VSSD.n990 VSSD.t918 238.083
R6581 VSSD.n990 VSSD.t1151 238.083
R6582 VSSD.n956 VSSD.t1140 238.083
R6583 VSSD.n956 VSSD.t107 238.083
R6584 VSSD.n161 VSSD.t226 233.732
R6585 VSSD.n178 VSSD.t101 233.732
R6586 VSSD.n194 VSSD.t484 233.732
R6587 VSSD.n213 VSSD.t780 233.732
R6588 VSSD.n229 VSSD.t461 233.732
R6589 VSSD.n245 VSSD.t892 233.732
R6590 VSSD.n159 VSSD.t723 233.732
R6591 VSSD.n535 VSSD.t54 233.732
R6592 VSSD.n135 VSSD.t407 233.732
R6593 VSSD.n123 VSSD.t251 233.732
R6594 VSSD.n627 VSSD.t49 233.732
R6595 VSSD.n643 VSSD.t1163 233.732
R6596 VSSD.t108 VSSD.t577 229.254
R6597 VSSD.t330 VSSD.t1166 229.254
R6598 VSSD.t93 VSSD.t737 229.254
R6599 VSSD.t197 VSSD.t451 229.254
R6600 VSSD.t888 VSSD.t563 229.254
R6601 VSSD.n1673 VSSD.t144 226.882
R6602 VSSD.n1708 VSSD.t907 226.882
R6603 VSSD.n1744 VSSD.t664 226.882
R6604 VSSD.n1779 VSSD.t253 226.882
R6605 VSSD.n1815 VSSD.t636 226.882
R6606 VSSD.n1477 VSSD.t314 226.882
R6607 VSSD.n1511 VSSD.t599 226.882
R6608 VSSD.n1547 VSSD.t435 226.882
R6609 VSSD.n1583 VSSD.t265 226.882
R6610 VSSD.n1617 VSSD.t482 226.882
R6611 VSSD.n1854 VSSD.t915 226.882
R6612 VSSD.n88 VSSD.t218 226.882
R6613 VSSD.n2008 VSSD.t291 226.882
R6614 VSSD.n1982 VSSD.t383 226.882
R6615 VSSD.n1977 VSSD.t848 226.882
R6616 VSSD.n1951 VSSD.t815 226.882
R6617 VSSD.n1946 VSSD.t181 226.882
R6618 VSSD.n1920 VSSD.t990 226.882
R6619 VSSD.n1915 VSSD.t1139 226.882
R6620 VSSD.n1889 VSSD.t789 226.882
R6621 VSSD.n1272 VSSD.t964 226.882
R6622 VSSD.n1272 VSSD.t33 226.882
R6623 VSSD.n1237 VSSD.t348 226.882
R6624 VSSD.n1237 VSSD.t289 226.882
R6625 VSSD.n1202 VSSD.t503 226.882
R6626 VSSD.n1202 VSSD.t686 226.882
R6627 VSSD.n1167 VSSD.t88 226.882
R6628 VSSD.n1167 VSSD.t129 226.882
R6629 VSSD.n1132 VSSD.t736 226.882
R6630 VSSD.n1132 VSSD.t140 226.882
R6631 VSSD.n1097 VSSD.t586 226.882
R6632 VSSD.n1097 VSSD.t958 226.882
R6633 VSSD.n1062 VSSD.t42 226.882
R6634 VSSD.n1062 VSSD.t620 226.882
R6635 VSSD.n1027 VSSD.t565 226.882
R6636 VSSD.n1027 VSSD.t755 226.882
R6637 VSSD.n992 VSSD.t734 226.882
R6638 VSSD.n992 VSSD.t1150 226.882
R6639 VSSD.n957 VSSD.t1141 226.882
R6640 VSSD.n957 VSSD.t799 226.882
R6641 VSSD VSSD.t174 226.383
R6642 VSSD.n464 VSSD.t224 223.315
R6643 VSSD.n429 VSSD.t103 223.315
R6644 VSSD.n394 VSSD.t750 223.315
R6645 VSSD.n359 VSSD.t782 223.315
R6646 VSSD.n324 VSSD.t463 223.315
R6647 VSSD.n289 VSSD.t894 223.315
R6648 VSSD.n499 VSSD.t358 223.315
R6649 VSSD.n537 VSSD.t56 223.315
R6650 VSSD.n577 VSSD.t153 223.315
R6651 VSSD.n757 VSSD.t809 223.315
R6652 VSSD.n722 VSSD.t51 223.315
R6653 VSSD.n687 VSSD.t185 223.315
R6654 VSSD.t981 VSSD.t338 213.256
R6655 VSSD.t156 VSSD.t6 213.256
R6656 VSSD.t741 VSSD.t771 213.256
R6657 VSSD.t300 VSSD.t367 213.256
R6658 VSSD VSSD.t616 212.767
R6659 VSSD.n2013 VSSD 210.728
R6660 VSSD.n1667 VSSD.n1666 209.254
R6661 VSSD.n1702 VSSD.n1701 209.254
R6662 VSSD.n1738 VSSD.n1737 209.254
R6663 VSSD.n1773 VSSD.n1772 209.254
R6664 VSSD.n1809 VSSD.n1808 209.254
R6665 VSSD.n1471 VSSD.n1470 209.254
R6666 VSSD.n1429 VSSD.n1428 209.254
R6667 VSSD.n1541 VSSD.n1540 209.254
R6668 VSSD.n1577 VSSD.n1576 209.254
R6669 VSSD.n1394 VSSD.n1393 209.254
R6670 VSSD.n1861 VSSD.n1860 209.254
R6671 VSSD.n92 VSSD.n91 209.254
R6672 VSSD.n11 VSSD.n10 209.254
R6673 VSSD.n1988 VSSD.n19 209.254
R6674 VSSD.n32 VSSD.n31 209.254
R6675 VSSD.n1957 VSSD.n40 209.254
R6676 VSSD.n53 VSSD.n52 209.254
R6677 VSSD.n1926 VSSD.n61 209.254
R6678 VSSD.n74 VSSD.n73 209.254
R6679 VSSD.n1895 VSSD.n82 209.254
R6680 VSSD.n1278 VSSD.n818 209.254
R6681 VSSD.n1278 VSSD.n819 209.254
R6682 VSSD.n1243 VSSD.n833 209.254
R6683 VSSD.n1243 VSSD.n834 209.254
R6684 VSSD.n1208 VSSD.n848 209.254
R6685 VSSD.n1208 VSSD.n849 209.254
R6686 VSSD.n1173 VSSD.n863 209.254
R6687 VSSD.n1173 VSSD.n864 209.254
R6688 VSSD.n1138 VSSD.n878 209.254
R6689 VSSD.n1138 VSSD.n879 209.254
R6690 VSSD.n1103 VSSD.n893 209.254
R6691 VSSD.n1103 VSSD.n894 209.254
R6692 VSSD.n1068 VSSD.n908 209.254
R6693 VSSD.n1068 VSSD.n909 209.254
R6694 VSSD.n1033 VSSD.n923 209.254
R6695 VSSD.n1033 VSSD.n924 209.254
R6696 VSSD.n998 VSSD.n938 209.254
R6697 VSSD.n998 VSSD.n939 209.254
R6698 VSSD.n963 VSSD.n953 209.254
R6699 VSSD.n963 VSSD.n954 209.254
R6700 VSSD.n776 VSSD.n117 207.213
R6701 VSSD.n486 VSSD.n475 207.213
R6702 VSSD.n477 VSSD.n476 207.213
R6703 VSSD.n480 VSSD.n479 207.213
R6704 VSSD.t699 VSSD.t43 206.387
R6705 VSSD.t938 VSSD.t767 206.387
R6706 VSSD.t704 VSSD.t703 206.387
R6707 VSSD.t842 VSSD.t52 206.387
R6708 VSSD.t746 VSSD.t783 206.387
R6709 VSSD.t1000 VSSD.t479 205.775
R6710 VSSD.t517 VSSD.t532 205.775
R6711 VSSD.t1167 VSSD.t430 205.775
R6712 VSSD.t280 VSSD.t596 205.775
R6713 VSSD.t166 VSSD.t868 205.775
R6714 VSSD.t145 VSSD 205.143
R6715 VSSD.t902 VSSD 205.143
R6716 VSSD.t661 VSSD 205.143
R6717 VSSD.t713 VSSD 205.143
R6718 VSSD.n1637 VSSD.n1636 204.457
R6719 VSSD.n1388 VSSD.n1387 204.457
R6720 VSSD.n457 VSSD.n165 203.526
R6721 VSSD.n422 VSSD.n181 203.526
R6722 VSSD.n387 VSSD.n197 203.526
R6723 VSSD.n352 VSSD.n216 203.526
R6724 VSSD.n317 VSSD.n232 203.526
R6725 VSSD.n282 VSSD.n248 203.526
R6726 VSSD.n506 VSSD.n156 203.526
R6727 VSSD.n544 VSSD.n144 203.526
R6728 VSSD.n584 VSSD.n132 203.526
R6729 VSSD.n750 VSSD.n614 203.526
R6730 VSSD.n715 VSSD.n630 203.526
R6731 VSSD.n680 VSSD.n646 203.526
R6732 VSSD.n449 VSSD.n168 202.843
R6733 VSSD.n414 VSSD.n184 202.843
R6734 VSSD.n379 VSSD.n200 202.843
R6735 VSSD.n344 VSSD.n219 202.843
R6736 VSSD.n309 VSSD.n235 202.843
R6737 VSSD.n274 VSSD.n251 202.843
R6738 VSSD.n515 VSSD.n514 202.843
R6739 VSSD.n552 VSSD.n551 202.843
R6740 VSSD.n593 VSSD.n592 202.843
R6741 VSSD.n742 VSSD.n617 202.843
R6742 VSSD.n707 VSSD.n633 202.843
R6743 VSSD.n672 VSSD.n649 202.843
R6744 VSSD.n109 VSSD.n108 200.516
R6745 VSSD.n1837 VSSD.n1836 200.516
R6746 VSSD.n107 VSSD.n106 200.516
R6747 VSSD.n1844 VSSD.n1843 200.516
R6748 VSSD.n1847 VSSD.n1846 200.516
R6749 VSSD.n1320 VSSD.n792 200.516
R6750 VSSD.n1320 VSSD.n793 200.516
R6751 VSSD.n1318 VSSD.n794 200.516
R6752 VSSD.n1318 VSSD.n796 200.516
R6753 VSSD.n799 VSSD.n797 200.516
R6754 VSSD.n799 VSSD.n798 200.516
R6755 VSSD.n1312 VSSD.n801 200.516
R6756 VSSD.n1312 VSSD.n802 200.516
R6757 VSSD.n805 VSSD.n803 200.516
R6758 VSSD.n805 VSSD.n804 200.516
R6759 VSSD.n1644 VSSD.n1643 199.739
R6760 VSSD.n1378 VSSD.n1377 199.739
R6761 VSSD.n1679 VSSD.n1371 199.739
R6762 VSSD.n1693 VSSD.n1692 199.739
R6763 VSSD.n1715 VSSD.n1714 199.739
R6764 VSSD.n1355 VSSD.n1354 199.739
R6765 VSSD.n1750 VSSD.n1348 199.739
R6766 VSSD.n1764 VSSD.n1763 199.739
R6767 VSSD.n1786 VSSD.n1785 199.739
R6768 VSSD.n1332 VSSD.n1331 199.739
R6769 VSSD.n1448 VSSD.n1447 199.739
R6770 VSSD.n1462 VSSD.n1461 199.739
R6771 VSSD.n1484 VSSD.n1483 199.739
R6772 VSSD.n1498 VSSD.n1497 199.739
R6773 VSSD.n1518 VSSD.n1517 199.739
R6774 VSSD.n1418 VSSD.n1417 199.739
R6775 VSSD.n1554 VSSD.n1553 199.739
R6776 VSSD.n1568 VSSD.n1567 199.739
R6777 VSSD.n1590 VSSD.n1589 199.739
R6778 VSSD.n1604 VSSD.n1603 199.739
R6779 VSSD.n1853 VSSD.n1852 199.739
R6780 VSSD.n1869 VSSD.n1868 199.739
R6781 VSSD.n97 VSSD.n96 199.739
R6782 VSSD.n2009 VSSD.n5 199.739
R6783 VSSD.n15 VSSD.n14 199.739
R6784 VSSD.n1995 VSSD.n16 199.739
R6785 VSSD.n1981 VSSD.n22 199.739
R6786 VSSD.n1978 VSSD.n26 199.739
R6787 VSSD.n36 VSSD.n35 199.739
R6788 VSSD.n1964 VSSD.n37 199.739
R6789 VSSD.n1950 VSSD.n43 199.739
R6790 VSSD.n1947 VSSD.n47 199.739
R6791 VSSD.n57 VSSD.n56 199.739
R6792 VSSD.n1933 VSSD.n58 199.739
R6793 VSSD.n1919 VSSD.n64 199.739
R6794 VSSD.n1916 VSSD.n68 199.739
R6795 VSSD.n78 VSSD.n77 199.739
R6796 VSSD.n1902 VSSD.n79 199.739
R6797 VSSD.n1888 VSSD.n85 199.739
R6798 VSSD.n1885 VSSD.n89 199.739
R6799 VSSD.n174 VSSD.n173 199.739
R6800 VSSD.n190 VSSD.n189 199.739
R6801 VSSD.n206 VSSD.n205 199.739
R6802 VSSD.n225 VSSD.n224 199.739
R6803 VSSD.n241 VSSD.n240 199.739
R6804 VSSD.n257 VSSD.n256 199.739
R6805 VSSD.n530 VSSD.n149 199.739
R6806 VSSD.n569 VSSD.n568 199.739
R6807 VSSD.n608 VSSD.n125 199.739
R6808 VSSD.n623 VSSD.n622 199.739
R6809 VSSD.n639 VSSD.n638 199.739
R6810 VSSD.n655 VSSD.n654 199.739
R6811 VSSD.n1301 VSSD.n809 199.739
R6812 VSSD.n1301 VSSD.n810 199.739
R6813 VSSD.n1287 VSSD.n1285 199.739
R6814 VSSD.n1287 VSSD.n1286 199.739
R6815 VSSD.n825 VSSD.n823 199.739
R6816 VSSD.n825 VSSD.n824 199.739
R6817 VSSD.n1252 VSSD.n1250 199.739
R6818 VSSD.n1252 VSSD.n1251 199.739
R6819 VSSD.n840 VSSD.n838 199.739
R6820 VSSD.n840 VSSD.n839 199.739
R6821 VSSD.n1217 VSSD.n1215 199.739
R6822 VSSD.n1217 VSSD.n1216 199.739
R6823 VSSD.n855 VSSD.n853 199.739
R6824 VSSD.n855 VSSD.n854 199.739
R6825 VSSD.n1182 VSSD.n1180 199.739
R6826 VSSD.n1182 VSSD.n1181 199.739
R6827 VSSD.n870 VSSD.n868 199.739
R6828 VSSD.n870 VSSD.n869 199.739
R6829 VSSD.n1147 VSSD.n1145 199.739
R6830 VSSD.n1147 VSSD.n1146 199.739
R6831 VSSD.n885 VSSD.n883 199.739
R6832 VSSD.n885 VSSD.n884 199.739
R6833 VSSD.n1112 VSSD.n1110 199.739
R6834 VSSD.n1112 VSSD.n1111 199.739
R6835 VSSD.n900 VSSD.n898 199.739
R6836 VSSD.n900 VSSD.n899 199.739
R6837 VSSD.n1077 VSSD.n1075 199.739
R6838 VSSD.n1077 VSSD.n1076 199.739
R6839 VSSD.n915 VSSD.n913 199.739
R6840 VSSD.n915 VSSD.n914 199.739
R6841 VSSD.n1042 VSSD.n1040 199.739
R6842 VSSD.n1042 VSSD.n1041 199.739
R6843 VSSD.n930 VSSD.n928 199.739
R6844 VSSD.n930 VSSD.n929 199.739
R6845 VSSD.n1007 VSSD.n1005 199.739
R6846 VSSD.n1007 VSSD.n1006 199.739
R6847 VSSD.n945 VSSD.n943 199.739
R6848 VSSD.n945 VSSD.n944 199.739
R6849 VSSD.n972 VSSD.n970 199.739
R6850 VSSD.n972 VSSD.n971 199.739
R6851 VSSD.t1051 VSSD.t950 193.87
R6852 VSSD.t667 VSSD.t1093 193.87
R6853 VSSD.t1016 VSSD.t539 193.87
R6854 VSSD.t863 VSSD.t1069 193.87
R6855 VSSD.t1032 VSSD.t758 193.87
R6856 VSSD.t995 VSSD.t1076 193.87
R6857 VSSD.t1101 VSSD.t557 193.87
R6858 VSSD.t659 VSSD.t1049 193.87
R6859 VSSD.t1056 VSSD.t866 193.87
R6860 VSSD.t927 VSSD.t1010 193.87
R6861 VSSD.t691 VSSD.t355 191.417
R6862 VSSD.t278 VSSD.t580 191.417
R6863 VSSD.t1122 VSSD.t114 191.417
R6864 VSSD.t810 VSSD.t695 191.417
R6865 VSSD.t147 VSSD.t623 185.25
R6866 VSSD.t904 VSSD.t13 185.25
R6867 VSSD.t131 VSSD.t998 185.25
R6868 VSSD.t715 VSSD.t1126 185.25
R6869 VSSD.t637 VSSD.t274 185.25
R6870 VSSD.t476 VSSD.t188 182.298
R6871 VSSD.t487 VSSD.t1173 182.298
R6872 VSSD.t301 VSSD.t9 182.298
R6873 VSSD.t176 VSSD.t693 182.298
R6874 VSSD.t709 VSSD.t164 182.298
R6875 VSSD VSSD.t262 180.917
R6876 VSSD VSSD.t432 180.917
R6877 VSSD VSSD.t594 180.917
R6878 VSSD VSSD.t311 180.917
R6879 VSSD.t1014 VSSD 180.427
R6880 VSSD.t861 VSSD.t15 169.577
R6881 VSSD.t18 VSSD.t513 169.577
R6882 VSSD.t680 VSSD.t826 169.577
R6883 VSSD.t942 VSSD.t928 169.577
R6884 VSSD VSSD.t53 168.292
R6885 VSSD VSSD.t406 168.292
R6886 VSSD.t162 VSSD 166.81
R6887 VSSD.t270 VSSD.t240 164.114
R6888 VSSD.t266 VSSD.t485 164.114
R6889 VSSD.t511 VSSD.t605 164.114
R6890 VSSD.t726 VSSD.t1144 164.114
R6891 VSSD.t728 VSSD.t610 164.114
R6892 VSSD.n783 VSSD.t617 157.291
R6893 VSSD.n785 VSSD.t507 155.286
R6894 VSSD.n160 VSSD.t295 153.631
R6895 VSSD.n472 VSSD.t1015 153.631
R6896 VSSD.t408 VSSD.t763 150.535
R6897 VSSD.t490 VSSD.t576 150.535
R6898 VSSD.t94 VSSD.t738 150.535
R6899 VSSD.t1112 VSSD.t450 150.535
R6900 VSSD.t954 VSSD.t977 150.535
R6901 VSSD.n1830 VSSD.t856 149.762
R6902 VSSD.n1306 VSSD.t352 149.762
R6903 VSSD.n1306 VSSD.t721 149.762
R6904 VSSD.t1080 VSSD.t874 149.154
R6905 VSSD.t160 VSSD.t210 142.98
R6906 VSSD.t210 VSSD.t1182 142.98
R6907 VSSD.t1182 VSSD.t158 142.98
R6908 VSSD.t158 VSSD.t1184 142.98
R6909 VSSD.t1184 VSSD.t212 142.98
R6910 VSSD.t212 VSSD.t413 142.98
R6911 VSSD.t174 VSSD.t792 142.98
R6912 VSSD.t792 VSSD.t121 142.98
R6913 VSSD.t121 VSSD.t119 142.98
R6914 VSSD.t616 VSSD.t506 142.98
R6915 VSSD.t237 VSSD.t337 140.03
R6916 VSSD.t17 VSSD.t57 140.03
R6917 VSSD.t416 VSSD.t772 140.03
R6918 VSSD.t362 VSSD.t671 140.03
R6919 VSSD.t763 VSSD.t476 136.724
R6920 VSSD.t576 VSSD.t487 136.724
R6921 VSSD.t738 VSSD.t301 136.724
R6922 VSSD.t450 VSSD.t176 136.724
R6923 VSSD.t977 VSSD.t709 136.724
R6924 VSSD.t141 VSSD.t423 135.519
R6925 VSSD.t939 VSSD.t609 135.519
R6926 VSSD.t784 VSSD.t394 135.519
R6927 VSSD.t1178 VSSD.t919 135.519
R6928 VSSD.t745 VSSD.t993 135.519
R6929 VSSD.t1028 VSSD.t455 134.275
R6930 VSSD.t479 VSSD.t408 132.581
R6931 VSSD.t577 VSSD.t719 132.581
R6932 VSSD.t532 VSSD.t490 132.581
R6933 VSSD.t1166 VSSD.t604 132.581
R6934 VSSD.t430 VSSD.t94 132.581
R6935 VSSD.t737 VSSD.t374 132.581
R6936 VSSD.t596 VSSD.t1112 132.581
R6937 VSSD.t451 VSSD.t440 132.581
R6938 VSSD.t868 VSSD.t954 132.581
R6939 VSSD.t563 VSSD.t955 132.581
R6940 VSSD.t719 VSSD.t768 131.2
R6941 VSSD.t604 VSSD.t979 131.2
R6942 VSSD.t374 VSSD.t633 131.2
R6943 VSSD.t440 VSSD.t44 131.2
R6944 VSSD.t955 VSSD.t886 131.2
R6945 VSSD.t250 VSSD.n763 131.036
R6946 VSSD.t119 VSSD 127.66
R6947 VSSD.t337 VSSD.t861 127.183
R6948 VSSD.t57 VSSD.t18 127.183
R6949 VSSD.t772 VSSD.t680 127.183
R6950 VSSD.t928 VSSD.t362 127.183
R6951 VSSD.n2013 VSSD 125.898
R6952 VSSD.t242 VSSD.t1000 125.675
R6953 VSSD.t343 VSSD.t517 125.675
R6954 VSSD.t837 VSSD.t1167 125.675
R6955 VSSD.t988 VSSD.t280 125.675
R6956 VSSD.t764 VSSD.t166 125.675
R6957 VSSD.t355 VSSD.t237 123.329
R6958 VSSD.t338 VSSD.t923 123.329
R6959 VSSD.t580 VSSD.t17 123.329
R6960 VSSD.t6 VSSD.t321 123.329
R6961 VSSD.t114 VSSD.t416 123.329
R6962 VSSD.t771 VSSD.t417 123.329
R6963 VSSD.t671 VSSD.t810 123.329
R6964 VSSD.t395 VSSD.t300 123.329
R6965 VSSD.t240 VSSD.t141 123.087
R6966 VSSD.t485 VSSD.t939 123.087
R6967 VSSD.t605 VSSD.t784 123.087
R6968 VSSD.t1144 VSSD.t1178 123.087
R6969 VSSD.t610 VSSD.t745 123.087
R6970 VSSD.t923 VSSD.t117 122.044
R6971 VSSD.t321 VSSD.t1118 122.044
R6972 VSSD.t417 VSSD.t687 122.044
R6973 VSSD.t967 VSSD.t395 122.044
R6974 VSSD.t422 VSSD.t699 119.356
R6975 VSSD.t423 VSSD.t147 119.356
R6976 VSSD.t608 VSSD.t938 119.356
R6977 VSSD.t609 VSSD.t904 119.356
R6978 VSSD.t1142 VSSD.t704 119.356
R6979 VSSD.t394 VSSD.t131 119.356
R6980 VSSD.t922 VSSD.t842 119.356
R6981 VSSD.t919 VSSD.t715 119.356
R6982 VSSD.t994 VSSD.t746 119.356
R6983 VSSD.t993 VSSD.t637 119.356
R6984 VSSD.t982 VSSD.t422 118.112
R6985 VSSD.t652 VSSD.t608 118.112
R6986 VSSD.t104 VSSD.t1142 118.112
R6987 VSSD.t1152 VSSD.t922 118.112
R6988 VSSD.t975 VSSD.t994 118.112
R6989 VSSD.t555 VSSD.t691 116.906
R6990 VSSD.t627 VSSD.t278 116.906
R6991 VSSD.t296 VSSD.t1122 116.906
R6992 VSSD.t695 VSSD.t529 116.906
R6993 VSSD.t760 VSSD.t1080 116.008
R6994 VSSD.t751 VSSD.t481 116.008
R6995 VSSD.t409 VSSD.t206 116.008
R6996 VSSD.t262 VSSD.t264 116.008
R6997 VSSD.t491 VSSD.t1116 116.008
R6998 VSSD.t432 VSSD.t434 116.008
R6999 VSSD.t931 VSSD.t1114 116.008
R7000 VSSD.t594 VSSD.t598 116.008
R7001 VSSD.t438 VSSD.t1188 116.008
R7002 VSSD.t311 VSSD.t313 116.008
R7003 VSSD.t64 VSSD.t1157 116.008
R7004 VSSD.t506 VSSD 114.043
R7005 VSSD.t623 VSSD.t155 113.139
R7006 VSSD.t13 VSSD.t214 113.139
R7007 VSSD.t998 VSSD.t593 113.139
R7008 VSSD.t1126 VSSD.t940 113.139
R7009 VSSD.t274 VSSD.t628 113.139
R7010 VSSD.t1124 VSSD.t855 109.278
R7011 VSSD.t346 VSSD.t466 107.912
R7012 VSSD.t722 VSSD.t357 107.912
R7013 VSSD.t235 VSSD.t805 107.912
R7014 VSSD.t53 VSSD.t55 107.912
R7015 VSSD.t322 VSSD.t824 107.912
R7016 VSSD.t406 VSSD.t152 107.912
R7017 VSSD.t441 VSSD.t880 107.912
R7018 VSSD.t808 VSSD.t250 107.912
R7019 VSSD.t759 VSSD.t1028 104.436
R7020 VSSD.t73 VSSD.t420 104.436
R7021 VSSD.t143 VSSD.t145 104.436
R7022 VSSD.t208 VSSD.t765 104.436
R7023 VSSD.t906 VSSD.t902 104.436
R7024 VSSD.t71 VSSD.t453 104.436
R7025 VSSD.t663 VSSD.t661 104.436
R7026 VSSD.t1155 VSSD.t920 104.436
R7027 VSSD.t252 VSSD.t713 104.436
R7028 VSSD.t204 VSSD.t933 104.436
R7029 VSSD.t635 VSSD.t639 104.436
R7030 VSSD.n1666 VSSD.t624 100.001
R7031 VSSD.n1701 VSSD.t14 100.001
R7032 VSSD.n1737 VSSD.t999 100.001
R7033 VSSD.n1772 VSSD.t1127 100.001
R7034 VSSD.n1808 VSSD.t275 100.001
R7035 VSSD.n1470 VSSD.t167 100.001
R7036 VSSD.n1428 VSSD.t281 100.001
R7037 VSSD.n1540 VSSD.t1168 100.001
R7038 VSSD.n1576 VSSD.t518 100.001
R7039 VSSD.n1393 VSSD.t1001 100.001
R7040 VSSD.n1860 VSSD.t1084 100.001
R7041 VSSD.n91 VSSD.t1110 100.001
R7042 VSSD.n10 VSSD.t1087 100.001
R7043 VSSD.n19 VSSD.t1089 100.001
R7044 VSSD.n31 VSSD.t1092 100.001
R7045 VSSD.n40 VSSD.t1064 100.001
R7046 VSSD.n52 VSSD.t1068 100.001
R7047 VSSD.n61 VSSD.t1044 100.001
R7048 VSSD.n73 VSSD.t1105 100.001
R7049 VSSD.n82 VSSD.t1108 100.001
R7050 VSSD.n165 VSSD.t1170 100.001
R7051 VSSD.n181 VSSD.t731 100.001
R7052 VSSD.n197 VSSD.t698 100.001
R7053 VSSD.n216 VSSD.t725 100.001
R7054 VSSD.n232 VSSD.t1176 100.001
R7055 VSSD.n248 VSSD.t1172 100.001
R7056 VSSD.n156 VSSD.t692 100.001
R7057 VSSD.n144 VSSD.t279 100.001
R7058 VSSD.n132 VSSD.t1123 100.001
R7059 VSSD.n614 VSSD.t696 100.001
R7060 VSSD.n630 VSSD.t283 100.001
R7061 VSSD.n646 VSSD.t945 100.001
R7062 VSSD.n818 VSSD.t1027 100.001
R7063 VSSD.n819 VSSD.t1098 100.001
R7064 VSSD.n833 VSSD.t1100 100.001
R7065 VSSD.n834 VSSD.t1079 100.001
R7066 VSSD.n848 VSSD.t1066 100.001
R7067 VSSD.n849 VSSD.t1025 100.001
R7068 VSSD.n863 VSSD.t1073 100.001
R7069 VSSD.n864 VSSD.t1036 100.001
R7070 VSSD.n878 VSSD.t1055 100.001
R7071 VSSD.n879 VSSD.t1007 100.001
R7072 VSSD.n893 VSSD.t1090 100.001
R7073 VSSD.n894 VSSD.t1062 100.001
R7074 VSSD.n908 VSSD.t1085 100.001
R7075 VSSD.n909 VSSD.t1059 100.001
R7076 VSSD.n923 VSSD.t1040 100.001
R7077 VSSD.n924 VSSD.t1103 100.001
R7078 VSSD.n938 VSSD.t1013 100.001
R7079 VSSD.n939 VSSD.t1034 100.001
R7080 VSSD.n953 VSSD.t1065 100.001
R7081 VSSD.n954 VSSD.t1019 100.001
R7082 VSSD.t188 VSSD.t108 99.4355
R7083 VSSD.t1173 VSSD.t330 99.4355
R7084 VSSD.t9 VSSD.t93 99.4355
R7085 VSSD.t693 VSSD.t197 99.4355
R7086 VSSD.t164 VSSD.t888 99.4355
R7087 VSSD.t985 VSSD.t612 94.4449
R7088 VSSD VSSD.t760 92.5303
R7089 VSSD.t15 VSSD.t981 92.4969
R7090 VSSD.t513 VSSD.t156 92.4969
R7091 VSSD.t826 VSSD.t741 92.4969
R7092 VSSD.t367 VSSD.t942 92.4969
R7093 VSSD.t206 VSSD 89.7682
R7094 VSSD.t1116 VSSD 89.7682
R7095 VSSD.t1114 VSSD 89.7682
R7096 VSSD.t1188 VSSD 89.7682
R7097 VSSD.t1157 VSSD 89.7682
R7098 VSSD.t43 VSSD.t270 89.5173
R7099 VSSD.t767 VSSD.t266 89.5173
R7100 VSSD.t703 VSSD.t511 89.5173
R7101 VSSD.t52 VSSD.t726 89.5173
R7102 VSSD.t783 VSSD.t728 89.5173
R7103 VSSD.t377 VSSD.t372 86.5984
R7104 VSSD.t546 VSSD.t377 86.5984
R7105 VSSD.t857 VSSD.t548 86.5984
R7106 VSSD.t665 VSSD.t668 84.2917
R7107 VSSD.t949 VSSD.t386 84.2917
R7108 VSSD.t849 VSSD.t740 84.2917
R7109 VSSD.t62 VSSD.t818 84.2917
R7110 VSSD.t551 VSSD.t778 84.2917
R7111 VSSD.t757 VSSD.t965 84.2917
R7112 VSSD.t333 VSSD.t660 84.2917
R7113 VSSD.t556 VSSD.t970 84.2917
R7114 VSSD.t215 VSSD.t867 84.2917
R7115 VSSD.t865 VSSD.t912 84.2917
R7116 VSSD.t466 VSSD 83.5041
R7117 VSSD.t805 VSSD 83.5041
R7118 VSSD.t824 VSSD 83.5041
R7119 VSSD.t880 VSSD 83.5041
R7120 VSSD VSSD.t759 83.3009
R7121 VSSD.t853 VSSD.t1164 80.4129
R7122 VSSD.t550 VSSD.t1124 74.2273
R7123 VSSD.n1636 VSSD.t1029 72.8576
R7124 VSSD.n1377 VSSD.t271 72.8576
R7125 VSSD.n1692 VSSD.t267 72.8576
R7126 VSSD.n1354 VSSD.t512 72.8576
R7127 VSSD.n1763 VSSD.t727 72.8576
R7128 VSSD.n1331 VSSD.t729 72.8576
R7129 VSSD.n1461 VSSD.t165 72.8576
R7130 VSSD.n1497 VSSD.t694 72.8576
R7131 VSSD.n1417 VSSD.t10 72.8576
R7132 VSSD.n1567 VSSD.t1174 72.8576
R7133 VSSD.n1603 VSSD.t189 72.8576
R7134 VSSD.n1387 VSSD.t1081 72.8576
R7135 VSSD.n1868 VSSD.t1011 72.8576
R7136 VSSD.n96 VSSD.t1057 72.8576
R7137 VSSD.n14 VSSD.t1052 72.8576
R7138 VSSD.n16 VSSD.t1094 72.8576
R7139 VSSD.n35 VSSD.t1017 72.8576
R7140 VSSD.n37 VSSD.t1070 72.8576
R7141 VSSD.n56 VSSD.t1033 72.8576
R7142 VSSD.n58 VSSD.t1077 72.8576
R7143 VSSD.n77 VSSD.t1102 72.8576
R7144 VSSD.n79 VSSD.t1050 72.8576
R7145 VSSD.n168 VSSD.t516 72.8576
R7146 VSSD.n184 VSSD.t690 72.8576
R7147 VSSD.n200 VSSD.t277 72.8576
R7148 VSSD.n219 VSSD.t1121 72.8576
R7149 VSSD.n235 VSSD.t269 72.8576
R7150 VSSD.n251 VSSD.t622 72.8576
R7151 VSSD.n514 VSSD.t16 72.8576
R7152 VSSD.n551 VSSD.t514 72.8576
R7153 VSSD.n592 VSSD.t827 72.8576
R7154 VSSD.n617 VSSD.t943 72.8576
R7155 VSSD.n633 VSSD.t187 72.8576
R7156 VSSD.n649 VSSD.t1125 72.8576
R7157 VSSD.n1285 VSSD.t1097 72.8576
R7158 VSSD.n1286 VSSD.t1072 72.8576
R7159 VSSD.n1250 VSSD.t1075 72.8576
R7160 VSSD.n1251 VSSD.t1042 72.8576
R7161 VSSD.n1215 VSSD.t1048 72.8576
R7162 VSSD.n1216 VSSD.t1106 72.8576
R7163 VSSD.n1180 VSSD.t1054 72.8576
R7164 VSSD.n1181 VSSD.t1111 72.8576
R7165 VSSD.n1145 VSSD.t1021 72.8576
R7166 VSSD.n1146 VSSD.t1095 72.8576
R7167 VSSD.n1110 VSSD.t1031 72.8576
R7168 VSSD.n1111 VSSD.t1099 72.8576
R7169 VSSD.n1075 VSSD.t1023 72.8576
R7170 VSSD.n1076 VSSD.t1096 72.8576
R7171 VSSD.n1040 VSSD.t1060 72.8576
R7172 VSSD.n1041 VSSD.t1009 72.8576
R7173 VSSD.n1005 VSSD.t1082 72.8576
R7174 VSSD.n1006 VSSD.t1046 72.8576
R7175 VSSD.n970 VSSD.t1074 72.8576
R7176 VSSD.n971 VSSD.t1038 72.8576
R7177 VSSD.n766 VSSD.t413 71.4899
R7178 VSSD.n766 VSSD.t162 71.4899
R7179 VSSD.n1666 VSSD.t148 70.0005
R7180 VSSD.n1701 VSSD.t905 70.0005
R7181 VSSD.n1737 VSSD.t132 70.0005
R7182 VSSD.n1772 VSSD.t716 70.0005
R7183 VSSD.n1808 VSSD.t638 70.0005
R7184 VSSD.n1470 VSSD.t869 70.0005
R7185 VSSD.n1428 VSSD.t597 70.0005
R7186 VSSD.n1540 VSSD.t431 70.0005
R7187 VSSD.n1576 VSSD.t533 70.0005
R7188 VSSD.n1393 VSSD.t480 70.0005
R7189 VSSD.n1860 VSSD.t913 70.0005
R7190 VSSD.n91 VSSD.t216 70.0005
R7191 VSSD.n10 VSSD.t666 70.0005
R7192 VSSD.n19 VSSD.t387 70.0005
R7193 VSSD.n31 VSSD.t850 70.0005
R7194 VSSD.n40 VSSD.t819 70.0005
R7195 VSSD.n52 VSSD.t552 70.0005
R7196 VSSD.n61 VSSD.t966 70.0005
R7197 VSSD.n73 VSSD.t334 70.0005
R7198 VSSD.n82 VSSD.t971 70.0005
R7199 VSSD.n165 VSSD.t222 70.0005
R7200 VSSD.n181 VSSD.t1134 70.0005
R7201 VSSD.n197 VSSD.t748 70.0005
R7202 VSSD.n216 VSSD.t952 70.0005
R7203 VSSD.n232 VSSD.t342 70.0005
R7204 VSSD.n248 VSSD.t1131 70.0005
R7205 VSSD.n156 VSSD.t356 70.0005
R7206 VSSD.n144 VSSD.t581 70.0005
R7207 VSSD.n132 VSSD.t115 70.0005
R7208 VSSD.n614 VSSD.t811 70.0005
R7209 VSSD.n630 VSSD.t47 70.0005
R7210 VSSD.n646 VSSD.t1165 70.0005
R7211 VSSD.n818 VSSD.t136 70.0005
R7212 VSSD.n819 VSSD.t8 70.0005
R7213 VSSD.n833 VSSD.t600 70.0005
R7214 VSSD.n834 VSSD.t287 70.0005
R7215 VSSD.n848 VSSD.t1129 70.0005
R7216 VSSD.n849 VSSD.t78 70.0005
R7217 VSSD.n863 VSSD.t925 70.0005
R7218 VSSD.n864 VSSD.t128 70.0005
R7219 VSSD.n878 VSSD.t735 70.0005
R7220 VSSD.n879 VSSD.t138 70.0005
R7221 VSSD.n893 VSSD.t802 70.0005
R7222 VSSD.n894 VSSD.t961 70.0005
R7223 VSSD.n908 VSSD.t1149 70.0005
R7224 VSSD.n909 VSSD.t579 70.0005
R7225 VSSD.n923 VSSD.t567 70.0005
R7226 VSSD.n924 VSSD.t753 70.0005
R7227 VSSD.n938 VSSD.t732 70.0005
R7228 VSSD.n939 VSSD.t304 70.0005
R7229 VSSD.n953 VSSD.t499 70.0005
R7230 VSSD.n954 VSSD.t800 70.0005
R7231 VSSD.t851 VSSD.t381 68.0417
R7232 VSSD.t1190 VSSD.t930 68.0417
R7233 VSSD VSSD.n208 67.8232
R7234 VSSD.t292 VSSD.t650 67.4335
R7235 VSSD.t290 VSSD.t391 67.4335
R7236 VSSD.t509 VSSD.t382 67.4335
R7237 VSSD.t876 VSSD.t384 67.4335
R7238 VSSD.t845 VSSD.t646 67.4335
R7239 VSSD.t847 VSSD.t561 67.4335
R7240 VSSD.t682 VSSD.t814 67.4335
R7241 VSSD.t472 VSSD.t816 67.4335
R7242 VSSD.t553 VSSD.t822 67.4335
R7243 VSSD.t180 VSSD.t232 67.4335
R7244 VSSD.t110 VSSD.t989 67.4335
R7245 VSSD.t648 VSSD.t991 67.4335
R7246 VSSD.t1136 VSSD.t305 67.4335
R7247 VSSD.t1138 VSSD.t795 67.4335
R7248 VSSD.t36 VSSD.t788 67.4335
R7249 VSSD.t644 VSSD.t973 67.4335
R7250 VSSD.t219 VSSD.t470 67.4335
R7251 VSSD.t217 VSSD.t495 67.4335
R7252 VSSD.t326 VSSD.t914 67.4335
R7253 VSSD.t878 VSSD.t910 67.4335
R7254 VSSD.t184 VSSD.t375 63.918
R7255 VSSD.t548 VSSD.t944 60.8252
R7256 VSSD.n1377 VSSD.t241 60.5809
R7257 VSSD.n1692 VSSD.t486 60.5809
R7258 VSSD.n1354 VSSD.t606 60.5809
R7259 VSSD.n1763 VSSD.t1145 60.5809
R7260 VSSD.n1331 VSSD.t611 60.5809
R7261 VSSD.n1461 VSSD.t710 60.5809
R7262 VSSD.n1497 VSSD.t177 60.5809
R7263 VSSD.n1417 VSSD.t302 60.5809
R7264 VSSD.n1567 VSSD.t488 60.5809
R7265 VSSD.n1603 VSSD.t477 60.5809
R7266 VSSD.n1868 VSSD.t403 60.5809
R7267 VSSD.n96 VSSD.t1003 60.5809
R7268 VSSD.n14 VSSD.t92 60.5809
R7269 VSSD.n16 VSSD.t401 60.5809
R7270 VSSD.n35 VSSD.t541 60.5809
R7271 VSSD.n37 VSSD.t40 60.5809
R7272 VSSD.n56 VSSD.t702 60.5809
R7273 VSSD.n58 VSSD.t196 60.5809
R7274 VSSD.n77 VSSD.t412 60.5809
R7275 VSSD.n79 VSSD.t718 60.5809
R7276 VSSD.n168 VSSD.t369 60.5809
R7277 VSSD.n184 VSSD.t360 60.5809
R7278 VSSD.n200 VSSD.t706 60.5809
R7279 VSSD.n219 VSSD.t316 60.5809
R7280 VSSD.n235 VSSD.t299 60.5809
R7281 VSSD.n251 VSSD.t844 60.5809
R7282 VSSD.n514 VSSD.t862 60.5809
R7283 VSSD.n551 VSSD.t19 60.5809
R7284 VSSD.n592 VSSD.t681 60.5809
R7285 VSSD.n617 VSSD.t929 60.5809
R7286 VSSD.n633 VSSD.t909 60.5809
R7287 VSSD.n649 VSSD.t459 60.5809
R7288 VSSD.n1285 VSSD.t336 60.5809
R7289 VSSD.n1286 VSSD.t86 60.5809
R7290 VSSD.n1250 VSSD.t405 60.5809
R7291 VSSD.n1251 VSSD.t984 60.5809
R7292 VSSD.n1215 VSSD.t836 60.5809
R7293 VSSD.n1216 VSSD.t835 60.5809
R7294 VSSD.n1180 VSSD.t63 60.5809
R7295 VSSD.n1181 VSSD.t35 60.5809
R7296 VSSD.n1145 VSSD.t389 60.5809
R7297 VSSD.n1146 VSSD.t489 60.5809
R7298 VSSD.n1110 VSSD.t828 60.5809
R7299 VSSD.n1111 VSSD.t494 60.5809
R7300 VSSD.n1075 VSSD.t607 60.5809
R7301 VSSD.n1076 VSSD.t179 60.5809
R7302 VSSD.n1040 VSSD.t957 60.5809
R7303 VSSD.n1041 VSSD.t679 60.5809
R7304 VSSD.n1005 VSSD.t841 60.5809
R7305 VSSD.n1006 VSSD.t941 60.5809
R7306 VSSD.n970 VSSD.t962 60.5809
R7307 VSSD.n971 VSSD.t345 60.5809
R7308 VSSD.t458 VSSD.t859 59.7943
R7309 VSSD.t916 VSSD.n2014 50.3709
R7310 VSSD.t379 VSSD.t1190 44.3304
R7311 VSSD.n1634 VSSD.n1632 43.9358
R7312 VSSD.n1628 VSSD.n1627 43.9358
R7313 VSSD.n767 VSSD.n766 43.3338
R7314 VSSD.t859 VSSD.t379 42.2685
R7315 VSSD.n1643 VSSD.t74 38.5719
R7316 VSSD.n1643 VSSD.t421 38.5719
R7317 VSSD.n1371 VSSD.t209 38.5719
R7318 VSSD.n1371 VSSD.t766 38.5719
R7319 VSSD.n1714 VSSD.t72 38.5719
R7320 VSSD.n1714 VSSD.t454 38.5719
R7321 VSSD.n1348 VSSD.t1156 38.5719
R7322 VSSD.n1348 VSSD.t921 38.5719
R7323 VSSD.n1785 VSSD.t205 38.5719
R7324 VSSD.n1785 VSSD.t934 38.5719
R7325 VSSD.n1447 VSSD.t65 38.5719
R7326 VSSD.n1447 VSSD.t1158 38.5719
R7327 VSSD.n1483 VSSD.t439 38.5719
R7328 VSSD.n1483 VSSD.t1189 38.5719
R7329 VSSD.n1517 VSSD.t932 38.5719
R7330 VSSD.n1517 VSSD.t1115 38.5719
R7331 VSSD.n1553 VSSD.t492 38.5719
R7332 VSSD.n1553 VSSD.t1117 38.5719
R7333 VSSD.n1589 VSSD.t410 38.5719
R7334 VSSD.n1589 VSSD.t207 38.5719
R7335 VSSD.n1852 VSSD.t327 38.5719
R7336 VSSD.n1852 VSSD.t879 38.5719
R7337 VSSD.n5 VSSD.t651 38.5719
R7338 VSSD.n5 VSSD.t392 38.5719
R7339 VSSD.n22 VSSD.t510 38.5719
R7340 VSSD.n22 VSSD.t877 38.5719
R7341 VSSD.n26 VSSD.t647 38.5719
R7342 VSSD.n26 VSSD.t562 38.5719
R7343 VSSD.n43 VSSD.t683 38.5719
R7344 VSSD.n43 VSSD.t473 38.5719
R7345 VSSD.n47 VSSD.t823 38.5719
R7346 VSSD.n47 VSSD.t233 38.5719
R7347 VSSD.n64 VSSD.t111 38.5719
R7348 VSSD.n64 VSSD.t649 38.5719
R7349 VSSD.n68 VSSD.t306 38.5719
R7350 VSSD.n68 VSSD.t796 38.5719
R7351 VSSD.n85 VSSD.t37 38.5719
R7352 VSSD.n85 VSSD.t645 38.5719
R7353 VSSD.n89 VSSD.t471 38.5719
R7354 VSSD.n89 VSSD.t496 38.5719
R7355 VSSD.n173 VSSD.t947 38.5719
R7356 VSSD.n173 VSSD.t308 38.5719
R7357 VSSD.n189 VSSD.t67 38.5719
R7358 VSSD.n189 VSSD.t883 38.5719
R7359 VSSD.n205 VSSD.t677 38.5719
R7360 VSSD.n205 VSSD.t804 38.5719
R7361 VSSD.n224 VSSD.t428 38.5719
R7362 VSSD.n224 VSSD.t559 38.5719
R7363 VSSD.n240 VSSD.t774 38.5719
R7364 VSSD.n240 VSSD.t310 38.5719
R7365 VSSD.n256 VSSD.t831 38.5719
R7366 VSSD.n256 VSSD.t469 38.5719
R7367 VSSD.n149 VSSD.t236 38.5719
R7368 VSSD.n149 VSSD.t806 38.5719
R7369 VSSD.n568 VSSD.t323 38.5719
R7370 VSSD.n568 VSSD.t825 38.5719
R7371 VSSD.n125 VSSD.t442 38.5719
R7372 VSSD.n125 VSSD.t881 38.5719
R7373 VSSD.n622 VSSD.t397 38.5719
R7374 VSSD.n622 VSSD.t475 38.5719
R7375 VSSD.n638 VSSD.t347 38.5719
R7376 VSSD.n638 VSSD.t467 38.5719
R7377 VSSD.n654 VSSD.t986 38.5719
R7378 VSSD.n654 VSSD.t821 38.5719
R7379 VSSD.n809 VSSD.t632 38.5719
R7380 VSSD.n809 VSSD.t371 38.5719
R7381 VSSD.n810 VSSD.t742 38.5719
R7382 VSSD.n810 VSSD.t1177 38.5719
R7383 VSSD.n823 VSSD.t572 38.5719
R7384 VSSD.n823 VSSD.t895 38.5719
R7385 VSSD.n824 VSSD.t522 38.5719
R7386 VSSD.n824 VSSD.t82 38.5719
R7387 VSSD.n838 VSSD.t658 38.5719
R7388 VSSD.n838 VSSD.t963 38.5719
R7389 VSSD.n839 VSSD.t425 38.5719
R7390 VSSD.n839 VSSD.t674 38.5719
R7391 VSSD.n853 VSSD.t978 38.5719
R7392 VSSD.n853 VSSD.t655 38.5719
R7393 VSSD.n854 VSSD.t60 38.5719
R7394 VSSD.n854 VSSD.t987 38.5719
R7395 VSSD.n868 VSSD.t1159 38.5719
R7396 VSSD.n868 VSSD.t3 38.5719
R7397 VSSD.n869 VSSD.t871 38.5719
R7398 VSSD.n869 VSSD.t5 38.5719
R7399 VSSD.n883 VSSD.t29 38.5719
R7400 VSSD.n883 VSSD.t449 38.5719
R7401 VSSD.n884 VSSD.t113 38.5719
R7402 VSSD.n884 VSSD.t448 38.5719
R7403 VSSD.n898 VSSD.t838 38.5719
R7404 VSSD.n898 VSSD.t124 38.5719
R7405 VSSD.n899 VSSD.t791 38.5719
R7406 VSSD.n899 VSSD.t125 38.5719
R7407 VSSD.n913 VSSD.t739 38.5719
R7408 VSSD.n913 VSSD.t230 38.5719
R7409 VSSD.n914 VSSD.t437 38.5719
R7410 VSSD.n914 VSSD.t231 38.5719
R7411 VSSD.n928 VSSD.t997 38.5719
R7412 VSSD.n928 VSSD.t524 38.5719
R7413 VSSD.n929 VSSD.t203 38.5719
R7414 VSSD.n929 VSSD.t527 38.5719
R7415 VSSD.n943 VSSD.t25 38.5719
R7416 VSSD.n943 VSSD.t257 38.5719
R7417 VSSD.n944 VSSD.t762 38.5719
R7418 VSSD.n944 VSSD.t1146 38.5719
R7419 VSSD VSSD.t73 38.5425
R7420 VSSD VSSD.t208 38.5425
R7421 VSSD VSSD.t71 38.5425
R7422 VSSD VSSD.t1155 38.5425
R7423 VSSD VSSD.t204 38.5425
R7424 VSSD.n763 VSSD 37.256
R7425 VSSD.n765 VSSD.t346 35.9713
R7426 VSSD.t398 VSSD.t916 35.5561
R7427 VSSD.t612 VSSD.t398 35.1857
R7428 VSSD.n764 VSSD.t967 34.6866
R7429 VSSD.n1635 VSSD.n1634 34.6358
R7430 VSSD.n1638 VSSD.n1383 34.6358
R7431 VSSD.n1650 VSSD.n1649 34.6358
R7432 VSSD.n1650 VSSD.n1380 34.6358
R7433 VSSD.n1654 VSSD.n1380 34.6358
R7434 VSSD.n1655 VSSD.n1654 34.6358
R7435 VSSD.n1656 VSSD.n1655 34.6358
R7436 VSSD.n1660 VSSD.n1659 34.6358
R7437 VSSD.n1661 VSSD.n1660 34.6358
R7438 VSSD.n1661 VSSD.n1375 34.6358
R7439 VSSD.n1665 VSSD.n1375 34.6358
R7440 VSSD.n1669 VSSD.n1668 34.6358
R7441 VSSD.n1669 VSSD.n1373 34.6358
R7442 VSSD.n1685 VSSD.n1368 34.6358
R7443 VSSD.n1686 VSSD.n1685 34.6358
R7444 VSSD.n1687 VSSD.n1686 34.6358
R7445 VSSD.n1687 VSSD.n1366 34.6358
R7446 VSSD.n1691 VSSD.n1366 34.6358
R7447 VSSD.n1695 VSSD.n1694 34.6358
R7448 VSSD.n1695 VSSD.n1364 34.6358
R7449 VSSD.n1699 VSSD.n1364 34.6358
R7450 VSSD.n1700 VSSD.n1699 34.6358
R7451 VSSD.n1703 VSSD.n1362 34.6358
R7452 VSSD.n1707 VSSD.n1362 34.6358
R7453 VSSD.n1721 VSSD.n1720 34.6358
R7454 VSSD.n1721 VSSD.n1357 34.6358
R7455 VSSD.n1725 VSSD.n1357 34.6358
R7456 VSSD.n1726 VSSD.n1725 34.6358
R7457 VSSD.n1727 VSSD.n1726 34.6358
R7458 VSSD.n1731 VSSD.n1730 34.6358
R7459 VSSD.n1732 VSSD.n1731 34.6358
R7460 VSSD.n1732 VSSD.n1352 34.6358
R7461 VSSD.n1736 VSSD.n1352 34.6358
R7462 VSSD.n1740 VSSD.n1739 34.6358
R7463 VSSD.n1740 VSSD.n1350 34.6358
R7464 VSSD.n1756 VSSD.n1345 34.6358
R7465 VSSD.n1757 VSSD.n1756 34.6358
R7466 VSSD.n1758 VSSD.n1757 34.6358
R7467 VSSD.n1758 VSSD.n1343 34.6358
R7468 VSSD.n1762 VSSD.n1343 34.6358
R7469 VSSD.n1766 VSSD.n1765 34.6358
R7470 VSSD.n1766 VSSD.n1341 34.6358
R7471 VSSD.n1770 VSSD.n1341 34.6358
R7472 VSSD.n1771 VSSD.n1770 34.6358
R7473 VSSD.n1774 VSSD.n1339 34.6358
R7474 VSSD.n1778 VSSD.n1339 34.6358
R7475 VSSD.n1792 VSSD.n1791 34.6358
R7476 VSSD.n1792 VSSD.n1334 34.6358
R7477 VSSD.n1796 VSSD.n1334 34.6358
R7478 VSSD.n1797 VSSD.n1796 34.6358
R7479 VSSD.n1798 VSSD.n1797 34.6358
R7480 VSSD.n1802 VSSD.n1801 34.6358
R7481 VSSD.n1803 VSSD.n1802 34.6358
R7482 VSSD.n1803 VSSD.n1329 34.6358
R7483 VSSD.n1807 VSSD.n1329 34.6358
R7484 VSSD.n1811 VSSD.n1810 34.6358
R7485 VSSD.n1811 VSSD.n1327 34.6358
R7486 VSSD.n1460 VSSD.n1442 34.6358
R7487 VSSD.n1456 VSSD.n1442 34.6358
R7488 VSSD.n1456 VSSD.n1455 34.6358
R7489 VSSD.n1455 VSSD.n1454 34.6358
R7490 VSSD.n1454 VSSD.n1444 34.6358
R7491 VSSD.n1469 VSSD.n1468 34.6358
R7492 VSSD.n1468 VSSD.n1440 34.6358
R7493 VSSD.n1464 VSSD.n1440 34.6358
R7494 VSSD.n1464 VSSD.n1463 34.6358
R7495 VSSD.n1476 VSSD.n1438 34.6358
R7496 VSSD.n1472 VSSD.n1438 34.6358
R7497 VSSD.n1496 VSSD.n1495 34.6358
R7498 VSSD.n1495 VSSD.n1432 34.6358
R7499 VSSD.n1491 VSSD.n1432 34.6358
R7500 VSSD.n1491 VSSD.n1490 34.6358
R7501 VSSD.n1490 VSSD.n1489 34.6358
R7502 VSSD.n1505 VSSD.n1504 34.6358
R7503 VSSD.n1504 VSSD.n1503 34.6358
R7504 VSSD.n1503 VSSD.n1430 34.6358
R7505 VSSD.n1499 VSSD.n1430 34.6358
R7506 VSSD.n1510 VSSD.n1509 34.6358
R7507 VSSD.n1509 VSSD.n1426 34.6358
R7508 VSSD.n1530 VSSD.n1529 34.6358
R7509 VSSD.n1529 VSSD.n1528 34.6358
R7510 VSSD.n1528 VSSD.n1420 34.6358
R7511 VSSD.n1524 VSSD.n1420 34.6358
R7512 VSSD.n1524 VSSD.n1523 34.6358
R7513 VSSD.n1539 VSSD.n1415 34.6358
R7514 VSSD.n1535 VSSD.n1415 34.6358
R7515 VSSD.n1535 VSSD.n1534 34.6358
R7516 VSSD.n1534 VSSD.n1533 34.6358
R7517 VSSD.n1543 VSSD.n1413 34.6358
R7518 VSSD.n1543 VSSD.n1542 34.6358
R7519 VSSD.n1566 VSSD.n1407 34.6358
R7520 VSSD.n1562 VSSD.n1407 34.6358
R7521 VSSD.n1562 VSSD.n1561 34.6358
R7522 VSSD.n1561 VSSD.n1560 34.6358
R7523 VSSD.n1560 VSSD.n1409 34.6358
R7524 VSSD.n1575 VSSD.n1574 34.6358
R7525 VSSD.n1574 VSSD.n1405 34.6358
R7526 VSSD.n1570 VSSD.n1405 34.6358
R7527 VSSD.n1570 VSSD.n1569 34.6358
R7528 VSSD.n1582 VSSD.n1403 34.6358
R7529 VSSD.n1578 VSSD.n1403 34.6358
R7530 VSSD.n1602 VSSD.n1601 34.6358
R7531 VSSD.n1601 VSSD.n1397 34.6358
R7532 VSSD.n1597 VSSD.n1397 34.6358
R7533 VSSD.n1597 VSSD.n1596 34.6358
R7534 VSSD.n1596 VSSD.n1595 34.6358
R7535 VSSD.n1611 VSSD.n1610 34.6358
R7536 VSSD.n1610 VSSD.n1609 34.6358
R7537 VSSD.n1609 VSSD.n1395 34.6358
R7538 VSSD.n1605 VSSD.n1395 34.6358
R7539 VSSD.n1616 VSSD.n1615 34.6358
R7540 VSSD.n1615 VSSD.n1391 34.6358
R7541 VSSD.n1623 VSSD.n1622 34.6358
R7542 VSSD.n1627 VSSD.n1385 34.6358
R7543 VSSD.n1839 VSSD.n1838 34.6358
R7544 VSSD.n1859 VSSD.n1858 34.6358
R7545 VSSD.n1867 VSSD.n1866 34.6358
R7546 VSSD.n1866 VSSD.n98 34.6358
R7547 VSSD.n1862 VSSD.n98 34.6358
R7548 VSSD.n1876 VSSD.n1875 34.6358
R7549 VSSD.n1875 VSSD.n1874 34.6358
R7550 VSSD.n1874 VSSD.n94 34.6358
R7551 VSSD.n1880 VSSD.n1879 34.6358
R7552 VSSD.n2006 VSSD.n8 34.6358
R7553 VSSD.n2002 VSSD.n2001 34.6358
R7554 VSSD.n2001 VSSD.n2000 34.6358
R7555 VSSD.n2000 VSSD.n12 34.6358
R7556 VSSD.n1994 VSSD.n1993 34.6358
R7557 VSSD.n1993 VSSD.n17 34.6358
R7558 VSSD.n1989 VSSD.n17 34.6358
R7559 VSSD.n1987 VSSD.n1986 34.6358
R7560 VSSD.n1975 VSSD.n29 34.6358
R7561 VSSD.n1971 VSSD.n1970 34.6358
R7562 VSSD.n1970 VSSD.n1969 34.6358
R7563 VSSD.n1969 VSSD.n33 34.6358
R7564 VSSD.n1963 VSSD.n1962 34.6358
R7565 VSSD.n1962 VSSD.n38 34.6358
R7566 VSSD.n1958 VSSD.n38 34.6358
R7567 VSSD.n1956 VSSD.n1955 34.6358
R7568 VSSD.n1944 VSSD.n50 34.6358
R7569 VSSD.n1940 VSSD.n1939 34.6358
R7570 VSSD.n1939 VSSD.n1938 34.6358
R7571 VSSD.n1938 VSSD.n54 34.6358
R7572 VSSD.n1932 VSSD.n1931 34.6358
R7573 VSSD.n1931 VSSD.n59 34.6358
R7574 VSSD.n1927 VSSD.n59 34.6358
R7575 VSSD.n1925 VSSD.n1924 34.6358
R7576 VSSD.n1913 VSSD.n71 34.6358
R7577 VSSD.n1909 VSSD.n1908 34.6358
R7578 VSSD.n1908 VSSD.n1907 34.6358
R7579 VSSD.n1907 VSSD.n75 34.6358
R7580 VSSD.n1901 VSSD.n1900 34.6358
R7581 VSSD.n1900 VSSD.n80 34.6358
R7582 VSSD.n1896 VSSD.n80 34.6358
R7583 VSSD.n1894 VSSD.n1893 34.6358
R7584 VSSD.n1314 VSSD.n1313 34.6358
R7585 VSSD.n1305 VSSD.n807 34.6358
R7586 VSSD.n1292 VSSD.n814 34.6358
R7587 VSSD.n1293 VSSD.n1292 34.6358
R7588 VSSD.n1294 VSSD.n1293 34.6358
R7589 VSSD.n1294 VSSD.n812 34.6358
R7590 VSSD.n1298 VSSD.n812 34.6358
R7591 VSSD.n1279 VSSD.n816 34.6358
R7592 VSSD.n1283 VSSD.n816 34.6358
R7593 VSSD.n1284 VSSD.n1283 34.6358
R7594 VSSD.n1288 VSSD.n1284 34.6358
R7595 VSSD.n1276 VSSD.n820 34.6358
R7596 VSSD.n1277 VSSD.n1276 34.6358
R7597 VSSD.n1257 VSSD.n829 34.6358
R7598 VSSD.n1258 VSSD.n1257 34.6358
R7599 VSSD.n1259 VSSD.n1258 34.6358
R7600 VSSD.n1259 VSSD.n827 34.6358
R7601 VSSD.n1263 VSSD.n827 34.6358
R7602 VSSD.n1244 VSSD.n831 34.6358
R7603 VSSD.n1248 VSSD.n831 34.6358
R7604 VSSD.n1249 VSSD.n1248 34.6358
R7605 VSSD.n1253 VSSD.n1249 34.6358
R7606 VSSD.n1241 VSSD.n835 34.6358
R7607 VSSD.n1242 VSSD.n1241 34.6358
R7608 VSSD.n1222 VSSD.n844 34.6358
R7609 VSSD.n1223 VSSD.n1222 34.6358
R7610 VSSD.n1224 VSSD.n1223 34.6358
R7611 VSSD.n1224 VSSD.n842 34.6358
R7612 VSSD.n1228 VSSD.n842 34.6358
R7613 VSSD.n1209 VSSD.n846 34.6358
R7614 VSSD.n1213 VSSD.n846 34.6358
R7615 VSSD.n1214 VSSD.n1213 34.6358
R7616 VSSD.n1218 VSSD.n1214 34.6358
R7617 VSSD.n1206 VSSD.n850 34.6358
R7618 VSSD.n1207 VSSD.n1206 34.6358
R7619 VSSD.n1187 VSSD.n859 34.6358
R7620 VSSD.n1188 VSSD.n1187 34.6358
R7621 VSSD.n1189 VSSD.n1188 34.6358
R7622 VSSD.n1189 VSSD.n857 34.6358
R7623 VSSD.n1193 VSSD.n857 34.6358
R7624 VSSD.n1174 VSSD.n861 34.6358
R7625 VSSD.n1178 VSSD.n861 34.6358
R7626 VSSD.n1179 VSSD.n1178 34.6358
R7627 VSSD.n1183 VSSD.n1179 34.6358
R7628 VSSD.n1171 VSSD.n865 34.6358
R7629 VSSD.n1172 VSSD.n1171 34.6358
R7630 VSSD.n1152 VSSD.n874 34.6358
R7631 VSSD.n1153 VSSD.n1152 34.6358
R7632 VSSD.n1154 VSSD.n1153 34.6358
R7633 VSSD.n1154 VSSD.n872 34.6358
R7634 VSSD.n1158 VSSD.n872 34.6358
R7635 VSSD.n1139 VSSD.n876 34.6358
R7636 VSSD.n1143 VSSD.n876 34.6358
R7637 VSSD.n1144 VSSD.n1143 34.6358
R7638 VSSD.n1148 VSSD.n1144 34.6358
R7639 VSSD.n1136 VSSD.n880 34.6358
R7640 VSSD.n1137 VSSD.n1136 34.6358
R7641 VSSD.n1117 VSSD.n889 34.6358
R7642 VSSD.n1118 VSSD.n1117 34.6358
R7643 VSSD.n1119 VSSD.n1118 34.6358
R7644 VSSD.n1119 VSSD.n887 34.6358
R7645 VSSD.n1123 VSSD.n887 34.6358
R7646 VSSD.n1104 VSSD.n891 34.6358
R7647 VSSD.n1108 VSSD.n891 34.6358
R7648 VSSD.n1109 VSSD.n1108 34.6358
R7649 VSSD.n1113 VSSD.n1109 34.6358
R7650 VSSD.n1101 VSSD.n895 34.6358
R7651 VSSD.n1102 VSSD.n1101 34.6358
R7652 VSSD.n1082 VSSD.n904 34.6358
R7653 VSSD.n1083 VSSD.n1082 34.6358
R7654 VSSD.n1084 VSSD.n1083 34.6358
R7655 VSSD.n1084 VSSD.n902 34.6358
R7656 VSSD.n1088 VSSD.n902 34.6358
R7657 VSSD.n1069 VSSD.n906 34.6358
R7658 VSSD.n1073 VSSD.n906 34.6358
R7659 VSSD.n1074 VSSD.n1073 34.6358
R7660 VSSD.n1078 VSSD.n1074 34.6358
R7661 VSSD.n1066 VSSD.n910 34.6358
R7662 VSSD.n1067 VSSD.n1066 34.6358
R7663 VSSD.n1047 VSSD.n919 34.6358
R7664 VSSD.n1048 VSSD.n1047 34.6358
R7665 VSSD.n1049 VSSD.n1048 34.6358
R7666 VSSD.n1049 VSSD.n917 34.6358
R7667 VSSD.n1053 VSSD.n917 34.6358
R7668 VSSD.n1034 VSSD.n921 34.6358
R7669 VSSD.n1038 VSSD.n921 34.6358
R7670 VSSD.n1039 VSSD.n1038 34.6358
R7671 VSSD.n1043 VSSD.n1039 34.6358
R7672 VSSD.n1031 VSSD.n925 34.6358
R7673 VSSD.n1032 VSSD.n1031 34.6358
R7674 VSSD.n1012 VSSD.n934 34.6358
R7675 VSSD.n1013 VSSD.n1012 34.6358
R7676 VSSD.n1014 VSSD.n1013 34.6358
R7677 VSSD.n1014 VSSD.n932 34.6358
R7678 VSSD.n1018 VSSD.n932 34.6358
R7679 VSSD.n999 VSSD.n936 34.6358
R7680 VSSD.n1003 VSSD.n936 34.6358
R7681 VSSD.n1004 VSSD.n1003 34.6358
R7682 VSSD.n1008 VSSD.n1004 34.6358
R7683 VSSD.n996 VSSD.n940 34.6358
R7684 VSSD.n997 VSSD.n996 34.6358
R7685 VSSD.n977 VSSD.n949 34.6358
R7686 VSSD.n978 VSSD.n977 34.6358
R7687 VSSD.n979 VSSD.n978 34.6358
R7688 VSSD.n979 VSSD.n947 34.6358
R7689 VSSD.n983 VSSD.n947 34.6358
R7690 VSSD.n964 VSSD.n951 34.6358
R7691 VSSD.n968 VSSD.n951 34.6358
R7692 VSSD.n969 VSSD.n968 34.6358
R7693 VSSD.n973 VSSD.n969 34.6358
R7694 VSSD.n961 VSSD.n955 34.6358
R7695 VSSD.n962 VSSD.n961 34.6358
R7696 VSSD.n1642 VSSD.n1383 34.2593
R7697 VSSD.n2018 VSSD.n0 33.8829
R7698 VSSD.n1835 VSSD.n109 32.0005
R7699 VSSD.n1311 VSSD.n805 32.0005
R7700 VSSD.t820 VSSD.t985 31.1116
R7701 VSSD.n2014 VSSD.t550 30.9283
R7702 VSSD.n1648 VSSD.n1382 29.7417
R7703 VSSD.n1681 VSSD.n1680 29.7417
R7704 VSSD.n1719 VSSD.n1359 29.7417
R7705 VSSD.n1752 VSSD.n1751 29.7417
R7706 VSSD.n1790 VSSD.n1336 29.7417
R7707 VSSD.n1450 VSSD.n1449 29.7417
R7708 VSSD.n1485 VSSD.n1434 29.7417
R7709 VSSD.n1522 VSSD.n1422 29.7417
R7710 VSSD.n1556 VSSD.n1555 29.7417
R7711 VSSD.n1591 VSSD.n1399 29.7417
R7712 VSSD.n1300 VSSD.n1299 29.7417
R7713 VSSD.n1265 VSSD.n1264 29.7417
R7714 VSSD.n1230 VSSD.n1229 29.7417
R7715 VSSD.n1195 VSSD.n1194 29.7417
R7716 VSSD.n1160 VSSD.n1159 29.7417
R7717 VSSD.n1125 VSSD.n1124 29.7417
R7718 VSSD.n1090 VSSD.n1089 29.7417
R7719 VSSD.n1055 VSSD.n1054 29.7417
R7720 VSSD.n1020 VSSD.n1019 29.7417
R7721 VSSD.n985 VSSD.n984 29.7417
R7722 VSSD.n1844 VSSD.n104 28.9887
R7723 VSSD.n1318 VSSD.n1317 28.9887
R7724 VSSD.n1675 VSSD.n1370 27.4829
R7725 VSSD.n1713 VSSD.n1360 27.4829
R7726 VSSD.n1746 VSSD.n1347 27.4829
R7727 VSSD.n1784 VSSD.n1337 27.4829
R7728 VSSD.n1482 VSSD.n1436 27.4829
R7729 VSSD.n1516 VSSD.n1515 27.4829
R7730 VSSD.n1549 VSSD.n1411 27.4829
R7731 VSSD.n1588 VSSD.n1401 27.4829
R7732 VSSD.n1270 VSSD.n1269 27.4829
R7733 VSSD.n1235 VSSD.n1234 27.4829
R7734 VSSD.n1200 VSSD.n1199 27.4829
R7735 VSSD.n1165 VSSD.n1164 27.4829
R7736 VSSD.n1130 VSSD.n1129 27.4829
R7737 VSSD.n1095 VSSD.n1094 27.4829
R7738 VSSD.n1060 VSSD.n1059 27.4829
R7739 VSSD.n1025 VSSD.n1024 27.4829
R7740 VSSD.n990 VSSD.n989 27.4829
R7741 VSSD.n1622 VSSD.n1621 27.1064
R7742 VSSD.n1851 VSSD.n102 27.1064
R7743 VSSD.t855 VSSD.t458 26.8046
R7744 VSSD.n1831 VSSD.n1830 25.977
R7745 VSSD.n1307 VSSD.n1306 25.977
R7746 VSSD VSSD.n2013 25.7737
R7747 VSSD.t944 VSSD.t851 25.7737
R7748 VSSD.n108 VSSD.t1191 24.9236
R7749 VSSD.n108 VSSD.t860 24.9236
R7750 VSSD.n1836 VSSD.t858 24.9236
R7751 VSSD.n1836 VSSD.t854 24.9236
R7752 VSSD.n106 VSSD.t852 24.9236
R7753 VSSD.n106 VSSD.t549 24.9236
R7754 VSSD.n1843 VSSD.t378 24.9236
R7755 VSSD.n1843 VSSD.t547 24.9236
R7756 VSSD.n1846 VSSD.t376 24.9236
R7757 VSSD.n1846 VSSD.t373 24.9236
R7758 VSSD.n117 VSSD.t793 24.9236
R7759 VSSD.n117 VSSD.t122 24.9236
R7760 VSSD.n475 VSSD.t211 24.9236
R7761 VSSD.n475 VSSD.t1183 24.9236
R7762 VSSD.n476 VSSD.t159 24.9236
R7763 VSSD.n476 VSSD.t1185 24.9236
R7764 VSSD.n479 VSSD.t213 24.9236
R7765 VSSD.n479 VSSD.t414 24.9236
R7766 VSSD.n792 VSSD.t743 24.9236
R7767 VSSD.n792 VSSD.t543 24.9236
R7768 VSSD.n793 VSSD.t419 24.9236
R7769 VSSD.n793 VSSD.t261 24.9236
R7770 VSSD.n794 VSSD.t171 24.9236
R7771 VSSD.n794 VSSD.t542 24.9236
R7772 VSSD.n796 VSSD.t339 24.9236
R7773 VSSD.n796 VSSD.t259 24.9236
R7774 VSSD.n797 VSSD.t192 24.9236
R7775 VSSD.n797 VSSD.t173 24.9236
R7776 VSSD.n798 VSSD.t1193 24.9236
R7777 VSSD.n798 VSSD.t340 24.9236
R7778 VSSD.n801 VSSD.t247 24.9236
R7779 VSSD.n801 VSSD.t194 24.9236
R7780 VSSD.n802 VSSD.t353 24.9236
R7781 VSSD.n802 VSSD.t245 24.9236
R7782 VSSD.n803 VSSD.t720 24.9236
R7783 VSSD.n803 VSSD.t249 24.9236
R7784 VSSD.n804 VSSD.t350 24.9236
R7785 VSSD.n804 VSSD.t354 24.9236
R7786 VSSD.n1673 VSSD.n1373 24.8476
R7787 VSSD.n1708 VSSD.n1707 24.8476
R7788 VSSD.n1744 VSSD.n1350 24.8476
R7789 VSSD.n1779 VSSD.n1778 24.8476
R7790 VSSD.n1815 VSSD.n1327 24.8476
R7791 VSSD.n1477 VSSD.n1476 24.8476
R7792 VSSD.n1511 VSSD.n1510 24.8476
R7793 VSSD.n1547 VSSD.n1413 24.8476
R7794 VSSD.n1583 VSSD.n1582 24.8476
R7795 VSSD.n1617 VSSD.n1616 24.8476
R7796 VSSD.n1272 VSSD.n820 24.8476
R7797 VSSD.n1237 VSSD.n835 24.8476
R7798 VSSD.n1202 VSSD.n850 24.8476
R7799 VSSD.n1167 VSSD.n865 24.8476
R7800 VSSD.n1132 VSSD.n880 24.8476
R7801 VSSD.n1097 VSSD.n895 24.8476
R7802 VSSD.n1062 VSSD.n910 24.8476
R7803 VSSD.n1027 VSSD.n925 24.8476
R7804 VSSD.n992 VSSD.n940 24.8476
R7805 VSSD.n957 VSSD.n955 24.8476
R7806 VSSD.n2015 VSSD 24.8153
R7807 VSSD VSSD.t820 24.0746
R7808 VSSD.n1644 VSSD.n1382 22.9652
R7809 VSSD.n1675 VSSD.n1674 22.9652
R7810 VSSD.n1680 VSSD.n1679 22.9652
R7811 VSSD.n1709 VSSD.n1360 22.9652
R7812 VSSD.n1715 VSSD.n1359 22.9652
R7813 VSSD.n1746 VSSD.n1745 22.9652
R7814 VSSD.n1751 VSSD.n1750 22.9652
R7815 VSSD.n1780 VSSD.n1337 22.9652
R7816 VSSD.n1786 VSSD.n1336 22.9652
R7817 VSSD.n1817 VSSD.n1816 22.9652
R7818 VSSD.n1449 VSSD.n1448 22.9652
R7819 VSSD.n1478 VSSD.n1436 22.9652
R7820 VSSD.n1485 VSSD.n1484 22.9652
R7821 VSSD.n1515 VSSD.n1424 22.9652
R7822 VSSD.n1518 VSSD.n1422 22.9652
R7823 VSSD.n1549 VSSD.n1548 22.9652
R7824 VSSD.n1555 VSSD.n1554 22.9652
R7825 VSSD.n1584 VSSD.n1401 22.9652
R7826 VSSD.n1591 VSSD.n1590 22.9652
R7827 VSSD.n1621 VSSD.n1389 22.9652
R7828 VSSD.n1847 VSSD.n1845 22.9652
R7829 VSSD.n1320 VSSD.n1319 22.9652
R7830 VSSD.n1301 VSSD.n1300 22.9652
R7831 VSSD.n1271 VSSD.n1270 22.9652
R7832 VSSD.n1265 VSSD.n825 22.9652
R7833 VSSD.n1236 VSSD.n1235 22.9652
R7834 VSSD.n1230 VSSD.n840 22.9652
R7835 VSSD.n1201 VSSD.n1200 22.9652
R7836 VSSD.n1195 VSSD.n855 22.9652
R7837 VSSD.n1166 VSSD.n1165 22.9652
R7838 VSSD.n1160 VSSD.n870 22.9652
R7839 VSSD.n1131 VSSD.n1130 22.9652
R7840 VSSD.n1125 VSSD.n885 22.9652
R7841 VSSD.n1096 VSSD.n1095 22.9652
R7842 VSSD.n1090 VSSD.n900 22.9652
R7843 VSSD.n1061 VSSD.n1060 22.9652
R7844 VSSD.n1055 VSSD.n915 22.9652
R7845 VSSD.n1026 VSSD.n1025 22.9652
R7846 VSSD.n1020 VSSD.n930 22.9652
R7847 VSSD.n991 VSSD.n990 22.9652
R7848 VSSD.n985 VSSD.n945 22.9652
R7849 VSSD.t375 VSSD.t1162 22.6809
R7850 VSSD.t372 VSSD.t184 22.6809
R7851 VSSD.n1636 VSSD.t456 22.3257
R7852 VSSD.n1387 VSSD.t875 22.3257
R7853 VSSD.n1644 VSSD.n1642 21.4593
R7854 VSSD.n1674 VSSD.n1673 21.4593
R7855 VSSD.n1679 VSSD.n1370 21.4593
R7856 VSSD.n1709 VSSD.n1708 21.4593
R7857 VSSD.n1715 VSSD.n1713 21.4593
R7858 VSSD.n1745 VSSD.n1744 21.4593
R7859 VSSD.n1750 VSSD.n1347 21.4593
R7860 VSSD.n1780 VSSD.n1779 21.4593
R7861 VSSD.n1786 VSSD.n1784 21.4593
R7862 VSSD.n1816 VSSD.n1815 21.4593
R7863 VSSD.n1478 VSSD.n1477 21.4593
R7864 VSSD.n1484 VSSD.n1482 21.4593
R7865 VSSD.n1511 VSSD.n1424 21.4593
R7866 VSSD.n1518 VSSD.n1516 21.4593
R7867 VSSD.n1548 VSSD.n1547 21.4593
R7868 VSSD.n1554 VSSD.n1411 21.4593
R7869 VSSD.n1584 VSSD.n1583 21.4593
R7870 VSSD.n1590 VSSD.n1588 21.4593
R7871 VSSD.n1617 VSSD.n1389 21.4593
R7872 VSSD.n1847 VSSD.n102 21.4593
R7873 VSSD.n1320 VSSD.n0 21.4593
R7874 VSSD.n1301 VSSD.n807 21.4593
R7875 VSSD.n1272 VSSD.n1271 21.4593
R7876 VSSD.n1269 VSSD.n825 21.4593
R7877 VSSD.n1237 VSSD.n1236 21.4593
R7878 VSSD.n1234 VSSD.n840 21.4593
R7879 VSSD.n1202 VSSD.n1201 21.4593
R7880 VSSD.n1199 VSSD.n855 21.4593
R7881 VSSD.n1167 VSSD.n1166 21.4593
R7882 VSSD.n1164 VSSD.n870 21.4593
R7883 VSSD.n1132 VSSD.n1131 21.4593
R7884 VSSD.n1129 VSSD.n885 21.4593
R7885 VSSD.n1097 VSSD.n1096 21.4593
R7886 VSSD.n1094 VSSD.n900 21.4593
R7887 VSSD.n1062 VSSD.n1061 21.4593
R7888 VSSD.n1059 VSSD.n915 21.4593
R7889 VSSD.n1027 VSSD.n1026 21.4593
R7890 VSSD.n1024 VSSD.n930 21.4593
R7891 VSSD.n992 VSSD.n991 21.4593
R7892 VSSD.n989 VSSD.n945 21.4593
R7893 VSSD.n260 VSSD.n259 20.5251
R7894 VSSD.n658 VSSD.n657 20.5251
R7895 VSSD.n1980 VSSD.n1979 20.3299
R7896 VSSD.n1949 VSSD.n1948 20.3299
R7897 VSSD.n1918 VSSD.n1917 20.3299
R7898 VSSD.n1887 VSSD.n1886 20.3299
R7899 VSSD.n1854 VSSD.n100 19.9534
R7900 VSSD.n1881 VSSD.n88 19.9534
R7901 VSSD.n2008 VSSD.n2007 19.9534
R7902 VSSD.n1982 VSSD.n20 19.9534
R7903 VSSD.n1977 VSSD.n1976 19.9534
R7904 VSSD.n1951 VSSD.n41 19.9534
R7905 VSSD.n1946 VSSD.n1945 19.9534
R7906 VSSD.n1920 VSSD.n62 19.9534
R7907 VSSD.n1915 VSSD.n1914 19.9534
R7908 VSSD.n1889 VSSD.n83 19.9534
R7909 VSSD.n1825 VSSD 19.5877
R7910 VSSD.n1819 VSSD 19.5539
R7911 VSSD VSSD.n1828 18.8091
R7912 VSSD.t381 VSSD.t546 18.5572
R7913 VSSD.t930 VSSD.t853 18.5572
R7914 VSSD.n1306 VSSD.n1305 18.4476
R7915 VSSD.n469 VSSD.n468 18.1174
R7916 VSSD.n463 VSSD.n462 18.1174
R7917 VSSD.n462 VSSD.n163 18.1174
R7918 VSSD.n458 VSSD.n163 18.1174
R7919 VSSD.n456 VSSD.n455 18.1174
R7920 VSSD.n455 VSSD.n166 18.1174
R7921 VSSD.n451 VSSD.n166 18.1174
R7922 VSSD.n451 VSSD.n450 18.1174
R7923 VSSD.n448 VSSD.n169 18.1174
R7924 VSSD.n444 VSSD.n169 18.1174
R7925 VSSD.n444 VSSD.n443 18.1174
R7926 VSSD.n443 VSSD.n442 18.1174
R7927 VSSD.n442 VSSD.n171 18.1174
R7928 VSSD.n434 VSSD.n175 18.1174
R7929 VSSD.n428 VSSD.n427 18.1174
R7930 VSSD.n427 VSSD.n179 18.1174
R7931 VSSD.n423 VSSD.n179 18.1174
R7932 VSSD.n421 VSSD.n420 18.1174
R7933 VSSD.n420 VSSD.n182 18.1174
R7934 VSSD.n416 VSSD.n182 18.1174
R7935 VSSD.n416 VSSD.n415 18.1174
R7936 VSSD.n413 VSSD.n185 18.1174
R7937 VSSD.n409 VSSD.n185 18.1174
R7938 VSSD.n409 VSSD.n408 18.1174
R7939 VSSD.n408 VSSD.n407 18.1174
R7940 VSSD.n407 VSSD.n187 18.1174
R7941 VSSD.n399 VSSD.n191 18.1174
R7942 VSSD.n393 VSSD.n392 18.1174
R7943 VSSD.n392 VSSD.n195 18.1174
R7944 VSSD.n388 VSSD.n195 18.1174
R7945 VSSD.n386 VSSD.n385 18.1174
R7946 VSSD.n385 VSSD.n198 18.1174
R7947 VSSD.n381 VSSD.n198 18.1174
R7948 VSSD.n381 VSSD.n380 18.1174
R7949 VSSD.n378 VSSD.n201 18.1174
R7950 VSSD.n374 VSSD.n201 18.1174
R7951 VSSD.n374 VSSD.n373 18.1174
R7952 VSSD.n373 VSSD.n372 18.1174
R7953 VSSD.n372 VSSD.n203 18.1174
R7954 VSSD.n364 VSSD.n210 18.1174
R7955 VSSD.n358 VSSD.n357 18.1174
R7956 VSSD.n357 VSSD.n214 18.1174
R7957 VSSD.n353 VSSD.n214 18.1174
R7958 VSSD.n351 VSSD.n350 18.1174
R7959 VSSD.n350 VSSD.n217 18.1174
R7960 VSSD.n346 VSSD.n217 18.1174
R7961 VSSD.n346 VSSD.n345 18.1174
R7962 VSSD.n343 VSSD.n220 18.1174
R7963 VSSD.n339 VSSD.n220 18.1174
R7964 VSSD.n339 VSSD.n338 18.1174
R7965 VSSD.n338 VSSD.n337 18.1174
R7966 VSSD.n337 VSSD.n222 18.1174
R7967 VSSD.n329 VSSD.n226 18.1174
R7968 VSSD.n323 VSSD.n322 18.1174
R7969 VSSD.n322 VSSD.n230 18.1174
R7970 VSSD.n318 VSSD.n230 18.1174
R7971 VSSD.n316 VSSD.n315 18.1174
R7972 VSSD.n315 VSSD.n233 18.1174
R7973 VSSD.n311 VSSD.n233 18.1174
R7974 VSSD.n311 VSSD.n310 18.1174
R7975 VSSD.n308 VSSD.n236 18.1174
R7976 VSSD.n304 VSSD.n236 18.1174
R7977 VSSD.n304 VSSD.n303 18.1174
R7978 VSSD.n303 VSSD.n302 18.1174
R7979 VSSD.n302 VSSD.n238 18.1174
R7980 VSSD.n294 VSSD.n242 18.1174
R7981 VSSD.n288 VSSD.n287 18.1174
R7982 VSSD.n287 VSSD.n246 18.1174
R7983 VSSD.n283 VSSD.n246 18.1174
R7984 VSSD.n281 VSSD.n280 18.1174
R7985 VSSD.n280 VSSD.n249 18.1174
R7986 VSSD.n276 VSSD.n249 18.1174
R7987 VSSD.n276 VSSD.n275 18.1174
R7988 VSSD.n273 VSSD.n252 18.1174
R7989 VSSD.n269 VSSD.n252 18.1174
R7990 VSSD.n269 VSSD.n268 18.1174
R7991 VSSD.n268 VSSD.n267 18.1174
R7992 VSSD.n267 VSSD.n254 18.1174
R7993 VSSD.n492 VSSD.n491 18.1174
R7994 VSSD.n488 VSSD.n487 18.1174
R7995 VSSD.n482 VSSD.n481 18.1174
R7996 VSSD.n772 VSSD.n771 18.1174
R7997 VSSD.n776 VSSD.n775 18.1174
R7998 VSSD.n778 VSSD.n776 18.1174
R7999 VSSD.n782 VSSD.n115 18.1174
R8000 VSSD.n501 VSSD.n500 18.1174
R8001 VSSD.n501 VSSD.n157 18.1174
R8002 VSSD.n505 VSSD.n157 18.1174
R8003 VSSD.n508 VSSD.n507 18.1174
R8004 VSSD.n508 VSSD.n154 18.1174
R8005 VSSD.n512 VSSD.n154 18.1174
R8006 VSSD.n513 VSSD.n512 18.1174
R8007 VSSD.n516 VSSD.n152 18.1174
R8008 VSSD.n520 VSSD.n152 18.1174
R8009 VSSD.n521 VSSD.n520 18.1174
R8010 VSSD.n522 VSSD.n521 18.1174
R8011 VSSD.n522 VSSD.n150 18.1174
R8012 VSSD.n534 VSSD.n147 18.1174
R8013 VSSD.n538 VSSD.n145 18.1174
R8014 VSSD.n542 VSSD.n145 18.1174
R8015 VSSD.n543 VSSD.n542 18.1174
R8016 VSSD.n545 VSSD.n142 18.1174
R8017 VSSD.n549 VSSD.n142 18.1174
R8018 VSSD.n550 VSSD.n549 18.1174
R8019 VSSD.n553 VSSD.n550 18.1174
R8020 VSSD.n557 VSSD.n140 18.1174
R8021 VSSD.n558 VSSD.n557 18.1174
R8022 VSSD.n559 VSSD.n558 18.1174
R8023 VSSD.n559 VSSD.n138 18.1174
R8024 VSSD.n563 VSSD.n138 18.1174
R8025 VSSD.n573 VSSD.n572 18.1174
R8026 VSSD.n579 VSSD.n578 18.1174
R8027 VSSD.n579 VSSD.n133 18.1174
R8028 VSSD.n583 VSSD.n133 18.1174
R8029 VSSD.n586 VSSD.n585 18.1174
R8030 VSSD.n586 VSSD.n130 18.1174
R8031 VSSD.n590 VSSD.n130 18.1174
R8032 VSSD.n591 VSSD.n590 18.1174
R8033 VSSD.n594 VSSD.n128 18.1174
R8034 VSSD.n598 VSSD.n128 18.1174
R8035 VSSD.n599 VSSD.n598 18.1174
R8036 VSSD.n600 VSSD.n599 18.1174
R8037 VSSD.n600 VSSD.n126 18.1174
R8038 VSSD.n756 VSSD.n755 18.1174
R8039 VSSD.n755 VSSD.n612 18.1174
R8040 VSSD.n751 VSSD.n612 18.1174
R8041 VSSD.n749 VSSD.n748 18.1174
R8042 VSSD.n748 VSSD.n615 18.1174
R8043 VSSD.n744 VSSD.n615 18.1174
R8044 VSSD.n744 VSSD.n743 18.1174
R8045 VSSD.n741 VSSD.n618 18.1174
R8046 VSSD.n737 VSSD.n618 18.1174
R8047 VSSD.n737 VSSD.n736 18.1174
R8048 VSSD.n736 VSSD.n735 18.1174
R8049 VSSD.n735 VSSD.n620 18.1174
R8050 VSSD.n727 VSSD.n624 18.1174
R8051 VSSD.n721 VSSD.n720 18.1174
R8052 VSSD.n720 VSSD.n628 18.1174
R8053 VSSD.n716 VSSD.n628 18.1174
R8054 VSSD.n714 VSSD.n713 18.1174
R8055 VSSD.n713 VSSD.n631 18.1174
R8056 VSSD.n709 VSSD.n631 18.1174
R8057 VSSD.n709 VSSD.n708 18.1174
R8058 VSSD.n706 VSSD.n634 18.1174
R8059 VSSD.n702 VSSD.n634 18.1174
R8060 VSSD.n702 VSSD.n701 18.1174
R8061 VSSD.n701 VSSD.n700 18.1174
R8062 VSSD.n700 VSSD.n636 18.1174
R8063 VSSD.n692 VSSD.n640 18.1174
R8064 VSSD.n686 VSSD.n685 18.1174
R8065 VSSD.n685 VSSD.n644 18.1174
R8066 VSSD.n681 VSSD.n644 18.1174
R8067 VSSD.n679 VSSD.n678 18.1174
R8068 VSSD.n678 VSSD.n647 18.1174
R8069 VSSD.n674 VSSD.n647 18.1174
R8070 VSSD.n674 VSSD.n673 18.1174
R8071 VSSD.n671 VSSD.n650 18.1174
R8072 VSSD.n667 VSSD.n650 18.1174
R8073 VSSD.n667 VSSD.n666 18.1174
R8074 VSSD.n666 VSSD.n665 18.1174
R8075 VSSD.n665 VSSD.n652 18.1174
R8076 VSSD.n785 VSSD.n784 17.7236
R8077 VSSD.n1668 VSSD.n1667 17.6946
R8078 VSSD.n1703 VSSD.n1702 17.6946
R8079 VSSD.n1739 VSSD.n1738 17.6946
R8080 VSSD.n1774 VSSD.n1773 17.6946
R8081 VSSD.n1810 VSSD.n1809 17.6946
R8082 VSSD.n1472 VSSD.n1471 17.6946
R8083 VSSD.n1429 VSSD.n1426 17.6946
R8084 VSSD.n1542 VSSD.n1541 17.6946
R8085 VSSD.n1578 VSSD.n1577 17.6946
R8086 VSSD.n1394 VSSD.n1391 17.6946
R8087 VSSD.n1861 VSSD.n1859 17.6946
R8088 VSSD.n1879 VSSD.n92 17.6946
R8089 VSSD.n11 VSSD.n8 17.6946
R8090 VSSD.n1988 VSSD.n1987 17.6946
R8091 VSSD.n32 VSSD.n29 17.6946
R8092 VSSD.n1957 VSSD.n1956 17.6946
R8093 VSSD.n53 VSSD.n50 17.6946
R8094 VSSD.n1926 VSSD.n1925 17.6946
R8095 VSSD.n74 VSSD.n71 17.6946
R8096 VSSD.n1895 VSSD.n1894 17.6946
R8097 VSSD.n1278 VSSD.n1277 17.6946
R8098 VSSD.n1243 VSSD.n1242 17.6946
R8099 VSSD.n1208 VSSD.n1207 17.6946
R8100 VSSD.n1173 VSSD.n1172 17.6946
R8101 VSSD.n1138 VSSD.n1137 17.6946
R8102 VSSD.n1103 VSSD.n1102 17.6946
R8103 VSSD.n1068 VSSD.n1067 17.6946
R8104 VSSD.n1033 VSSD.n1032 17.6946
R8105 VSSD.n998 VSSD.n997 17.6946
R8106 VSSD.n963 VSSD.n962 17.6946
R8107 VSSD.n787 VSSD 17.5031
R8108 VSSD.n465 VSSD.n464 17.3297
R8109 VSSD.n430 VSSD.n429 17.3297
R8110 VSSD.n395 VSSD.n394 17.3297
R8111 VSSD.n360 VSSD.n359 17.3297
R8112 VSSD.n325 VSSD.n324 17.3297
R8113 VSSD.n290 VSSD.n289 17.3297
R8114 VSSD.n784 VSSD.n783 17.3297
R8115 VSSD.n499 VSSD.n498 17.3297
R8116 VSSD.n537 VSSD.n536 17.3297
R8117 VSSD.n577 VSSD.n576 17.3297
R8118 VSSD.n758 VSSD.n757 17.3297
R8119 VSSD.n723 VSSD.n722 17.3297
R8120 VSSD.n688 VSSD.n687 17.3297
R8121 VSSD.n471 VSSD.n160 16.9659
R8122 VSSD.n494 VSSD.n472 16.9659
R8123 VSSD.n465 VSSD.n161 16.9359
R8124 VSSD.n430 VSSD.n178 16.9359
R8125 VSSD.n395 VSSD.n194 16.9359
R8126 VSSD.n360 VSSD.n213 16.9359
R8127 VSSD.n325 VSSD.n229 16.9359
R8128 VSSD.n290 VSSD.n245 16.9359
R8129 VSSD.n778 VSSD.n777 16.9359
R8130 VSSD.n498 VSSD.n159 16.9359
R8131 VSSD.n536 VSSD.n535 16.9359
R8132 VSSD.n576 VSSD.n135 16.9359
R8133 VSSD.n758 VSSD.n123 16.9359
R8134 VSSD.n723 VSSD.n627 16.9359
R8135 VSSD.n688 VSSD.n643 16.9359
R8136 VSSD.n485 VSSD.n477 16.739
R8137 VSSD.n775 VSSD.n118 16.542
R8138 VSSD.n486 VSSD.n485 16.3451
R8139 VSSD.n488 VSSD.n473 15.7543
R8140 VSSD.n437 VSSD.n436 15.5574
R8141 VSSD.n402 VSSD.n401 15.5574
R8142 VSSD.n367 VSSD.n366 15.5574
R8143 VSSD.n332 VSSD.n331 15.5574
R8144 VSSD.n297 VSSD.n296 15.5574
R8145 VSSD.n262 VSSD.n261 15.5574
R8146 VSSD.n528 VSSD.n527 15.5574
R8147 VSSD.n566 VSSD.n565 15.5574
R8148 VSSD.n606 VSSD.n605 15.5574
R8149 VSSD.n730 VSSD.n729 15.5574
R8150 VSSD.n695 VSSD.n694 15.5574
R8151 VSSD.n660 VSSD.n659 15.5574
R8152 VSSD.n1845 VSSD.n1844 15.4358
R8153 VSSD.n1319 VSSD.n1318 15.4358
R8154 VSSD.n1649 VSSD.n1648 14.6829
R8155 VSSD.n1681 VSSD.n1368 14.6829
R8156 VSSD.n1720 VSSD.n1719 14.6829
R8157 VSSD.n1752 VSSD.n1345 14.6829
R8158 VSSD.n1791 VSSD.n1790 14.6829
R8159 VSSD.n1450 VSSD.n1444 14.6829
R8160 VSSD.n1489 VSSD.n1434 14.6829
R8161 VSSD.n1523 VSSD.n1522 14.6829
R8162 VSSD.n1556 VSSD.n1409 14.6829
R8163 VSSD.n1595 VSSD.n1399 14.6829
R8164 VSSD.n1858 VSSD.n100 14.6829
R8165 VSSD.n1881 VSSD.n1880 14.6829
R8166 VSSD.n2007 VSSD.n2006 14.6829
R8167 VSSD.n1986 VSSD.n20 14.6829
R8168 VSSD.n1976 VSSD.n1975 14.6829
R8169 VSSD.n1955 VSSD.n41 14.6829
R8170 VSSD.n1945 VSSD.n1944 14.6829
R8171 VSSD.n1924 VSSD.n62 14.6829
R8172 VSSD.n1914 VSSD.n1913 14.6829
R8173 VSSD.n1893 VSSD.n83 14.6829
R8174 VSSD.n1299 VSSD.n1298 14.6829
R8175 VSSD.n1264 VSSD.n1263 14.6829
R8176 VSSD.n1229 VSSD.n1228 14.6829
R8177 VSSD.n1194 VSSD.n1193 14.6829
R8178 VSSD.n1159 VSSD.n1158 14.6829
R8179 VSSD.n1124 VSSD.n1123 14.6829
R8180 VSSD.n1089 VSSD.n1088 14.6829
R8181 VSSD.n1054 VSSD.n1053 14.6829
R8182 VSSD.n1019 VSSD.n1018 14.6829
R8183 VSSD.n984 VSSD.n983 14.6829
R8184 VSSD.n481 VSSD.n480 13.5882
R8185 VSSD.n458 VSSD.n457 12.9974
R8186 VSSD.n423 VSSD.n422 12.9974
R8187 VSSD.n388 VSSD.n387 12.9974
R8188 VSSD.n353 VSSD.n352 12.9974
R8189 VSSD.n318 VSSD.n317 12.9974
R8190 VSSD.n283 VSSD.n282 12.9974
R8191 VSSD.n506 VSSD.n505 12.9974
R8192 VSSD.n544 VSSD.n543 12.9974
R8193 VSSD.n584 VSSD.n583 12.9974
R8194 VSSD.n751 VSSD.n750 12.9974
R8195 VSSD.n716 VSSD.n715 12.9974
R8196 VSSD.n681 VSSD.n680 12.9974
R8197 VSSD.n1831 VSSD.n109 12.424
R8198 VSSD.n1307 VSSD.n805 12.424
R8199 VSSD.n768 VSSD.n119 12.2097
R8200 VSSD.n436 VSSD.n435 12.0128
R8201 VSSD.n401 VSSD.n400 12.0128
R8202 VSSD.n366 VSSD.n365 12.0128
R8203 VSSD.n331 VSSD.n330 12.0128
R8204 VSSD.n296 VSSD.n295 12.0128
R8205 VSSD.n261 VSSD.n260 12.0128
R8206 VSSD.n767 VSSD.n121 12.0128
R8207 VSSD.n529 VSSD.n528 12.0128
R8208 VSSD.n566 VSSD.n136 12.0128
R8209 VSSD.n607 VSSD.n606 12.0128
R8210 VSSD.n729 VSSD.n728 12.0128
R8211 VSSD.n694 VSSD.n693 12.0128
R8212 VSSD.n659 VSSD.n658 12.0128
R8213 VSSD.n495 VSSD.n494 11.4222
R8214 VSSD.n435 VSSD.n434 11.2251
R8215 VSSD.n400 VSSD.n399 11.2251
R8216 VSSD.n365 VSSD.n364 11.2251
R8217 VSSD.n330 VSSD.n329 11.2251
R8218 VSSD.n295 VSSD.n294 11.2251
R8219 VSSD.n529 VSSD.n147 11.2251
R8220 VSSD.n572 VSSD.n136 11.2251
R8221 VSSD.n607 VSSD.n122 11.2251
R8222 VSSD.n728 VSSD.n727 11.2251
R8223 VSSD.n693 VSSD.n692 11.2251
R8224 VSSD.n1324 VSSD.n1323 11.0366
R8225 VSSD.n496 VSSD.n159 10.482
R8226 VSSD.n1853 VSSD.n1851 9.78874
R8227 VSSD.n1854 VSSD.n1853 9.78874
R8228 VSSD.n2010 VSSD.n2009 9.78874
R8229 VSSD.n2009 VSSD.n2008 9.78874
R8230 VSSD.n1982 VSSD.n1981 9.78874
R8231 VSSD.n1981 VSSD.n1980 9.78874
R8232 VSSD.n1979 VSSD.n1978 9.78874
R8233 VSSD.n1978 VSSD.n1977 9.78874
R8234 VSSD.n1951 VSSD.n1950 9.78874
R8235 VSSD.n1950 VSSD.n1949 9.78874
R8236 VSSD.n1948 VSSD.n1947 9.78874
R8237 VSSD.n1947 VSSD.n1946 9.78874
R8238 VSSD.n1920 VSSD.n1919 9.78874
R8239 VSSD.n1919 VSSD.n1918 9.78874
R8240 VSSD.n1917 VSSD.n1916 9.78874
R8241 VSSD.n1916 VSSD.n1915 9.78874
R8242 VSSD.n1889 VSSD.n1888 9.78874
R8243 VSSD.n1888 VSSD.n1887 9.78874
R8244 VSSD.n1886 VSSD.n1885 9.78874
R8245 VSSD.n1885 VSSD.n88 9.78874
R8246 VSSD.n786 VSSD.n785 9.69435
R8247 VSSD.n365 VSSD.n209 9.63373
R8248 VSSD.n1638 VSSD.n1637 9.41227
R8249 VSSD.n1623 VSSD.n1388 9.41227
R8250 VSSD.n107 VSSD.n104 9.41227
R8251 VSSD.n1317 VSSD.n799 9.41227
R8252 VSSD VSSD.n2018 9.35779
R8253 VSSD.n1885 VSSD.n1884 9.3005
R8254 VSSD.n1855 VSSD.n1854 9.3005
R8255 VSSD.n1851 VSSD.n1850 9.3005
R8256 VSSD.n1848 VSSD.n1847 9.3005
R8257 VSSD.n1832 VSSD.n1831 9.3005
R8258 VSSD.n1833 VSSD.n109 9.3005
R8259 VSSD.n1835 VSSD.n1834 9.3005
R8260 VSSD.n1838 VSSD.n105 9.3005
R8261 VSSD.n1840 VSSD.n1839 9.3005
R8262 VSSD.n1841 VSSD.n104 9.3005
R8263 VSSD.n1844 VSSD.n1842 9.3005
R8264 VSSD.n1845 VSSD.n103 9.3005
R8265 VSSD.n1849 VSSD.n102 9.3005
R8266 VSSD.n1853 VSSD.n101 9.3005
R8267 VSSD.n1856 VSSD.n100 9.3005
R8268 VSSD.n1858 VSSD.n1857 9.3005
R8269 VSSD.n1859 VSSD.n99 9.3005
R8270 VSSD.n1863 VSSD.n1862 9.3005
R8271 VSSD.n1864 VSSD.n98 9.3005
R8272 VSSD.n1866 VSSD.n1865 9.3005
R8273 VSSD.n1867 VSSD.n95 9.3005
R8274 VSSD.n1871 VSSD.n1870 9.3005
R8275 VSSD.n1872 VSSD.n94 9.3005
R8276 VSSD.n1874 VSSD.n1873 9.3005
R8277 VSSD.n1875 VSSD.n93 9.3005
R8278 VSSD.n1877 VSSD.n1876 9.3005
R8279 VSSD.n1879 VSSD.n1878 9.3005
R8280 VSSD.n1880 VSSD.n90 9.3005
R8281 VSSD.n1882 VSSD.n1881 9.3005
R8282 VSSD.n1883 VSSD.n88 9.3005
R8283 VSSD.n1886 VSSD.n87 9.3005
R8284 VSSD.n2011 VSSD.n2010 9.3005
R8285 VSSD.n2009 VSSD.n4 9.3005
R8286 VSSD.n2008 VSSD.n6 9.3005
R8287 VSSD.n2007 VSSD.n7 9.3005
R8288 VSSD.n2006 VSSD.n2005 9.3005
R8289 VSSD.n2004 VSSD.n8 9.3005
R8290 VSSD.n2003 VSSD.n2002 9.3005
R8291 VSSD.n2001 VSSD.n9 9.3005
R8292 VSSD.n2000 VSSD.n1999 9.3005
R8293 VSSD.n1998 VSSD.n12 9.3005
R8294 VSSD.n1997 VSSD.n1996 9.3005
R8295 VSSD.n1994 VSSD.n13 9.3005
R8296 VSSD.n1993 VSSD.n1992 9.3005
R8297 VSSD.n1991 VSSD.n17 9.3005
R8298 VSSD.n1990 VSSD.n1989 9.3005
R8299 VSSD.n1987 VSSD.n18 9.3005
R8300 VSSD.n1986 VSSD.n1985 9.3005
R8301 VSSD.n1984 VSSD.n20 9.3005
R8302 VSSD.n1983 VSSD.n1982 9.3005
R8303 VSSD.n1981 VSSD.n21 9.3005
R8304 VSSD.n1980 VSSD.n23 9.3005
R8305 VSSD.n1979 VSSD.n24 9.3005
R8306 VSSD.n1978 VSSD.n25 9.3005
R8307 VSSD.n1977 VSSD.n27 9.3005
R8308 VSSD.n1976 VSSD.n28 9.3005
R8309 VSSD.n1975 VSSD.n1974 9.3005
R8310 VSSD.n1973 VSSD.n29 9.3005
R8311 VSSD.n1972 VSSD.n1971 9.3005
R8312 VSSD.n1970 VSSD.n30 9.3005
R8313 VSSD.n1969 VSSD.n1968 9.3005
R8314 VSSD.n1967 VSSD.n33 9.3005
R8315 VSSD.n1966 VSSD.n1965 9.3005
R8316 VSSD.n1963 VSSD.n34 9.3005
R8317 VSSD.n1962 VSSD.n1961 9.3005
R8318 VSSD.n1960 VSSD.n38 9.3005
R8319 VSSD.n1959 VSSD.n1958 9.3005
R8320 VSSD.n1956 VSSD.n39 9.3005
R8321 VSSD.n1955 VSSD.n1954 9.3005
R8322 VSSD.n1953 VSSD.n41 9.3005
R8323 VSSD.n1952 VSSD.n1951 9.3005
R8324 VSSD.n1950 VSSD.n42 9.3005
R8325 VSSD.n1949 VSSD.n44 9.3005
R8326 VSSD.n1948 VSSD.n45 9.3005
R8327 VSSD.n1947 VSSD.n46 9.3005
R8328 VSSD.n1946 VSSD.n48 9.3005
R8329 VSSD.n1945 VSSD.n49 9.3005
R8330 VSSD.n1944 VSSD.n1943 9.3005
R8331 VSSD.n1942 VSSD.n50 9.3005
R8332 VSSD.n1941 VSSD.n1940 9.3005
R8333 VSSD.n1939 VSSD.n51 9.3005
R8334 VSSD.n1938 VSSD.n1937 9.3005
R8335 VSSD.n1936 VSSD.n54 9.3005
R8336 VSSD.n1935 VSSD.n1934 9.3005
R8337 VSSD.n1932 VSSD.n55 9.3005
R8338 VSSD.n1931 VSSD.n1930 9.3005
R8339 VSSD.n1929 VSSD.n59 9.3005
R8340 VSSD.n1928 VSSD.n1927 9.3005
R8341 VSSD.n1925 VSSD.n60 9.3005
R8342 VSSD.n1924 VSSD.n1923 9.3005
R8343 VSSD.n1922 VSSD.n62 9.3005
R8344 VSSD.n1921 VSSD.n1920 9.3005
R8345 VSSD.n1919 VSSD.n63 9.3005
R8346 VSSD.n1918 VSSD.n65 9.3005
R8347 VSSD.n1917 VSSD.n66 9.3005
R8348 VSSD.n1916 VSSD.n67 9.3005
R8349 VSSD.n1915 VSSD.n69 9.3005
R8350 VSSD.n1914 VSSD.n70 9.3005
R8351 VSSD.n1913 VSSD.n1912 9.3005
R8352 VSSD.n1911 VSSD.n71 9.3005
R8353 VSSD.n1910 VSSD.n1909 9.3005
R8354 VSSD.n1908 VSSD.n72 9.3005
R8355 VSSD.n1907 VSSD.n1906 9.3005
R8356 VSSD.n1905 VSSD.n75 9.3005
R8357 VSSD.n1904 VSSD.n1903 9.3005
R8358 VSSD.n1901 VSSD.n76 9.3005
R8359 VSSD.n1900 VSSD.n1899 9.3005
R8360 VSSD.n1898 VSSD.n80 9.3005
R8361 VSSD.n1897 VSSD.n1896 9.3005
R8362 VSSD.n1894 VSSD.n81 9.3005
R8363 VSSD.n1893 VSSD.n1892 9.3005
R8364 VSSD.n1891 VSSD.n83 9.3005
R8365 VSSD.n1890 VSSD.n1889 9.3005
R8366 VSSD.n1888 VSSD.n84 9.3005
R8367 VSSD.n1887 VSSD.n86 9.3005
R8368 VSSD.n258 VSSD.n257 9.3005
R8369 VSSD.n261 VSSD.n255 9.3005
R8370 VSSD.n264 VSSD.n263 9.3005
R8371 VSSD.n265 VSSD.n254 9.3005
R8372 VSSD.n267 VSSD.n266 9.3005
R8373 VSSD.n268 VSSD.n253 9.3005
R8374 VSSD.n270 VSSD.n269 9.3005
R8375 VSSD.n271 VSSD.n252 9.3005
R8376 VSSD.n273 VSSD.n272 9.3005
R8377 VSSD.n275 VSSD.n250 9.3005
R8378 VSSD.n277 VSSD.n276 9.3005
R8379 VSSD.n278 VSSD.n249 9.3005
R8380 VSSD.n280 VSSD.n279 9.3005
R8381 VSSD.n281 VSSD.n247 9.3005
R8382 VSSD.n284 VSSD.n283 9.3005
R8383 VSSD.n285 VSSD.n246 9.3005
R8384 VSSD.n287 VSSD.n286 9.3005
R8385 VSSD.n288 VSSD.n244 9.3005
R8386 VSSD.n291 VSSD.n290 9.3005
R8387 VSSD.n292 VSSD.n242 9.3005
R8388 VSSD.n470 VSSD.n469 9.3005
R8389 VSSD.n468 VSSD.n467 9.3005
R8390 VSSD.n466 VSSD.n465 9.3005
R8391 VSSD.n463 VSSD.n162 9.3005
R8392 VSSD.n462 VSSD.n461 9.3005
R8393 VSSD.n460 VSSD.n163 9.3005
R8394 VSSD.n459 VSSD.n458 9.3005
R8395 VSSD.n456 VSSD.n164 9.3005
R8396 VSSD.n455 VSSD.n454 9.3005
R8397 VSSD.n453 VSSD.n166 9.3005
R8398 VSSD.n452 VSSD.n451 9.3005
R8399 VSSD.n450 VSSD.n167 9.3005
R8400 VSSD.n448 VSSD.n447 9.3005
R8401 VSSD.n446 VSSD.n169 9.3005
R8402 VSSD.n445 VSSD.n444 9.3005
R8403 VSSD.n443 VSSD.n170 9.3005
R8404 VSSD.n442 VSSD.n441 9.3005
R8405 VSSD.n440 VSSD.n171 9.3005
R8406 VSSD.n439 VSSD.n438 9.3005
R8407 VSSD.n436 VSSD.n172 9.3005
R8408 VSSD.n176 VSSD.n174 9.3005
R8409 VSSD.n434 VSSD.n433 9.3005
R8410 VSSD.n432 VSSD.n175 9.3005
R8411 VSSD.n431 VSSD.n430 9.3005
R8412 VSSD.n428 VSSD.n177 9.3005
R8413 VSSD.n427 VSSD.n426 9.3005
R8414 VSSD.n425 VSSD.n179 9.3005
R8415 VSSD.n424 VSSD.n423 9.3005
R8416 VSSD.n421 VSSD.n180 9.3005
R8417 VSSD.n420 VSSD.n419 9.3005
R8418 VSSD.n418 VSSD.n182 9.3005
R8419 VSSD.n417 VSSD.n416 9.3005
R8420 VSSD.n415 VSSD.n183 9.3005
R8421 VSSD.n413 VSSD.n412 9.3005
R8422 VSSD.n411 VSSD.n185 9.3005
R8423 VSSD.n410 VSSD.n409 9.3005
R8424 VSSD.n408 VSSD.n186 9.3005
R8425 VSSD.n407 VSSD.n406 9.3005
R8426 VSSD.n405 VSSD.n187 9.3005
R8427 VSSD.n404 VSSD.n403 9.3005
R8428 VSSD.n401 VSSD.n188 9.3005
R8429 VSSD.n192 VSSD.n190 9.3005
R8430 VSSD.n399 VSSD.n398 9.3005
R8431 VSSD.n397 VSSD.n191 9.3005
R8432 VSSD.n396 VSSD.n395 9.3005
R8433 VSSD.n393 VSSD.n193 9.3005
R8434 VSSD.n392 VSSD.n391 9.3005
R8435 VSSD.n390 VSSD.n195 9.3005
R8436 VSSD.n389 VSSD.n388 9.3005
R8437 VSSD.n386 VSSD.n196 9.3005
R8438 VSSD.n385 VSSD.n384 9.3005
R8439 VSSD.n383 VSSD.n198 9.3005
R8440 VSSD.n382 VSSD.n381 9.3005
R8441 VSSD.n380 VSSD.n199 9.3005
R8442 VSSD.n378 VSSD.n377 9.3005
R8443 VSSD.n376 VSSD.n201 9.3005
R8444 VSSD.n375 VSSD.n374 9.3005
R8445 VSSD.n373 VSSD.n202 9.3005
R8446 VSSD.n372 VSSD.n371 9.3005
R8447 VSSD.n370 VSSD.n203 9.3005
R8448 VSSD.n369 VSSD.n368 9.3005
R8449 VSSD.n366 VSSD.n204 9.3005
R8450 VSSD.n211 VSSD.n206 9.3005
R8451 VSSD.n364 VSSD.n363 9.3005
R8452 VSSD.n362 VSSD.n210 9.3005
R8453 VSSD.n361 VSSD.n360 9.3005
R8454 VSSD.n358 VSSD.n212 9.3005
R8455 VSSD.n357 VSSD.n356 9.3005
R8456 VSSD.n355 VSSD.n214 9.3005
R8457 VSSD.n354 VSSD.n353 9.3005
R8458 VSSD.n351 VSSD.n215 9.3005
R8459 VSSD.n350 VSSD.n349 9.3005
R8460 VSSD.n348 VSSD.n217 9.3005
R8461 VSSD.n347 VSSD.n346 9.3005
R8462 VSSD.n345 VSSD.n218 9.3005
R8463 VSSD.n343 VSSD.n342 9.3005
R8464 VSSD.n341 VSSD.n220 9.3005
R8465 VSSD.n340 VSSD.n339 9.3005
R8466 VSSD.n338 VSSD.n221 9.3005
R8467 VSSD.n337 VSSD.n336 9.3005
R8468 VSSD.n335 VSSD.n222 9.3005
R8469 VSSD.n334 VSSD.n333 9.3005
R8470 VSSD.n331 VSSD.n223 9.3005
R8471 VSSD.n227 VSSD.n225 9.3005
R8472 VSSD.n329 VSSD.n328 9.3005
R8473 VSSD.n327 VSSD.n226 9.3005
R8474 VSSD.n326 VSSD.n325 9.3005
R8475 VSSD.n323 VSSD.n228 9.3005
R8476 VSSD.n322 VSSD.n321 9.3005
R8477 VSSD.n320 VSSD.n230 9.3005
R8478 VSSD.n319 VSSD.n318 9.3005
R8479 VSSD.n316 VSSD.n231 9.3005
R8480 VSSD.n315 VSSD.n314 9.3005
R8481 VSSD.n313 VSSD.n233 9.3005
R8482 VSSD.n312 VSSD.n311 9.3005
R8483 VSSD.n310 VSSD.n234 9.3005
R8484 VSSD.n308 VSSD.n307 9.3005
R8485 VSSD.n306 VSSD.n236 9.3005
R8486 VSSD.n305 VSSD.n304 9.3005
R8487 VSSD.n303 VSSD.n237 9.3005
R8488 VSSD.n302 VSSD.n301 9.3005
R8489 VSSD.n300 VSSD.n238 9.3005
R8490 VSSD.n299 VSSD.n298 9.3005
R8491 VSSD.n296 VSSD.n239 9.3005
R8492 VSSD.n243 VSSD.n241 9.3005
R8493 VSSD.n294 VSSD.n293 9.3005
R8494 VSSD.n656 VSSD.n655 9.3005
R8495 VSSD.n659 VSSD.n653 9.3005
R8496 VSSD.n662 VSSD.n661 9.3005
R8497 VSSD.n663 VSSD.n652 9.3005
R8498 VSSD.n665 VSSD.n664 9.3005
R8499 VSSD.n666 VSSD.n651 9.3005
R8500 VSSD.n668 VSSD.n667 9.3005
R8501 VSSD.n669 VSSD.n650 9.3005
R8502 VSSD.n671 VSSD.n670 9.3005
R8503 VSSD.n673 VSSD.n648 9.3005
R8504 VSSD.n675 VSSD.n674 9.3005
R8505 VSSD.n676 VSSD.n647 9.3005
R8506 VSSD.n678 VSSD.n677 9.3005
R8507 VSSD.n679 VSSD.n645 9.3005
R8508 VSSD.n682 VSSD.n681 9.3005
R8509 VSSD.n683 VSSD.n644 9.3005
R8510 VSSD.n685 VSSD.n684 9.3005
R8511 VSSD.n686 VSSD.n642 9.3005
R8512 VSSD.n689 VSSD.n688 9.3005
R8513 VSSD.n690 VSSD.n640 9.3005
R8514 VSSD.n498 VSSD.n497 9.3005
R8515 VSSD.n500 VSSD.n158 9.3005
R8516 VSSD.n502 VSSD.n501 9.3005
R8517 VSSD.n503 VSSD.n157 9.3005
R8518 VSSD.n505 VSSD.n504 9.3005
R8519 VSSD.n507 VSSD.n155 9.3005
R8520 VSSD.n509 VSSD.n508 9.3005
R8521 VSSD.n510 VSSD.n154 9.3005
R8522 VSSD.n512 VSSD.n511 9.3005
R8523 VSSD.n513 VSSD.n153 9.3005
R8524 VSSD.n517 VSSD.n516 9.3005
R8525 VSSD.n518 VSSD.n152 9.3005
R8526 VSSD.n520 VSSD.n519 9.3005
R8527 VSSD.n521 VSSD.n151 9.3005
R8528 VSSD.n523 VSSD.n522 9.3005
R8529 VSSD.n524 VSSD.n150 9.3005
R8530 VSSD.n526 VSSD.n525 9.3005
R8531 VSSD.n528 VSSD.n148 9.3005
R8532 VSSD.n531 VSSD.n530 9.3005
R8533 VSSD.n532 VSSD.n147 9.3005
R8534 VSSD.n534 VSSD.n533 9.3005
R8535 VSSD.n536 VSSD.n146 9.3005
R8536 VSSD.n539 VSSD.n538 9.3005
R8537 VSSD.n540 VSSD.n145 9.3005
R8538 VSSD.n542 VSSD.n541 9.3005
R8539 VSSD.n543 VSSD.n143 9.3005
R8540 VSSD.n546 VSSD.n545 9.3005
R8541 VSSD.n547 VSSD.n142 9.3005
R8542 VSSD.n549 VSSD.n548 9.3005
R8543 VSSD.n550 VSSD.n141 9.3005
R8544 VSSD.n554 VSSD.n553 9.3005
R8545 VSSD.n555 VSSD.n140 9.3005
R8546 VSSD.n557 VSSD.n556 9.3005
R8547 VSSD.n558 VSSD.n139 9.3005
R8548 VSSD.n560 VSSD.n559 9.3005
R8549 VSSD.n561 VSSD.n138 9.3005
R8550 VSSD.n563 VSSD.n562 9.3005
R8551 VSSD.n564 VSSD.n137 9.3005
R8552 VSSD.n567 VSSD.n566 9.3005
R8553 VSSD.n570 VSSD.n569 9.3005
R8554 VSSD.n572 VSSD.n571 9.3005
R8555 VSSD.n574 VSSD.n573 9.3005
R8556 VSSD.n576 VSSD.n575 9.3005
R8557 VSSD.n578 VSSD.n134 9.3005
R8558 VSSD.n580 VSSD.n579 9.3005
R8559 VSSD.n581 VSSD.n133 9.3005
R8560 VSSD.n583 VSSD.n582 9.3005
R8561 VSSD.n585 VSSD.n131 9.3005
R8562 VSSD.n587 VSSD.n586 9.3005
R8563 VSSD.n588 VSSD.n130 9.3005
R8564 VSSD.n590 VSSD.n589 9.3005
R8565 VSSD.n591 VSSD.n129 9.3005
R8566 VSSD.n595 VSSD.n594 9.3005
R8567 VSSD.n596 VSSD.n128 9.3005
R8568 VSSD.n598 VSSD.n597 9.3005
R8569 VSSD.n599 VSSD.n127 9.3005
R8570 VSSD.n601 VSSD.n600 9.3005
R8571 VSSD.n602 VSSD.n126 9.3005
R8572 VSSD.n604 VSSD.n603 9.3005
R8573 VSSD.n606 VSSD.n124 9.3005
R8574 VSSD.n609 VSSD.n608 9.3005
R8575 VSSD.n610 VSSD.n122 9.3005
R8576 VSSD.n761 VSSD.n760 9.3005
R8577 VSSD.n759 VSSD.n758 9.3005
R8578 VSSD.n756 VSSD.n611 9.3005
R8579 VSSD.n755 VSSD.n754 9.3005
R8580 VSSD.n753 VSSD.n612 9.3005
R8581 VSSD.n752 VSSD.n751 9.3005
R8582 VSSD.n749 VSSD.n613 9.3005
R8583 VSSD.n748 VSSD.n747 9.3005
R8584 VSSD.n746 VSSD.n615 9.3005
R8585 VSSD.n745 VSSD.n744 9.3005
R8586 VSSD.n743 VSSD.n616 9.3005
R8587 VSSD.n741 VSSD.n740 9.3005
R8588 VSSD.n739 VSSD.n618 9.3005
R8589 VSSD.n738 VSSD.n737 9.3005
R8590 VSSD.n736 VSSD.n619 9.3005
R8591 VSSD.n735 VSSD.n734 9.3005
R8592 VSSD.n733 VSSD.n620 9.3005
R8593 VSSD.n732 VSSD.n731 9.3005
R8594 VSSD.n729 VSSD.n621 9.3005
R8595 VSSD.n625 VSSD.n623 9.3005
R8596 VSSD.n727 VSSD.n726 9.3005
R8597 VSSD.n725 VSSD.n624 9.3005
R8598 VSSD.n724 VSSD.n723 9.3005
R8599 VSSD.n721 VSSD.n626 9.3005
R8600 VSSD.n720 VSSD.n719 9.3005
R8601 VSSD.n718 VSSD.n628 9.3005
R8602 VSSD.n717 VSSD.n716 9.3005
R8603 VSSD.n714 VSSD.n629 9.3005
R8604 VSSD.n713 VSSD.n712 9.3005
R8605 VSSD.n711 VSSD.n631 9.3005
R8606 VSSD.n710 VSSD.n709 9.3005
R8607 VSSD.n708 VSSD.n632 9.3005
R8608 VSSD.n706 VSSD.n705 9.3005
R8609 VSSD.n704 VSSD.n634 9.3005
R8610 VSSD.n703 VSSD.n702 9.3005
R8611 VSSD.n701 VSSD.n635 9.3005
R8612 VSSD.n700 VSSD.n699 9.3005
R8613 VSSD.n698 VSSD.n636 9.3005
R8614 VSSD.n697 VSSD.n696 9.3005
R8615 VSSD.n694 VSSD.n637 9.3005
R8616 VSSD.n641 VSSD.n639 9.3005
R8617 VSSD.n692 VSSD.n691 9.3005
R8618 VSSD.n493 VSSD.n492 9.3005
R8619 VSSD.n491 VSSD.n490 9.3005
R8620 VSSD.n489 VSSD.n488 9.3005
R8621 VSSD.n487 VSSD.n474 9.3005
R8622 VSSD.n485 VSSD.n484 9.3005
R8623 VSSD.n483 VSSD.n482 9.3005
R8624 VSSD.n481 VSSD.n478 9.3005
R8625 VSSD.n121 VSSD.n120 9.3005
R8626 VSSD.n769 VSSD.n768 9.3005
R8627 VSSD.n771 VSSD.n770 9.3005
R8628 VSSD.n773 VSSD.n772 9.3005
R8629 VSSD.n775 VSSD.n774 9.3005
R8630 VSSD.n776 VSSD.n116 9.3005
R8631 VSSD.n779 VSSD.n778 9.3005
R8632 VSSD.n780 VSSD.n115 9.3005
R8633 VSSD.n782 VSSD.n781 9.3005
R8634 VSSD.n784 VSSD.n114 9.3005
R8635 VSSD.n1627 VSSD.n1626 9.3005
R8636 VSSD.n1625 VSSD.n1385 9.3005
R8637 VSSD.n1624 VSSD.n1623 9.3005
R8638 VSSD.n1622 VSSD.n1386 9.3005
R8639 VSSD.n1621 VSSD.n1620 9.3005
R8640 VSSD.n1619 VSSD.n1389 9.3005
R8641 VSSD.n1618 VSSD.n1617 9.3005
R8642 VSSD.n1616 VSSD.n1390 9.3005
R8643 VSSD.n1615 VSSD.n1614 9.3005
R8644 VSSD.n1613 VSSD.n1391 9.3005
R8645 VSSD.n1612 VSSD.n1611 9.3005
R8646 VSSD.n1610 VSSD.n1392 9.3005
R8647 VSSD.n1609 VSSD.n1608 9.3005
R8648 VSSD.n1607 VSSD.n1395 9.3005
R8649 VSSD.n1606 VSSD.n1605 9.3005
R8650 VSSD.n1602 VSSD.n1396 9.3005
R8651 VSSD.n1601 VSSD.n1600 9.3005
R8652 VSSD.n1599 VSSD.n1397 9.3005
R8653 VSSD.n1598 VSSD.n1597 9.3005
R8654 VSSD.n1596 VSSD.n1398 9.3005
R8655 VSSD.n1595 VSSD.n1594 9.3005
R8656 VSSD.n1593 VSSD.n1399 9.3005
R8657 VSSD.n1592 VSSD.n1591 9.3005
R8658 VSSD.n1590 VSSD.n1400 9.3005
R8659 VSSD.n1588 VSSD.n1587 9.3005
R8660 VSSD.n1586 VSSD.n1401 9.3005
R8661 VSSD.n1585 VSSD.n1584 9.3005
R8662 VSSD.n1583 VSSD.n1402 9.3005
R8663 VSSD.n1582 VSSD.n1581 9.3005
R8664 VSSD.n1580 VSSD.n1403 9.3005
R8665 VSSD.n1579 VSSD.n1578 9.3005
R8666 VSSD.n1575 VSSD.n1404 9.3005
R8667 VSSD.n1574 VSSD.n1573 9.3005
R8668 VSSD.n1572 VSSD.n1405 9.3005
R8669 VSSD.n1571 VSSD.n1570 9.3005
R8670 VSSD.n1569 VSSD.n1406 9.3005
R8671 VSSD.n1566 VSSD.n1565 9.3005
R8672 VSSD.n1564 VSSD.n1407 9.3005
R8673 VSSD.n1563 VSSD.n1562 9.3005
R8674 VSSD.n1561 VSSD.n1408 9.3005
R8675 VSSD.n1560 VSSD.n1559 9.3005
R8676 VSSD.n1558 VSSD.n1409 9.3005
R8677 VSSD.n1557 VSSD.n1556 9.3005
R8678 VSSD.n1555 VSSD.n1410 9.3005
R8679 VSSD.n1554 VSSD.n1552 9.3005
R8680 VSSD.n1551 VSSD.n1411 9.3005
R8681 VSSD.n1550 VSSD.n1549 9.3005
R8682 VSSD.n1548 VSSD.n1412 9.3005
R8683 VSSD.n1547 VSSD.n1546 9.3005
R8684 VSSD.n1545 VSSD.n1413 9.3005
R8685 VSSD.n1544 VSSD.n1543 9.3005
R8686 VSSD.n1542 VSSD.n1414 9.3005
R8687 VSSD.n1539 VSSD.n1538 9.3005
R8688 VSSD.n1537 VSSD.n1415 9.3005
R8689 VSSD.n1536 VSSD.n1535 9.3005
R8690 VSSD.n1534 VSSD.n1416 9.3005
R8691 VSSD.n1533 VSSD.n1532 9.3005
R8692 VSSD.n1531 VSSD.n1530 9.3005
R8693 VSSD.n1529 VSSD.n1419 9.3005
R8694 VSSD.n1528 VSSD.n1527 9.3005
R8695 VSSD.n1526 VSSD.n1420 9.3005
R8696 VSSD.n1525 VSSD.n1524 9.3005
R8697 VSSD.n1523 VSSD.n1421 9.3005
R8698 VSSD.n1522 VSSD.n1521 9.3005
R8699 VSSD.n1520 VSSD.n1422 9.3005
R8700 VSSD.n1519 VSSD.n1518 9.3005
R8701 VSSD.n1516 VSSD.n1423 9.3005
R8702 VSSD.n1515 VSSD.n1514 9.3005
R8703 VSSD.n1513 VSSD.n1424 9.3005
R8704 VSSD.n1512 VSSD.n1511 9.3005
R8705 VSSD.n1510 VSSD.n1425 9.3005
R8706 VSSD.n1509 VSSD.n1508 9.3005
R8707 VSSD.n1507 VSSD.n1426 9.3005
R8708 VSSD.n1506 VSSD.n1505 9.3005
R8709 VSSD.n1504 VSSD.n1427 9.3005
R8710 VSSD.n1503 VSSD.n1502 9.3005
R8711 VSSD.n1501 VSSD.n1430 9.3005
R8712 VSSD.n1500 VSSD.n1499 9.3005
R8713 VSSD.n1496 VSSD.n1431 9.3005
R8714 VSSD.n1495 VSSD.n1494 9.3005
R8715 VSSD.n1493 VSSD.n1432 9.3005
R8716 VSSD.n1492 VSSD.n1491 9.3005
R8717 VSSD.n1490 VSSD.n1433 9.3005
R8718 VSSD.n1489 VSSD.n1488 9.3005
R8719 VSSD.n1487 VSSD.n1434 9.3005
R8720 VSSD.n1486 VSSD.n1485 9.3005
R8721 VSSD.n1484 VSSD.n1435 9.3005
R8722 VSSD.n1482 VSSD.n1481 9.3005
R8723 VSSD.n1480 VSSD.n1436 9.3005
R8724 VSSD.n1479 VSSD.n1478 9.3005
R8725 VSSD.n1477 VSSD.n1437 9.3005
R8726 VSSD.n1476 VSSD.n1475 9.3005
R8727 VSSD.n1474 VSSD.n1438 9.3005
R8728 VSSD.n1473 VSSD.n1472 9.3005
R8729 VSSD.n1469 VSSD.n1439 9.3005
R8730 VSSD.n1468 VSSD.n1467 9.3005
R8731 VSSD.n1466 VSSD.n1440 9.3005
R8732 VSSD.n1465 VSSD.n1464 9.3005
R8733 VSSD.n1463 VSSD.n1441 9.3005
R8734 VSSD.n1460 VSSD.n1459 9.3005
R8735 VSSD.n1458 VSSD.n1442 9.3005
R8736 VSSD.n1457 VSSD.n1456 9.3005
R8737 VSSD.n1455 VSSD.n1443 9.3005
R8738 VSSD.n1454 VSSD.n1453 9.3005
R8739 VSSD.n1452 VSSD.n1444 9.3005
R8740 VSSD.n1451 VSSD.n1450 9.3005
R8741 VSSD.n1449 VSSD.n1445 9.3005
R8742 VSSD.n1818 VSSD.n1817 9.3005
R8743 VSSD.n1634 VSSD.n1633 9.3005
R8744 VSSD.n1635 VSSD.n1384 9.3005
R8745 VSSD.n1639 VSSD.n1638 9.3005
R8746 VSSD.n1640 VSSD.n1383 9.3005
R8747 VSSD.n1642 VSSD.n1641 9.3005
R8748 VSSD.n1645 VSSD.n1644 9.3005
R8749 VSSD.n1646 VSSD.n1382 9.3005
R8750 VSSD.n1648 VSSD.n1647 9.3005
R8751 VSSD.n1649 VSSD.n1381 9.3005
R8752 VSSD.n1651 VSSD.n1650 9.3005
R8753 VSSD.n1652 VSSD.n1380 9.3005
R8754 VSSD.n1654 VSSD.n1653 9.3005
R8755 VSSD.n1655 VSSD.n1379 9.3005
R8756 VSSD.n1657 VSSD.n1656 9.3005
R8757 VSSD.n1659 VSSD.n1658 9.3005
R8758 VSSD.n1660 VSSD.n1376 9.3005
R8759 VSSD.n1662 VSSD.n1661 9.3005
R8760 VSSD.n1663 VSSD.n1375 9.3005
R8761 VSSD.n1665 VSSD.n1664 9.3005
R8762 VSSD.n1668 VSSD.n1374 9.3005
R8763 VSSD.n1670 VSSD.n1669 9.3005
R8764 VSSD.n1671 VSSD.n1373 9.3005
R8765 VSSD.n1673 VSSD.n1672 9.3005
R8766 VSSD.n1674 VSSD.n1372 9.3005
R8767 VSSD.n1676 VSSD.n1675 9.3005
R8768 VSSD.n1677 VSSD.n1370 9.3005
R8769 VSSD.n1679 VSSD.n1678 9.3005
R8770 VSSD.n1680 VSSD.n1369 9.3005
R8771 VSSD.n1682 VSSD.n1681 9.3005
R8772 VSSD.n1683 VSSD.n1368 9.3005
R8773 VSSD.n1685 VSSD.n1684 9.3005
R8774 VSSD.n1686 VSSD.n1367 9.3005
R8775 VSSD.n1688 VSSD.n1687 9.3005
R8776 VSSD.n1689 VSSD.n1366 9.3005
R8777 VSSD.n1691 VSSD.n1690 9.3005
R8778 VSSD.n1694 VSSD.n1365 9.3005
R8779 VSSD.n1696 VSSD.n1695 9.3005
R8780 VSSD.n1697 VSSD.n1364 9.3005
R8781 VSSD.n1699 VSSD.n1698 9.3005
R8782 VSSD.n1700 VSSD.n1363 9.3005
R8783 VSSD.n1704 VSSD.n1703 9.3005
R8784 VSSD.n1705 VSSD.n1362 9.3005
R8785 VSSD.n1707 VSSD.n1706 9.3005
R8786 VSSD.n1708 VSSD.n1361 9.3005
R8787 VSSD.n1710 VSSD.n1709 9.3005
R8788 VSSD.n1711 VSSD.n1360 9.3005
R8789 VSSD.n1713 VSSD.n1712 9.3005
R8790 VSSD.n1716 VSSD.n1715 9.3005
R8791 VSSD.n1717 VSSD.n1359 9.3005
R8792 VSSD.n1719 VSSD.n1718 9.3005
R8793 VSSD.n1720 VSSD.n1358 9.3005
R8794 VSSD.n1722 VSSD.n1721 9.3005
R8795 VSSD.n1723 VSSD.n1357 9.3005
R8796 VSSD.n1725 VSSD.n1724 9.3005
R8797 VSSD.n1726 VSSD.n1356 9.3005
R8798 VSSD.n1728 VSSD.n1727 9.3005
R8799 VSSD.n1730 VSSD.n1729 9.3005
R8800 VSSD.n1731 VSSD.n1353 9.3005
R8801 VSSD.n1733 VSSD.n1732 9.3005
R8802 VSSD.n1734 VSSD.n1352 9.3005
R8803 VSSD.n1736 VSSD.n1735 9.3005
R8804 VSSD.n1739 VSSD.n1351 9.3005
R8805 VSSD.n1741 VSSD.n1740 9.3005
R8806 VSSD.n1742 VSSD.n1350 9.3005
R8807 VSSD.n1744 VSSD.n1743 9.3005
R8808 VSSD.n1745 VSSD.n1349 9.3005
R8809 VSSD.n1747 VSSD.n1746 9.3005
R8810 VSSD.n1748 VSSD.n1347 9.3005
R8811 VSSD.n1750 VSSD.n1749 9.3005
R8812 VSSD.n1751 VSSD.n1346 9.3005
R8813 VSSD.n1753 VSSD.n1752 9.3005
R8814 VSSD.n1754 VSSD.n1345 9.3005
R8815 VSSD.n1756 VSSD.n1755 9.3005
R8816 VSSD.n1757 VSSD.n1344 9.3005
R8817 VSSD.n1759 VSSD.n1758 9.3005
R8818 VSSD.n1760 VSSD.n1343 9.3005
R8819 VSSD.n1762 VSSD.n1761 9.3005
R8820 VSSD.n1765 VSSD.n1342 9.3005
R8821 VSSD.n1767 VSSD.n1766 9.3005
R8822 VSSD.n1768 VSSD.n1341 9.3005
R8823 VSSD.n1770 VSSD.n1769 9.3005
R8824 VSSD.n1771 VSSD.n1340 9.3005
R8825 VSSD.n1775 VSSD.n1774 9.3005
R8826 VSSD.n1776 VSSD.n1339 9.3005
R8827 VSSD.n1778 VSSD.n1777 9.3005
R8828 VSSD.n1779 VSSD.n1338 9.3005
R8829 VSSD.n1781 VSSD.n1780 9.3005
R8830 VSSD.n1782 VSSD.n1337 9.3005
R8831 VSSD.n1784 VSSD.n1783 9.3005
R8832 VSSD.n1787 VSSD.n1786 9.3005
R8833 VSSD.n1788 VSSD.n1336 9.3005
R8834 VSSD.n1790 VSSD.n1789 9.3005
R8835 VSSD.n1791 VSSD.n1335 9.3005
R8836 VSSD.n1793 VSSD.n1792 9.3005
R8837 VSSD.n1794 VSSD.n1334 9.3005
R8838 VSSD.n1796 VSSD.n1795 9.3005
R8839 VSSD.n1797 VSSD.n1333 9.3005
R8840 VSSD.n1799 VSSD.n1798 9.3005
R8841 VSSD.n1801 VSSD.n1800 9.3005
R8842 VSSD.n1802 VSSD.n1330 9.3005
R8843 VSSD.n1804 VSSD.n1803 9.3005
R8844 VSSD.n1805 VSSD.n1329 9.3005
R8845 VSSD.n1807 VSSD.n1806 9.3005
R8846 VSSD.n1810 VSSD.n1328 9.3005
R8847 VSSD.n1812 VSSD.n1811 9.3005
R8848 VSSD.n1813 VSSD.n1327 9.3005
R8849 VSSD.n1815 VSSD.n1814 9.3005
R8850 VSSD.n1816 VSSD.n1326 9.3005
R8851 VSSD.n959 VSSD.n955 9.3005
R8852 VSSD.n961 VSSD.n960 9.3005
R8853 VSSD.n962 VSSD.n952 9.3005
R8854 VSSD.n965 VSSD.n964 9.3005
R8855 VSSD.n966 VSSD.n951 9.3005
R8856 VSSD.n968 VSSD.n967 9.3005
R8857 VSSD.n969 VSSD.n950 9.3005
R8858 VSSD.n974 VSSD.n973 9.3005
R8859 VSSD.n975 VSSD.n949 9.3005
R8860 VSSD.n977 VSSD.n976 9.3005
R8861 VSSD.n978 VSSD.n948 9.3005
R8862 VSSD.n980 VSSD.n979 9.3005
R8863 VSSD.n981 VSSD.n947 9.3005
R8864 VSSD.n983 VSSD.n982 9.3005
R8865 VSSD.n984 VSSD.n946 9.3005
R8866 VSSD.n986 VSSD.n985 9.3005
R8867 VSSD.n987 VSSD.n945 9.3005
R8868 VSSD.n989 VSSD.n988 9.3005
R8869 VSSD.n990 VSSD.n942 9.3005
R8870 VSSD.n991 VSSD.n941 9.3005
R8871 VSSD.n993 VSSD.n992 9.3005
R8872 VSSD.n994 VSSD.n940 9.3005
R8873 VSSD.n996 VSSD.n995 9.3005
R8874 VSSD.n997 VSSD.n937 9.3005
R8875 VSSD.n1000 VSSD.n999 9.3005
R8876 VSSD.n1001 VSSD.n936 9.3005
R8877 VSSD.n1003 VSSD.n1002 9.3005
R8878 VSSD.n1004 VSSD.n935 9.3005
R8879 VSSD.n1009 VSSD.n1008 9.3005
R8880 VSSD.n1010 VSSD.n934 9.3005
R8881 VSSD.n1012 VSSD.n1011 9.3005
R8882 VSSD.n1013 VSSD.n933 9.3005
R8883 VSSD.n1015 VSSD.n1014 9.3005
R8884 VSSD.n1016 VSSD.n932 9.3005
R8885 VSSD.n1018 VSSD.n1017 9.3005
R8886 VSSD.n1019 VSSD.n931 9.3005
R8887 VSSD.n1021 VSSD.n1020 9.3005
R8888 VSSD.n1022 VSSD.n930 9.3005
R8889 VSSD.n1024 VSSD.n1023 9.3005
R8890 VSSD.n1025 VSSD.n927 9.3005
R8891 VSSD.n1026 VSSD.n926 9.3005
R8892 VSSD.n1028 VSSD.n1027 9.3005
R8893 VSSD.n1029 VSSD.n925 9.3005
R8894 VSSD.n1031 VSSD.n1030 9.3005
R8895 VSSD.n1032 VSSD.n922 9.3005
R8896 VSSD.n1035 VSSD.n1034 9.3005
R8897 VSSD.n1036 VSSD.n921 9.3005
R8898 VSSD.n1038 VSSD.n1037 9.3005
R8899 VSSD.n1039 VSSD.n920 9.3005
R8900 VSSD.n1044 VSSD.n1043 9.3005
R8901 VSSD.n1045 VSSD.n919 9.3005
R8902 VSSD.n1047 VSSD.n1046 9.3005
R8903 VSSD.n1048 VSSD.n918 9.3005
R8904 VSSD.n1050 VSSD.n1049 9.3005
R8905 VSSD.n1051 VSSD.n917 9.3005
R8906 VSSD.n1053 VSSD.n1052 9.3005
R8907 VSSD.n1054 VSSD.n916 9.3005
R8908 VSSD.n1056 VSSD.n1055 9.3005
R8909 VSSD.n1057 VSSD.n915 9.3005
R8910 VSSD.n1059 VSSD.n1058 9.3005
R8911 VSSD.n1060 VSSD.n912 9.3005
R8912 VSSD.n1061 VSSD.n911 9.3005
R8913 VSSD.n1063 VSSD.n1062 9.3005
R8914 VSSD.n1064 VSSD.n910 9.3005
R8915 VSSD.n1066 VSSD.n1065 9.3005
R8916 VSSD.n1067 VSSD.n907 9.3005
R8917 VSSD.n1070 VSSD.n1069 9.3005
R8918 VSSD.n1071 VSSD.n906 9.3005
R8919 VSSD.n1073 VSSD.n1072 9.3005
R8920 VSSD.n1074 VSSD.n905 9.3005
R8921 VSSD.n1079 VSSD.n1078 9.3005
R8922 VSSD.n1080 VSSD.n904 9.3005
R8923 VSSD.n1082 VSSD.n1081 9.3005
R8924 VSSD.n1083 VSSD.n903 9.3005
R8925 VSSD.n1085 VSSD.n1084 9.3005
R8926 VSSD.n1086 VSSD.n902 9.3005
R8927 VSSD.n1088 VSSD.n1087 9.3005
R8928 VSSD.n1089 VSSD.n901 9.3005
R8929 VSSD.n1091 VSSD.n1090 9.3005
R8930 VSSD.n1092 VSSD.n900 9.3005
R8931 VSSD.n1094 VSSD.n1093 9.3005
R8932 VSSD.n1095 VSSD.n897 9.3005
R8933 VSSD.n1096 VSSD.n896 9.3005
R8934 VSSD.n1098 VSSD.n1097 9.3005
R8935 VSSD.n1099 VSSD.n895 9.3005
R8936 VSSD.n1101 VSSD.n1100 9.3005
R8937 VSSD.n1102 VSSD.n892 9.3005
R8938 VSSD.n1105 VSSD.n1104 9.3005
R8939 VSSD.n1106 VSSD.n891 9.3005
R8940 VSSD.n1108 VSSD.n1107 9.3005
R8941 VSSD.n1109 VSSD.n890 9.3005
R8942 VSSD.n1114 VSSD.n1113 9.3005
R8943 VSSD.n1115 VSSD.n889 9.3005
R8944 VSSD.n1117 VSSD.n1116 9.3005
R8945 VSSD.n1118 VSSD.n888 9.3005
R8946 VSSD.n1120 VSSD.n1119 9.3005
R8947 VSSD.n1121 VSSD.n887 9.3005
R8948 VSSD.n1123 VSSD.n1122 9.3005
R8949 VSSD.n1124 VSSD.n886 9.3005
R8950 VSSD.n1126 VSSD.n1125 9.3005
R8951 VSSD.n1127 VSSD.n885 9.3005
R8952 VSSD.n1129 VSSD.n1128 9.3005
R8953 VSSD.n1130 VSSD.n882 9.3005
R8954 VSSD.n1131 VSSD.n881 9.3005
R8955 VSSD.n1133 VSSD.n1132 9.3005
R8956 VSSD.n1134 VSSD.n880 9.3005
R8957 VSSD.n1136 VSSD.n1135 9.3005
R8958 VSSD.n1137 VSSD.n877 9.3005
R8959 VSSD.n1140 VSSD.n1139 9.3005
R8960 VSSD.n1141 VSSD.n876 9.3005
R8961 VSSD.n1143 VSSD.n1142 9.3005
R8962 VSSD.n1144 VSSD.n875 9.3005
R8963 VSSD.n1149 VSSD.n1148 9.3005
R8964 VSSD.n1150 VSSD.n874 9.3005
R8965 VSSD.n1152 VSSD.n1151 9.3005
R8966 VSSD.n1153 VSSD.n873 9.3005
R8967 VSSD.n1155 VSSD.n1154 9.3005
R8968 VSSD.n1156 VSSD.n872 9.3005
R8969 VSSD.n1158 VSSD.n1157 9.3005
R8970 VSSD.n1159 VSSD.n871 9.3005
R8971 VSSD.n1161 VSSD.n1160 9.3005
R8972 VSSD.n1162 VSSD.n870 9.3005
R8973 VSSD.n1164 VSSD.n1163 9.3005
R8974 VSSD.n1165 VSSD.n867 9.3005
R8975 VSSD.n1166 VSSD.n866 9.3005
R8976 VSSD.n1168 VSSD.n1167 9.3005
R8977 VSSD.n1169 VSSD.n865 9.3005
R8978 VSSD.n1171 VSSD.n1170 9.3005
R8979 VSSD.n1172 VSSD.n862 9.3005
R8980 VSSD.n1175 VSSD.n1174 9.3005
R8981 VSSD.n1176 VSSD.n861 9.3005
R8982 VSSD.n1178 VSSD.n1177 9.3005
R8983 VSSD.n1179 VSSD.n860 9.3005
R8984 VSSD.n1184 VSSD.n1183 9.3005
R8985 VSSD.n1185 VSSD.n859 9.3005
R8986 VSSD.n1187 VSSD.n1186 9.3005
R8987 VSSD.n1188 VSSD.n858 9.3005
R8988 VSSD.n1190 VSSD.n1189 9.3005
R8989 VSSD.n1191 VSSD.n857 9.3005
R8990 VSSD.n1193 VSSD.n1192 9.3005
R8991 VSSD.n1194 VSSD.n856 9.3005
R8992 VSSD.n1196 VSSD.n1195 9.3005
R8993 VSSD.n1197 VSSD.n855 9.3005
R8994 VSSD.n1199 VSSD.n1198 9.3005
R8995 VSSD.n1200 VSSD.n852 9.3005
R8996 VSSD.n1201 VSSD.n851 9.3005
R8997 VSSD.n1203 VSSD.n1202 9.3005
R8998 VSSD.n1204 VSSD.n850 9.3005
R8999 VSSD.n1206 VSSD.n1205 9.3005
R9000 VSSD.n1207 VSSD.n847 9.3005
R9001 VSSD.n1210 VSSD.n1209 9.3005
R9002 VSSD.n1211 VSSD.n846 9.3005
R9003 VSSD.n1213 VSSD.n1212 9.3005
R9004 VSSD.n1214 VSSD.n845 9.3005
R9005 VSSD.n1219 VSSD.n1218 9.3005
R9006 VSSD.n1220 VSSD.n844 9.3005
R9007 VSSD.n1222 VSSD.n1221 9.3005
R9008 VSSD.n1223 VSSD.n843 9.3005
R9009 VSSD.n1225 VSSD.n1224 9.3005
R9010 VSSD.n1226 VSSD.n842 9.3005
R9011 VSSD.n1228 VSSD.n1227 9.3005
R9012 VSSD.n1229 VSSD.n841 9.3005
R9013 VSSD.n1231 VSSD.n1230 9.3005
R9014 VSSD.n1232 VSSD.n840 9.3005
R9015 VSSD.n1234 VSSD.n1233 9.3005
R9016 VSSD.n1235 VSSD.n837 9.3005
R9017 VSSD.n1236 VSSD.n836 9.3005
R9018 VSSD.n1238 VSSD.n1237 9.3005
R9019 VSSD.n1239 VSSD.n835 9.3005
R9020 VSSD.n1241 VSSD.n1240 9.3005
R9021 VSSD.n1242 VSSD.n832 9.3005
R9022 VSSD.n1245 VSSD.n1244 9.3005
R9023 VSSD.n1246 VSSD.n831 9.3005
R9024 VSSD.n1248 VSSD.n1247 9.3005
R9025 VSSD.n1249 VSSD.n830 9.3005
R9026 VSSD.n1254 VSSD.n1253 9.3005
R9027 VSSD.n1255 VSSD.n829 9.3005
R9028 VSSD.n1257 VSSD.n1256 9.3005
R9029 VSSD.n1258 VSSD.n828 9.3005
R9030 VSSD.n1260 VSSD.n1259 9.3005
R9031 VSSD.n1261 VSSD.n827 9.3005
R9032 VSSD.n1263 VSSD.n1262 9.3005
R9033 VSSD.n1264 VSSD.n826 9.3005
R9034 VSSD.n1266 VSSD.n1265 9.3005
R9035 VSSD.n1267 VSSD.n825 9.3005
R9036 VSSD.n1269 VSSD.n1268 9.3005
R9037 VSSD.n1270 VSSD.n822 9.3005
R9038 VSSD.n1271 VSSD.n821 9.3005
R9039 VSSD.n1273 VSSD.n1272 9.3005
R9040 VSSD.n1274 VSSD.n820 9.3005
R9041 VSSD.n1276 VSSD.n1275 9.3005
R9042 VSSD.n1277 VSSD.n817 9.3005
R9043 VSSD.n1280 VSSD.n1279 9.3005
R9044 VSSD.n1281 VSSD.n816 9.3005
R9045 VSSD.n1283 VSSD.n1282 9.3005
R9046 VSSD.n1284 VSSD.n815 9.3005
R9047 VSSD.n1289 VSSD.n1288 9.3005
R9048 VSSD.n1290 VSSD.n814 9.3005
R9049 VSSD.n1292 VSSD.n1291 9.3005
R9050 VSSD.n1293 VSSD.n813 9.3005
R9051 VSSD.n1295 VSSD.n1294 9.3005
R9052 VSSD.n1296 VSSD.n812 9.3005
R9053 VSSD.n1298 VSSD.n1297 9.3005
R9054 VSSD.n1299 VSSD.n811 9.3005
R9055 VSSD.n1300 VSSD.n808 9.3005
R9056 VSSD.n1302 VSSD.n1301 9.3005
R9057 VSSD.n1303 VSSD.n807 9.3005
R9058 VSSD.n1305 VSSD.n1304 9.3005
R9059 VSSD.n1306 VSSD.n806 9.3005
R9060 VSSD.n1308 VSSD.n1307 9.3005
R9061 VSSD.n1309 VSSD.n805 9.3005
R9062 VSSD.n1311 VSSD.n1310 9.3005
R9063 VSSD.n1313 VSSD.n800 9.3005
R9064 VSSD.n1315 VSSD.n1314 9.3005
R9065 VSSD.n1317 VSSD.n1316 9.3005
R9066 VSSD.n1318 VSSD.n795 9.3005
R9067 VSSD.n1319 VSSD.n791 9.3005
R9068 VSSD.n1321 VSSD.n1320 9.3005
R9069 VSSD.n1322 VSSD.n0 9.3005
R9070 VSSD.n762 VSSD.n122 9.05896
R9071 VSSD.n762 VSSD.n761 9.05896
R9072 VSSD.n789 VSSD.n788 8.65442
R9073 VSSD.n1820 VSSD.n1325 8.56446
R9074 VSSD.n1822 VSSD.n1325 8.338
R9075 VSSD.n1324 VSSD.n112 8.338
R9076 VSSD.t1162 VSSD 8.24792
R9077 VSSD.n790 VSSD.n789 8.133
R9078 VSSD.n469 VSSD.n160 8.07435
R9079 VSSD.n492 VSSD.n472 8.07435
R9080 VSSD.n1656 VSSD.n1378 7.90638
R9081 VSSD.n1693 VSSD.n1691 7.90638
R9082 VSSD.n1727 VSSD.n1355 7.90638
R9083 VSSD.n1764 VSSD.n1762 7.90638
R9084 VSSD.n1798 VSSD.n1332 7.90638
R9085 VSSD.n1462 VSSD.n1460 7.90638
R9086 VSSD.n1498 VSSD.n1496 7.90638
R9087 VSSD.n1530 VSSD.n1418 7.90638
R9088 VSSD.n1568 VSSD.n1566 7.90638
R9089 VSSD.n1604 VSSD.n1602 7.90638
R9090 VSSD.n1869 VSSD.n1867 7.90638
R9091 VSSD.n97 VSSD.n94 7.90638
R9092 VSSD.n15 VSSD.n12 7.90638
R9093 VSSD.n1995 VSSD.n1994 7.90638
R9094 VSSD.n36 VSSD.n33 7.90638
R9095 VSSD.n1964 VSSD.n1963 7.90638
R9096 VSSD.n57 VSSD.n54 7.90638
R9097 VSSD.n1933 VSSD.n1932 7.90638
R9098 VSSD.n78 VSSD.n75 7.90638
R9099 VSSD.n1902 VSSD.n1901 7.90638
R9100 VSSD.n1287 VSSD.n814 7.90638
R9101 VSSD.n1252 VSSD.n829 7.90638
R9102 VSSD.n1217 VSSD.n844 7.90638
R9103 VSSD.n1182 VSSD.n859 7.90638
R9104 VSSD.n1147 VSSD.n874 7.90638
R9105 VSSD.n1112 VSSD.n889 7.90638
R9106 VSSD.n1077 VSSD.n904 7.90638
R9107 VSSD.n1042 VSSD.n919 7.90638
R9108 VSSD.n1007 VSSD.n934 7.90638
R9109 VSSD.n972 VSSD.n949 7.90638
R9110 VSSD.n437 VSSD.n171 7.6805
R9111 VSSD.n402 VSSD.n187 7.6805
R9112 VSSD.n367 VSSD.n203 7.6805
R9113 VSSD.n332 VSSD.n222 7.6805
R9114 VSSD.n297 VSSD.n238 7.6805
R9115 VSSD.n262 VSSD.n254 7.6805
R9116 VSSD.n527 VSSD.n150 7.6805
R9117 VSSD.n565 VSSD.n563 7.6805
R9118 VSSD.n605 VSSD.n126 7.6805
R9119 VSSD.n730 VSSD.n620 7.6805
R9120 VSSD.n695 VSSD.n636 7.6805
R9121 VSSD.n660 VSSD.n652 7.6805
R9122 VSSD.n1448 VSSD.n1446 7.12063
R9123 VSSD.n1830 VSSD.n1829 6.94395
R9124 VSSD.n763 VSSD.n762 6.88285
R9125 VSSD.n958 VSSD.n956 6.74107
R9126 VSSD.n958 VSSD.n957 6.48892
R9127 VSSD.n1637 VSSD.n1635 6.4005
R9128 VSSD.n1388 VSSD.n1385 6.4005
R9129 VSSD.n1837 VSSD.n1835 6.4005
R9130 VSSD.n1312 VSSD.n1311 6.4005
R9131 VSSD.t1164 VSSD.t857 6.18607
R9132 VSSD.n768 VSSD.n767 6.10512
R9133 VSSD.n771 VSSD.n119 5.90819
R9134 VSSD.n457 VSSD.n456 5.1205
R9135 VSSD.n422 VSSD.n421 5.1205
R9136 VSSD.n387 VSSD.n386 5.1205
R9137 VSSD.n352 VSSD.n351 5.1205
R9138 VSSD.n317 VSSD.n316 5.1205
R9139 VSSD.n282 VSSD.n281 5.1205
R9140 VSSD.n507 VSSD.n506 5.1205
R9141 VSSD.n545 VSSD.n544 5.1205
R9142 VSSD.n585 VSSD.n584 5.1205
R9143 VSSD.n750 VSSD.n749 5.1205
R9144 VSSD.n715 VSSD.n714 5.1205
R9145 VSSD.n680 VSSD.n679 5.1205
R9146 VSSD.n1821 VSSD.n1820 5.02915
R9147 VSSD.n788 VSSD.n110 5.02264
R9148 VSSD.n1824 VSSD.n113 5.02264
R9149 VSSD.n480 VSSD.n121 4.52973
R9150 VSSD.n1824 VSSD.n1823 4.5005
R9151 VSSD.n790 VSSD.n110 4.5005
R9152 VSSD.n1822 VSSD.n1821 4.5005
R9153 VSSD.n1819 VSSD.n112 4.5005
R9154 VSSD.n1826 VSSD.n1825 4.5005
R9155 VSSD.n1828 VSSD.n1827 4.5005
R9156 VSSD.n787 VSSD.n111 4.5005
R9157 VSSD.n1823 VSSD.n790 4.38425
R9158 VSSD.n1827 VSSD.n1826 4.38425
R9159 VSSD.n788 VSSD.n113 4.38353
R9160 VSSD.n449 VSSD.n448 4.13588
R9161 VSSD.n414 VSSD.n413 4.13588
R9162 VSSD.n379 VSSD.n378 4.13588
R9163 VSSD.n344 VSSD.n343 4.13588
R9164 VSSD.n309 VSSD.n308 4.13588
R9165 VSSD.n274 VSSD.n273 4.13588
R9166 VSSD.n516 VSSD.n515 4.13588
R9167 VSSD.n552 VSSD.n140 4.13588
R9168 VSSD.n594 VSSD.n593 4.13588
R9169 VSSD.n742 VSSD.n741 4.13588
R9170 VSSD.n707 VSSD.n706 4.13588
R9171 VSSD.n672 VSSD.n671 4.13588
R9172 VSSD.n1827 VSSD.n111 3.633
R9173 VSSD.n1838 VSSD.n1837 3.38874
R9174 VSSD.n1313 VSSD.n1312 3.38874
R9175 VSSD.n111 VSSD 3.2355
R9176 VSSD.n438 VSSD.n437 3.10353
R9177 VSSD.n435 VSSD.n174 3.10353
R9178 VSSD.n403 VSSD.n402 3.10353
R9179 VSSD.n400 VSSD.n190 3.10353
R9180 VSSD.n368 VSSD.n367 3.10353
R9181 VSSD.n365 VSSD.n206 3.10353
R9182 VSSD.n333 VSSD.n332 3.10353
R9183 VSSD.n330 VSSD.n225 3.10353
R9184 VSSD.n298 VSSD.n297 3.10353
R9185 VSSD.n295 VSSD.n241 3.10353
R9186 VSSD.n263 VSSD.n262 3.10353
R9187 VSSD.n260 VSSD.n257 3.10353
R9188 VSSD.n527 VSSD.n526 3.10353
R9189 VSSD.n530 VSSD.n529 3.10353
R9190 VSSD.n565 VSSD.n564 3.10353
R9191 VSSD.n569 VSSD.n136 3.10353
R9192 VSSD.n605 VSSD.n604 3.10353
R9193 VSSD.n608 VSSD.n607 3.10353
R9194 VSSD.n731 VSSD.n730 3.10353
R9195 VSSD.n728 VSSD.n623 3.10353
R9196 VSSD.n696 VSSD.n695 3.10353
R9197 VSSD.n693 VSSD.n639 3.10353
R9198 VSSD.n661 VSSD.n660 3.10353
R9199 VSSD.n658 VSSD.n655 3.10353
R9200 VSSD.n1667 VSSD.n1665 2.63579
R9201 VSSD.n1702 VSSD.n1700 2.63579
R9202 VSSD.n1738 VSSD.n1736 2.63579
R9203 VSSD.n1773 VSSD.n1771 2.63579
R9204 VSSD.n1809 VSSD.n1807 2.63579
R9205 VSSD.n1471 VSSD.n1469 2.63579
R9206 VSSD.n1505 VSSD.n1429 2.63579
R9207 VSSD.n1541 VSSD.n1539 2.63579
R9208 VSSD.n1577 VSSD.n1575 2.63579
R9209 VSSD.n1611 VSSD.n1394 2.63579
R9210 VSSD.n1862 VSSD.n1861 2.63579
R9211 VSSD.n1876 VSSD.n92 2.63579
R9212 VSSD.n2002 VSSD.n11 2.63579
R9213 VSSD.n1989 VSSD.n1988 2.63579
R9214 VSSD.n1971 VSSD.n32 2.63579
R9215 VSSD.n1958 VSSD.n1957 2.63579
R9216 VSSD.n1940 VSSD.n53 2.63579
R9217 VSSD.n1927 VSSD.n1926 2.63579
R9218 VSSD.n1909 VSSD.n74 2.63579
R9219 VSSD.n1896 VSSD.n1895 2.63579
R9220 VSSD.n1279 VSSD.n1278 2.63579
R9221 VSSD.n1244 VSSD.n1243 2.63579
R9222 VSSD.n1209 VSSD.n1208 2.63579
R9223 VSSD.n1174 VSSD.n1173 2.63579
R9224 VSSD.n1139 VSSD.n1138 2.63579
R9225 VSSD.n1104 VSSD.n1103 2.63579
R9226 VSSD.n1069 VSSD.n1068 2.63579
R9227 VSSD.n1034 VSSD.n1033 2.63579
R9228 VSSD.n999 VSSD.n998 2.63579
R9229 VSSD.n964 VSSD.n963 2.63579
R9230 VSSD.n491 VSSD.n473 2.36358
R9231 VSSD.n1659 VSSD.n1378 1.88285
R9232 VSSD.n1694 VSSD.n1693 1.88285
R9233 VSSD.n1730 VSSD.n1355 1.88285
R9234 VSSD.n1765 VSSD.n1764 1.88285
R9235 VSSD.n1801 VSSD.n1332 1.88285
R9236 VSSD.n1463 VSSD.n1462 1.88285
R9237 VSSD.n1499 VSSD.n1498 1.88285
R9238 VSSD.n1533 VSSD.n1418 1.88285
R9239 VSSD.n1569 VSSD.n1568 1.88285
R9240 VSSD.n1605 VSSD.n1604 1.88285
R9241 VSSD.n1870 VSSD.n97 1.88285
R9242 VSSD.n1870 VSSD.n1869 1.88285
R9243 VSSD.n1996 VSSD.n15 1.88285
R9244 VSSD.n1996 VSSD.n1995 1.88285
R9245 VSSD.n1965 VSSD.n36 1.88285
R9246 VSSD.n1965 VSSD.n1964 1.88285
R9247 VSSD.n1934 VSSD.n57 1.88285
R9248 VSSD.n1934 VSSD.n1933 1.88285
R9249 VSSD.n1903 VSSD.n78 1.88285
R9250 VSSD.n1903 VSSD.n1902 1.88285
R9251 VSSD.n1288 VSSD.n1287 1.88285
R9252 VSSD.n1253 VSSD.n1252 1.88285
R9253 VSSD.n1218 VSSD.n1217 1.88285
R9254 VSSD.n1183 VSSD.n1182 1.88285
R9255 VSSD.n1148 VSSD.n1147 1.88285
R9256 VSSD.n1113 VSSD.n1112 1.88285
R9257 VSSD.n1078 VSSD.n1077 1.88285
R9258 VSSD.n1043 VSSD.n1042 1.88285
R9259 VSSD.n1008 VSSD.n1007 1.88285
R9260 VSSD.n973 VSSD.n972 1.88285
R9261 VSSD.n487 VSSD.n486 1.77281
R9262 VSSD.n772 VSSD.n118 1.57588
R9263 VSSD.n495 VSSD.n471 1.47818
R9264 VSSD.n482 VSSD.n477 1.37896
R9265 VSSD.n1823 VSSD.n1822 1.3605
R9266 VSSD.n1826 VSSD.n112 1.3605
R9267 VSSD.n1820 VSSD.n113 1.35908
R9268 VSSD.n468 VSSD.n161 1.18204
R9269 VSSD.n178 VSSD.n175 1.18204
R9270 VSSD.n194 VSSD.n191 1.18204
R9271 VSSD.n213 VSSD.n210 1.18204
R9272 VSSD.n229 VSSD.n226 1.18204
R9273 VSSD.n245 VSSD.n242 1.18204
R9274 VSSD.n777 VSSD.n115 1.18204
R9275 VSSD.n535 VSSD.n534 1.18204
R9276 VSSD.n573 VSSD.n135 1.18204
R9277 VSSD.n761 VSSD.n123 1.18204
R9278 VSSD.n627 VSSD.n624 1.18204
R9279 VSSD.n643 VSSD.n640 1.18204
R9280 VSSD.n450 VSSD.n449 0.985115
R9281 VSSD.n415 VSSD.n414 0.985115
R9282 VSSD.n380 VSSD.n379 0.985115
R9283 VSSD.n345 VSSD.n344 0.985115
R9284 VSSD.n310 VSSD.n309 0.985115
R9285 VSSD.n275 VSSD.n274 0.985115
R9286 VSSD.n515 VSSD.n513 0.985115
R9287 VSSD.n553 VSSD.n552 0.985115
R9288 VSSD.n593 VSSD.n591 0.985115
R9289 VSSD.n743 VSSD.n742 0.985115
R9290 VSSD.n708 VSSD.n707 0.985115
R9291 VSSD.n673 VSSD.n672 0.985115
R9292 VSSD.n464 VSSD.n463 0.788192
R9293 VSSD.n429 VSSD.n428 0.788192
R9294 VSSD.n394 VSSD.n393 0.788192
R9295 VSSD.n359 VSSD.n358 0.788192
R9296 VSSD.n324 VSSD.n323 0.788192
R9297 VSSD.n289 VSSD.n288 0.788192
R9298 VSSD.n783 VSSD.n782 0.788192
R9299 VSSD.n500 VSSD.n499 0.788192
R9300 VSSD.n538 VSSD.n537 0.788192
R9301 VSSD.n578 VSSD.n577 0.788192
R9302 VSSD.n757 VSSD.n756 0.788192
R9303 VSSD.n722 VSSD.n721 0.788192
R9304 VSSD.n687 VSSD.n686 0.788192
R9305 VSSD.n496 VSSD.n495 0.780448
R9306 VSSD.n959 VSSD.n958 0.663075
R9307 VSSD.n1825 VSSD.n1824 0.523938
R9308 VSSD.n1828 VSSD.n110 0.521333
R9309 VSSD.n1821 VSSD.n1819 0.520031
R9310 VSSD.n789 VSSD.n787 0.518729
R9311 VSSD.n1839 VSSD.n107 0.376971
R9312 VSSD.n1314 VSSD.n799 0.376971
R9313 VSSD.n1325 VSSD.n1324 0.234847
R9314 VSSD.n471 VSSD.n470 0.151035
R9315 VSSD.n494 VSSD.n493 0.151035
R9316 VSSD.n1832 VSSD.n1829 0.150766
R9317 VSSD.n1829 VSSD 0.150327
R9318 VSSD.n1446 VSSD.n1445 0.148519
R9319 VSSD.n6 VSSD.n4 0.120292
R9320 VSSD.n7 VSSD.n6 0.120292
R9321 VSSD.n2005 VSSD.n7 0.120292
R9322 VSSD.n2005 VSSD.n2004 0.120292
R9323 VSSD.n2004 VSSD.n2003 0.120292
R9324 VSSD.n2003 VSSD.n9 0.120292
R9325 VSSD.n1999 VSSD.n9 0.120292
R9326 VSSD.n1999 VSSD.n1998 0.120292
R9327 VSSD.n1998 VSSD.n1997 0.120292
R9328 VSSD.n1997 VSSD.n13 0.120292
R9329 VSSD.n1992 VSSD.n13 0.120292
R9330 VSSD.n1992 VSSD.n1991 0.120292
R9331 VSSD.n1991 VSSD.n1990 0.120292
R9332 VSSD.n1990 VSSD.n18 0.120292
R9333 VSSD.n1985 VSSD.n18 0.120292
R9334 VSSD.n1985 VSSD.n1984 0.120292
R9335 VSSD.n1984 VSSD.n1983 0.120292
R9336 VSSD.n1983 VSSD.n21 0.120292
R9337 VSSD.n23 VSSD.n21 0.120292
R9338 VSSD.n27 VSSD.n25 0.120292
R9339 VSSD.n28 VSSD.n27 0.120292
R9340 VSSD.n1974 VSSD.n28 0.120292
R9341 VSSD.n1974 VSSD.n1973 0.120292
R9342 VSSD.n1973 VSSD.n1972 0.120292
R9343 VSSD.n1972 VSSD.n30 0.120292
R9344 VSSD.n1968 VSSD.n30 0.120292
R9345 VSSD.n1968 VSSD.n1967 0.120292
R9346 VSSD.n1967 VSSD.n1966 0.120292
R9347 VSSD.n1966 VSSD.n34 0.120292
R9348 VSSD.n1961 VSSD.n34 0.120292
R9349 VSSD.n1961 VSSD.n1960 0.120292
R9350 VSSD.n1960 VSSD.n1959 0.120292
R9351 VSSD.n1959 VSSD.n39 0.120292
R9352 VSSD.n1954 VSSD.n39 0.120292
R9353 VSSD.n1954 VSSD.n1953 0.120292
R9354 VSSD.n1953 VSSD.n1952 0.120292
R9355 VSSD.n1952 VSSD.n42 0.120292
R9356 VSSD.n44 VSSD.n42 0.120292
R9357 VSSD.n48 VSSD.n46 0.120292
R9358 VSSD.n49 VSSD.n48 0.120292
R9359 VSSD.n1943 VSSD.n49 0.120292
R9360 VSSD.n1943 VSSD.n1942 0.120292
R9361 VSSD.n1942 VSSD.n1941 0.120292
R9362 VSSD.n1941 VSSD.n51 0.120292
R9363 VSSD.n1937 VSSD.n51 0.120292
R9364 VSSD.n1937 VSSD.n1936 0.120292
R9365 VSSD.n1936 VSSD.n1935 0.120292
R9366 VSSD.n1935 VSSD.n55 0.120292
R9367 VSSD.n1930 VSSD.n55 0.120292
R9368 VSSD.n1930 VSSD.n1929 0.120292
R9369 VSSD.n1929 VSSD.n1928 0.120292
R9370 VSSD.n1928 VSSD.n60 0.120292
R9371 VSSD.n1923 VSSD.n60 0.120292
R9372 VSSD.n1923 VSSD.n1922 0.120292
R9373 VSSD.n1922 VSSD.n1921 0.120292
R9374 VSSD.n1921 VSSD.n63 0.120292
R9375 VSSD.n65 VSSD.n63 0.120292
R9376 VSSD.n69 VSSD.n67 0.120292
R9377 VSSD.n70 VSSD.n69 0.120292
R9378 VSSD.n1912 VSSD.n70 0.120292
R9379 VSSD.n1912 VSSD.n1911 0.120292
R9380 VSSD.n1911 VSSD.n1910 0.120292
R9381 VSSD.n1910 VSSD.n72 0.120292
R9382 VSSD.n1906 VSSD.n72 0.120292
R9383 VSSD.n1906 VSSD.n1905 0.120292
R9384 VSSD.n1905 VSSD.n1904 0.120292
R9385 VSSD.n1904 VSSD.n76 0.120292
R9386 VSSD.n1899 VSSD.n76 0.120292
R9387 VSSD.n1899 VSSD.n1898 0.120292
R9388 VSSD.n1898 VSSD.n1897 0.120292
R9389 VSSD.n1897 VSSD.n81 0.120292
R9390 VSSD.n1892 VSSD.n81 0.120292
R9391 VSSD.n1892 VSSD.n1891 0.120292
R9392 VSSD.n1891 VSSD.n1890 0.120292
R9393 VSSD.n1890 VSSD.n84 0.120292
R9394 VSSD.n86 VSSD.n84 0.120292
R9395 VSSD.n1884 VSSD.n1883 0.120292
R9396 VSSD.n1883 VSSD.n1882 0.120292
R9397 VSSD.n1882 VSSD.n90 0.120292
R9398 VSSD.n1878 VSSD.n90 0.120292
R9399 VSSD.n1878 VSSD.n1877 0.120292
R9400 VSSD.n1877 VSSD.n93 0.120292
R9401 VSSD.n1873 VSSD.n93 0.120292
R9402 VSSD.n1873 VSSD.n1872 0.120292
R9403 VSSD.n1872 VSSD.n1871 0.120292
R9404 VSSD.n1871 VSSD.n95 0.120292
R9405 VSSD.n1865 VSSD.n95 0.120292
R9406 VSSD.n1865 VSSD.n1864 0.120292
R9407 VSSD.n1864 VSSD.n1863 0.120292
R9408 VSSD.n1863 VSSD.n99 0.120292
R9409 VSSD.n1857 VSSD.n99 0.120292
R9410 VSSD.n1857 VSSD.n1856 0.120292
R9411 VSSD.n1856 VSSD.n1855 0.120292
R9412 VSSD.n1855 VSSD.n101 0.120292
R9413 VSSD.n1850 VSSD.n101 0.120292
R9414 VSSD.n1848 VSSD.n103 0.120292
R9415 VSSD.n1842 VSSD.n103 0.120292
R9416 VSSD.n1842 VSSD.n1841 0.120292
R9417 VSSD.n1841 VSSD.n1840 0.120292
R9418 VSSD.n1840 VSSD.n105 0.120292
R9419 VSSD.n1834 VSSD.n105 0.120292
R9420 VSSD.n1834 VSSD.n1833 0.120292
R9421 VSSD.n1833 VSSD.n1832 0.120292
R9422 VSSD.n467 VSSD.n466 0.120292
R9423 VSSD.n466 VSSD.n162 0.120292
R9424 VSSD.n461 VSSD.n162 0.120292
R9425 VSSD.n461 VSSD.n460 0.120292
R9426 VSSD.n460 VSSD.n459 0.120292
R9427 VSSD.n459 VSSD.n164 0.120292
R9428 VSSD.n454 VSSD.n164 0.120292
R9429 VSSD.n454 VSSD.n453 0.120292
R9430 VSSD.n453 VSSD.n452 0.120292
R9431 VSSD.n452 VSSD.n167 0.120292
R9432 VSSD.n447 VSSD.n167 0.120292
R9433 VSSD.n447 VSSD.n446 0.120292
R9434 VSSD.n446 VSSD.n445 0.120292
R9435 VSSD.n445 VSSD.n170 0.120292
R9436 VSSD.n441 VSSD.n170 0.120292
R9437 VSSD.n441 VSSD.n440 0.120292
R9438 VSSD.n440 VSSD.n439 0.120292
R9439 VSSD.n439 VSSD.n172 0.120292
R9440 VSSD.n176 VSSD.n172 0.120292
R9441 VSSD.n433 VSSD.n176 0.120292
R9442 VSSD.n432 VSSD.n431 0.120292
R9443 VSSD.n431 VSSD.n177 0.120292
R9444 VSSD.n426 VSSD.n177 0.120292
R9445 VSSD.n426 VSSD.n425 0.120292
R9446 VSSD.n425 VSSD.n424 0.120292
R9447 VSSD.n424 VSSD.n180 0.120292
R9448 VSSD.n419 VSSD.n180 0.120292
R9449 VSSD.n419 VSSD.n418 0.120292
R9450 VSSD.n418 VSSD.n417 0.120292
R9451 VSSD.n417 VSSD.n183 0.120292
R9452 VSSD.n412 VSSD.n183 0.120292
R9453 VSSD.n412 VSSD.n411 0.120292
R9454 VSSD.n411 VSSD.n410 0.120292
R9455 VSSD.n410 VSSD.n186 0.120292
R9456 VSSD.n406 VSSD.n186 0.120292
R9457 VSSD.n406 VSSD.n405 0.120292
R9458 VSSD.n405 VSSD.n404 0.120292
R9459 VSSD.n404 VSSD.n188 0.120292
R9460 VSSD.n192 VSSD.n188 0.120292
R9461 VSSD.n398 VSSD.n192 0.120292
R9462 VSSD.n397 VSSD.n396 0.120292
R9463 VSSD.n396 VSSD.n193 0.120292
R9464 VSSD.n391 VSSD.n193 0.120292
R9465 VSSD.n391 VSSD.n390 0.120292
R9466 VSSD.n390 VSSD.n389 0.120292
R9467 VSSD.n389 VSSD.n196 0.120292
R9468 VSSD.n384 VSSD.n196 0.120292
R9469 VSSD.n384 VSSD.n383 0.120292
R9470 VSSD.n383 VSSD.n382 0.120292
R9471 VSSD.n382 VSSD.n199 0.120292
R9472 VSSD.n377 VSSD.n199 0.120292
R9473 VSSD.n377 VSSD.n376 0.120292
R9474 VSSD.n376 VSSD.n375 0.120292
R9475 VSSD.n375 VSSD.n202 0.120292
R9476 VSSD.n371 VSSD.n202 0.120292
R9477 VSSD.n371 VSSD.n370 0.120292
R9478 VSSD.n370 VSSD.n369 0.120292
R9479 VSSD.n369 VSSD.n204 0.120292
R9480 VSSD.n211 VSSD.n204 0.120292
R9481 VSSD.n363 VSSD.n211 0.120292
R9482 VSSD.n362 VSSD.n361 0.120292
R9483 VSSD.n361 VSSD.n212 0.120292
R9484 VSSD.n356 VSSD.n212 0.120292
R9485 VSSD.n356 VSSD.n355 0.120292
R9486 VSSD.n355 VSSD.n354 0.120292
R9487 VSSD.n354 VSSD.n215 0.120292
R9488 VSSD.n349 VSSD.n215 0.120292
R9489 VSSD.n349 VSSD.n348 0.120292
R9490 VSSD.n348 VSSD.n347 0.120292
R9491 VSSD.n347 VSSD.n218 0.120292
R9492 VSSD.n342 VSSD.n218 0.120292
R9493 VSSD.n342 VSSD.n341 0.120292
R9494 VSSD.n341 VSSD.n340 0.120292
R9495 VSSD.n340 VSSD.n221 0.120292
R9496 VSSD.n336 VSSD.n221 0.120292
R9497 VSSD.n336 VSSD.n335 0.120292
R9498 VSSD.n335 VSSD.n334 0.120292
R9499 VSSD.n334 VSSD.n223 0.120292
R9500 VSSD.n227 VSSD.n223 0.120292
R9501 VSSD.n328 VSSD.n227 0.120292
R9502 VSSD.n327 VSSD.n326 0.120292
R9503 VSSD.n326 VSSD.n228 0.120292
R9504 VSSD.n321 VSSD.n228 0.120292
R9505 VSSD.n321 VSSD.n320 0.120292
R9506 VSSD.n320 VSSD.n319 0.120292
R9507 VSSD.n319 VSSD.n231 0.120292
R9508 VSSD.n314 VSSD.n231 0.120292
R9509 VSSD.n314 VSSD.n313 0.120292
R9510 VSSD.n313 VSSD.n312 0.120292
R9511 VSSD.n312 VSSD.n234 0.120292
R9512 VSSD.n307 VSSD.n234 0.120292
R9513 VSSD.n307 VSSD.n306 0.120292
R9514 VSSD.n306 VSSD.n305 0.120292
R9515 VSSD.n305 VSSD.n237 0.120292
R9516 VSSD.n301 VSSD.n237 0.120292
R9517 VSSD.n301 VSSD.n300 0.120292
R9518 VSSD.n300 VSSD.n299 0.120292
R9519 VSSD.n299 VSSD.n239 0.120292
R9520 VSSD.n243 VSSD.n239 0.120292
R9521 VSSD.n293 VSSD.n243 0.120292
R9522 VSSD.n292 VSSD.n291 0.120292
R9523 VSSD.n291 VSSD.n244 0.120292
R9524 VSSD.n286 VSSD.n244 0.120292
R9525 VSSD.n286 VSSD.n285 0.120292
R9526 VSSD.n285 VSSD.n284 0.120292
R9527 VSSD.n284 VSSD.n247 0.120292
R9528 VSSD.n279 VSSD.n247 0.120292
R9529 VSSD.n279 VSSD.n278 0.120292
R9530 VSSD.n278 VSSD.n277 0.120292
R9531 VSSD.n277 VSSD.n250 0.120292
R9532 VSSD.n272 VSSD.n250 0.120292
R9533 VSSD.n272 VSSD.n271 0.120292
R9534 VSSD.n271 VSSD.n270 0.120292
R9535 VSSD.n270 VSSD.n253 0.120292
R9536 VSSD.n266 VSSD.n253 0.120292
R9537 VSSD.n266 VSSD.n265 0.120292
R9538 VSSD.n265 VSSD.n264 0.120292
R9539 VSSD.n264 VSSD.n255 0.120292
R9540 VSSD.n258 VSSD.n255 0.120292
R9541 VSSD.n259 VSSD.n258 0.120292
R9542 VSSD.n497 VSSD.n496 0.120292
R9543 VSSD.n497 VSSD.n158 0.120292
R9544 VSSD.n502 VSSD.n158 0.120292
R9545 VSSD.n503 VSSD.n502 0.120292
R9546 VSSD.n504 VSSD.n503 0.120292
R9547 VSSD.n504 VSSD.n155 0.120292
R9548 VSSD.n509 VSSD.n155 0.120292
R9549 VSSD.n510 VSSD.n509 0.120292
R9550 VSSD.n511 VSSD.n510 0.120292
R9551 VSSD.n511 VSSD.n153 0.120292
R9552 VSSD.n517 VSSD.n153 0.120292
R9553 VSSD.n518 VSSD.n517 0.120292
R9554 VSSD.n519 VSSD.n518 0.120292
R9555 VSSD.n519 VSSD.n151 0.120292
R9556 VSSD.n523 VSSD.n151 0.120292
R9557 VSSD.n524 VSSD.n523 0.120292
R9558 VSSD.n525 VSSD.n524 0.120292
R9559 VSSD.n525 VSSD.n148 0.120292
R9560 VSSD.n531 VSSD.n148 0.120292
R9561 VSSD.n532 VSSD.n531 0.120292
R9562 VSSD.n533 VSSD.n146 0.120292
R9563 VSSD.n539 VSSD.n146 0.120292
R9564 VSSD.n540 VSSD.n539 0.120292
R9565 VSSD.n541 VSSD.n540 0.120292
R9566 VSSD.n541 VSSD.n143 0.120292
R9567 VSSD.n546 VSSD.n143 0.120292
R9568 VSSD.n547 VSSD.n546 0.120292
R9569 VSSD.n548 VSSD.n547 0.120292
R9570 VSSD.n548 VSSD.n141 0.120292
R9571 VSSD.n554 VSSD.n141 0.120292
R9572 VSSD.n555 VSSD.n554 0.120292
R9573 VSSD.n556 VSSD.n555 0.120292
R9574 VSSD.n556 VSSD.n139 0.120292
R9575 VSSD.n560 VSSD.n139 0.120292
R9576 VSSD.n561 VSSD.n560 0.120292
R9577 VSSD.n562 VSSD.n561 0.120292
R9578 VSSD.n562 VSSD.n137 0.120292
R9579 VSSD.n567 VSSD.n137 0.120292
R9580 VSSD.n570 VSSD.n567 0.120292
R9581 VSSD.n571 VSSD.n570 0.120292
R9582 VSSD.n575 VSSD.n574 0.120292
R9583 VSSD.n575 VSSD.n134 0.120292
R9584 VSSD.n580 VSSD.n134 0.120292
R9585 VSSD.n581 VSSD.n580 0.120292
R9586 VSSD.n582 VSSD.n581 0.120292
R9587 VSSD.n582 VSSD.n131 0.120292
R9588 VSSD.n587 VSSD.n131 0.120292
R9589 VSSD.n588 VSSD.n587 0.120292
R9590 VSSD.n589 VSSD.n588 0.120292
R9591 VSSD.n589 VSSD.n129 0.120292
R9592 VSSD.n595 VSSD.n129 0.120292
R9593 VSSD.n596 VSSD.n595 0.120292
R9594 VSSD.n597 VSSD.n596 0.120292
R9595 VSSD.n597 VSSD.n127 0.120292
R9596 VSSD.n601 VSSD.n127 0.120292
R9597 VSSD.n602 VSSD.n601 0.120292
R9598 VSSD.n603 VSSD.n602 0.120292
R9599 VSSD.n603 VSSD.n124 0.120292
R9600 VSSD.n609 VSSD.n124 0.120292
R9601 VSSD.n610 VSSD.n609 0.120292
R9602 VSSD.n760 VSSD.n759 0.120292
R9603 VSSD.n759 VSSD.n611 0.120292
R9604 VSSD.n754 VSSD.n611 0.120292
R9605 VSSD.n754 VSSD.n753 0.120292
R9606 VSSD.n753 VSSD.n752 0.120292
R9607 VSSD.n752 VSSD.n613 0.120292
R9608 VSSD.n747 VSSD.n613 0.120292
R9609 VSSD.n747 VSSD.n746 0.120292
R9610 VSSD.n746 VSSD.n745 0.120292
R9611 VSSD.n745 VSSD.n616 0.120292
R9612 VSSD.n740 VSSD.n616 0.120292
R9613 VSSD.n740 VSSD.n739 0.120292
R9614 VSSD.n739 VSSD.n738 0.120292
R9615 VSSD.n738 VSSD.n619 0.120292
R9616 VSSD.n734 VSSD.n619 0.120292
R9617 VSSD.n734 VSSD.n733 0.120292
R9618 VSSD.n733 VSSD.n732 0.120292
R9619 VSSD.n732 VSSD.n621 0.120292
R9620 VSSD.n625 VSSD.n621 0.120292
R9621 VSSD.n726 VSSD.n625 0.120292
R9622 VSSD.n725 VSSD.n724 0.120292
R9623 VSSD.n724 VSSD.n626 0.120292
R9624 VSSD.n719 VSSD.n626 0.120292
R9625 VSSD.n719 VSSD.n718 0.120292
R9626 VSSD.n718 VSSD.n717 0.120292
R9627 VSSD.n717 VSSD.n629 0.120292
R9628 VSSD.n712 VSSD.n629 0.120292
R9629 VSSD.n712 VSSD.n711 0.120292
R9630 VSSD.n711 VSSD.n710 0.120292
R9631 VSSD.n710 VSSD.n632 0.120292
R9632 VSSD.n705 VSSD.n632 0.120292
R9633 VSSD.n705 VSSD.n704 0.120292
R9634 VSSD.n704 VSSD.n703 0.120292
R9635 VSSD.n703 VSSD.n635 0.120292
R9636 VSSD.n699 VSSD.n635 0.120292
R9637 VSSD.n699 VSSD.n698 0.120292
R9638 VSSD.n698 VSSD.n697 0.120292
R9639 VSSD.n697 VSSD.n637 0.120292
R9640 VSSD.n641 VSSD.n637 0.120292
R9641 VSSD.n691 VSSD.n641 0.120292
R9642 VSSD.n690 VSSD.n689 0.120292
R9643 VSSD.n689 VSSD.n642 0.120292
R9644 VSSD.n684 VSSD.n642 0.120292
R9645 VSSD.n684 VSSD.n683 0.120292
R9646 VSSD.n683 VSSD.n682 0.120292
R9647 VSSD.n682 VSSD.n645 0.120292
R9648 VSSD.n677 VSSD.n645 0.120292
R9649 VSSD.n677 VSSD.n676 0.120292
R9650 VSSD.n676 VSSD.n675 0.120292
R9651 VSSD.n675 VSSD.n648 0.120292
R9652 VSSD.n670 VSSD.n648 0.120292
R9653 VSSD.n670 VSSD.n669 0.120292
R9654 VSSD.n669 VSSD.n668 0.120292
R9655 VSSD.n668 VSSD.n651 0.120292
R9656 VSSD.n664 VSSD.n651 0.120292
R9657 VSSD.n664 VSSD.n663 0.120292
R9658 VSSD.n663 VSSD.n662 0.120292
R9659 VSSD.n662 VSSD.n653 0.120292
R9660 VSSD.n656 VSSD.n653 0.120292
R9661 VSSD.n657 VSSD.n656 0.120292
R9662 VSSD.n490 VSSD.n489 0.120292
R9663 VSSD.n489 VSSD.n474 0.120292
R9664 VSSD.n484 VSSD.n474 0.120292
R9665 VSSD.n484 VSSD.n483 0.120292
R9666 VSSD.n483 VSSD.n478 0.120292
R9667 VSSD.n478 VSSD.n120 0.120292
R9668 VSSD.n769 VSSD.n120 0.120292
R9669 VSSD.n770 VSSD.n769 0.120292
R9670 VSSD.n774 VSSD.n773 0.120292
R9671 VSSD.n774 VSSD.n116 0.120292
R9672 VSSD.n779 VSSD.n116 0.120292
R9673 VSSD.n780 VSSD.n779 0.120292
R9674 VSSD.n781 VSSD.n114 0.120292
R9675 VSSD.n786 VSSD.n114 0.120292
R9676 VSSD.n1626 VSSD.n1625 0.120292
R9677 VSSD.n1625 VSSD.n1624 0.120292
R9678 VSSD.n1624 VSSD.n1386 0.120292
R9679 VSSD.n1620 VSSD.n1619 0.120292
R9680 VSSD.n1619 VSSD.n1618 0.120292
R9681 VSSD.n1618 VSSD.n1390 0.120292
R9682 VSSD.n1614 VSSD.n1390 0.120292
R9683 VSSD.n1614 VSSD.n1613 0.120292
R9684 VSSD.n1613 VSSD.n1612 0.120292
R9685 VSSD.n1612 VSSD.n1392 0.120292
R9686 VSSD.n1608 VSSD.n1392 0.120292
R9687 VSSD.n1608 VSSD.n1607 0.120292
R9688 VSSD.n1607 VSSD.n1606 0.120292
R9689 VSSD.n1606 VSSD.n1396 0.120292
R9690 VSSD.n1600 VSSD.n1396 0.120292
R9691 VSSD.n1600 VSSD.n1599 0.120292
R9692 VSSD.n1599 VSSD.n1598 0.120292
R9693 VSSD.n1598 VSSD.n1398 0.120292
R9694 VSSD.n1594 VSSD.n1398 0.120292
R9695 VSSD.n1594 VSSD.n1593 0.120292
R9696 VSSD.n1593 VSSD.n1592 0.120292
R9697 VSSD.n1592 VSSD.n1400 0.120292
R9698 VSSD.n1587 VSSD.n1400 0.120292
R9699 VSSD.n1586 VSSD.n1585 0.120292
R9700 VSSD.n1585 VSSD.n1402 0.120292
R9701 VSSD.n1581 VSSD.n1402 0.120292
R9702 VSSD.n1581 VSSD.n1580 0.120292
R9703 VSSD.n1580 VSSD.n1579 0.120292
R9704 VSSD.n1579 VSSD.n1404 0.120292
R9705 VSSD.n1573 VSSD.n1404 0.120292
R9706 VSSD.n1573 VSSD.n1572 0.120292
R9707 VSSD.n1572 VSSD.n1571 0.120292
R9708 VSSD.n1571 VSSD.n1406 0.120292
R9709 VSSD.n1565 VSSD.n1406 0.120292
R9710 VSSD.n1565 VSSD.n1564 0.120292
R9711 VSSD.n1564 VSSD.n1563 0.120292
R9712 VSSD.n1563 VSSD.n1408 0.120292
R9713 VSSD.n1559 VSSD.n1408 0.120292
R9714 VSSD.n1559 VSSD.n1558 0.120292
R9715 VSSD.n1558 VSSD.n1557 0.120292
R9716 VSSD.n1557 VSSD.n1410 0.120292
R9717 VSSD.n1552 VSSD.n1410 0.120292
R9718 VSSD.n1552 VSSD.n1551 0.120292
R9719 VSSD.n1550 VSSD.n1412 0.120292
R9720 VSSD.n1546 VSSD.n1412 0.120292
R9721 VSSD.n1546 VSSD.n1545 0.120292
R9722 VSSD.n1545 VSSD.n1544 0.120292
R9723 VSSD.n1544 VSSD.n1414 0.120292
R9724 VSSD.n1538 VSSD.n1414 0.120292
R9725 VSSD.n1538 VSSD.n1537 0.120292
R9726 VSSD.n1537 VSSD.n1536 0.120292
R9727 VSSD.n1536 VSSD.n1416 0.120292
R9728 VSSD.n1532 VSSD.n1416 0.120292
R9729 VSSD.n1532 VSSD.n1531 0.120292
R9730 VSSD.n1531 VSSD.n1419 0.120292
R9731 VSSD.n1527 VSSD.n1419 0.120292
R9732 VSSD.n1527 VSSD.n1526 0.120292
R9733 VSSD.n1526 VSSD.n1525 0.120292
R9734 VSSD.n1525 VSSD.n1421 0.120292
R9735 VSSD.n1521 VSSD.n1421 0.120292
R9736 VSSD.n1521 VSSD.n1520 0.120292
R9737 VSSD.n1520 VSSD.n1519 0.120292
R9738 VSSD.n1519 VSSD.n1423 0.120292
R9739 VSSD.n1514 VSSD.n1513 0.120292
R9740 VSSD.n1513 VSSD.n1512 0.120292
R9741 VSSD.n1512 VSSD.n1425 0.120292
R9742 VSSD.n1508 VSSD.n1425 0.120292
R9743 VSSD.n1508 VSSD.n1507 0.120292
R9744 VSSD.n1507 VSSD.n1506 0.120292
R9745 VSSD.n1506 VSSD.n1427 0.120292
R9746 VSSD.n1502 VSSD.n1427 0.120292
R9747 VSSD.n1502 VSSD.n1501 0.120292
R9748 VSSD.n1501 VSSD.n1500 0.120292
R9749 VSSD.n1500 VSSD.n1431 0.120292
R9750 VSSD.n1494 VSSD.n1431 0.120292
R9751 VSSD.n1494 VSSD.n1493 0.120292
R9752 VSSD.n1493 VSSD.n1492 0.120292
R9753 VSSD.n1492 VSSD.n1433 0.120292
R9754 VSSD.n1488 VSSD.n1433 0.120292
R9755 VSSD.n1488 VSSD.n1487 0.120292
R9756 VSSD.n1487 VSSD.n1486 0.120292
R9757 VSSD.n1486 VSSD.n1435 0.120292
R9758 VSSD.n1481 VSSD.n1435 0.120292
R9759 VSSD.n1480 VSSD.n1479 0.120292
R9760 VSSD.n1479 VSSD.n1437 0.120292
R9761 VSSD.n1475 VSSD.n1437 0.120292
R9762 VSSD.n1475 VSSD.n1474 0.120292
R9763 VSSD.n1474 VSSD.n1473 0.120292
R9764 VSSD.n1473 VSSD.n1439 0.120292
R9765 VSSD.n1467 VSSD.n1439 0.120292
R9766 VSSD.n1467 VSSD.n1466 0.120292
R9767 VSSD.n1466 VSSD.n1465 0.120292
R9768 VSSD.n1465 VSSD.n1441 0.120292
R9769 VSSD.n1459 VSSD.n1441 0.120292
R9770 VSSD.n1459 VSSD.n1458 0.120292
R9771 VSSD.n1458 VSSD.n1457 0.120292
R9772 VSSD.n1457 VSSD.n1443 0.120292
R9773 VSSD.n1453 VSSD.n1443 0.120292
R9774 VSSD.n1453 VSSD.n1452 0.120292
R9775 VSSD.n1452 VSSD.n1451 0.120292
R9776 VSSD.n1451 VSSD.n1445 0.120292
R9777 VSSD.n1633 VSSD.n1384 0.120292
R9778 VSSD.n1639 VSSD.n1384 0.120292
R9779 VSSD.n1640 VSSD.n1639 0.120292
R9780 VSSD.n1646 VSSD.n1645 0.120292
R9781 VSSD.n1647 VSSD.n1646 0.120292
R9782 VSSD.n1647 VSSD.n1381 0.120292
R9783 VSSD.n1651 VSSD.n1381 0.120292
R9784 VSSD.n1652 VSSD.n1651 0.120292
R9785 VSSD.n1653 VSSD.n1652 0.120292
R9786 VSSD.n1653 VSSD.n1379 0.120292
R9787 VSSD.n1657 VSSD.n1379 0.120292
R9788 VSSD.n1658 VSSD.n1657 0.120292
R9789 VSSD.n1658 VSSD.n1376 0.120292
R9790 VSSD.n1662 VSSD.n1376 0.120292
R9791 VSSD.n1663 VSSD.n1662 0.120292
R9792 VSSD.n1664 VSSD.n1663 0.120292
R9793 VSSD.n1664 VSSD.n1374 0.120292
R9794 VSSD.n1670 VSSD.n1374 0.120292
R9795 VSSD.n1671 VSSD.n1670 0.120292
R9796 VSSD.n1672 VSSD.n1671 0.120292
R9797 VSSD.n1672 VSSD.n1372 0.120292
R9798 VSSD.n1676 VSSD.n1372 0.120292
R9799 VSSD.n1678 VSSD.n1369 0.120292
R9800 VSSD.n1682 VSSD.n1369 0.120292
R9801 VSSD.n1683 VSSD.n1682 0.120292
R9802 VSSD.n1684 VSSD.n1683 0.120292
R9803 VSSD.n1684 VSSD.n1367 0.120292
R9804 VSSD.n1688 VSSD.n1367 0.120292
R9805 VSSD.n1689 VSSD.n1688 0.120292
R9806 VSSD.n1690 VSSD.n1689 0.120292
R9807 VSSD.n1690 VSSD.n1365 0.120292
R9808 VSSD.n1696 VSSD.n1365 0.120292
R9809 VSSD.n1697 VSSD.n1696 0.120292
R9810 VSSD.n1698 VSSD.n1697 0.120292
R9811 VSSD.n1698 VSSD.n1363 0.120292
R9812 VSSD.n1704 VSSD.n1363 0.120292
R9813 VSSD.n1705 VSSD.n1704 0.120292
R9814 VSSD.n1706 VSSD.n1705 0.120292
R9815 VSSD.n1706 VSSD.n1361 0.120292
R9816 VSSD.n1710 VSSD.n1361 0.120292
R9817 VSSD.n1711 VSSD.n1710 0.120292
R9818 VSSD.n1717 VSSD.n1716 0.120292
R9819 VSSD.n1718 VSSD.n1717 0.120292
R9820 VSSD.n1718 VSSD.n1358 0.120292
R9821 VSSD.n1722 VSSD.n1358 0.120292
R9822 VSSD.n1723 VSSD.n1722 0.120292
R9823 VSSD.n1724 VSSD.n1723 0.120292
R9824 VSSD.n1724 VSSD.n1356 0.120292
R9825 VSSD.n1728 VSSD.n1356 0.120292
R9826 VSSD.n1729 VSSD.n1728 0.120292
R9827 VSSD.n1729 VSSD.n1353 0.120292
R9828 VSSD.n1733 VSSD.n1353 0.120292
R9829 VSSD.n1734 VSSD.n1733 0.120292
R9830 VSSD.n1735 VSSD.n1734 0.120292
R9831 VSSD.n1735 VSSD.n1351 0.120292
R9832 VSSD.n1741 VSSD.n1351 0.120292
R9833 VSSD.n1742 VSSD.n1741 0.120292
R9834 VSSD.n1743 VSSD.n1742 0.120292
R9835 VSSD.n1743 VSSD.n1349 0.120292
R9836 VSSD.n1747 VSSD.n1349 0.120292
R9837 VSSD.n1749 VSSD.n1346 0.120292
R9838 VSSD.n1753 VSSD.n1346 0.120292
R9839 VSSD.n1754 VSSD.n1753 0.120292
R9840 VSSD.n1755 VSSD.n1754 0.120292
R9841 VSSD.n1755 VSSD.n1344 0.120292
R9842 VSSD.n1759 VSSD.n1344 0.120292
R9843 VSSD.n1760 VSSD.n1759 0.120292
R9844 VSSD.n1761 VSSD.n1760 0.120292
R9845 VSSD.n1761 VSSD.n1342 0.120292
R9846 VSSD.n1767 VSSD.n1342 0.120292
R9847 VSSD.n1768 VSSD.n1767 0.120292
R9848 VSSD.n1769 VSSD.n1768 0.120292
R9849 VSSD.n1769 VSSD.n1340 0.120292
R9850 VSSD.n1775 VSSD.n1340 0.120292
R9851 VSSD.n1776 VSSD.n1775 0.120292
R9852 VSSD.n1777 VSSD.n1776 0.120292
R9853 VSSD.n1777 VSSD.n1338 0.120292
R9854 VSSD.n1781 VSSD.n1338 0.120292
R9855 VSSD.n1782 VSSD.n1781 0.120292
R9856 VSSD.n1788 VSSD.n1787 0.120292
R9857 VSSD.n1789 VSSD.n1788 0.120292
R9858 VSSD.n1789 VSSD.n1335 0.120292
R9859 VSSD.n1793 VSSD.n1335 0.120292
R9860 VSSD.n1794 VSSD.n1793 0.120292
R9861 VSSD.n1795 VSSD.n1794 0.120292
R9862 VSSD.n1795 VSSD.n1333 0.120292
R9863 VSSD.n1799 VSSD.n1333 0.120292
R9864 VSSD.n1800 VSSD.n1799 0.120292
R9865 VSSD.n1800 VSSD.n1330 0.120292
R9866 VSSD.n1804 VSSD.n1330 0.120292
R9867 VSSD.n1805 VSSD.n1804 0.120292
R9868 VSSD.n1806 VSSD.n1805 0.120292
R9869 VSSD.n1806 VSSD.n1328 0.120292
R9870 VSSD.n1812 VSSD.n1328 0.120292
R9871 VSSD.n1813 VSSD.n1812 0.120292
R9872 VSSD.n1814 VSSD.n1813 0.120292
R9873 VSSD.n1814 VSSD.n1326 0.120292
R9874 VSSD.n1818 VSSD.n1326 0.120292
R9875 VSSD.n960 VSSD.n959 0.120292
R9876 VSSD.n960 VSSD.n952 0.120292
R9877 VSSD.n965 VSSD.n952 0.120292
R9878 VSSD.n966 VSSD.n965 0.120292
R9879 VSSD.n967 VSSD.n966 0.120292
R9880 VSSD.n967 VSSD.n950 0.120292
R9881 VSSD.n974 VSSD.n950 0.120292
R9882 VSSD.n975 VSSD.n974 0.120292
R9883 VSSD.n976 VSSD.n975 0.120292
R9884 VSSD.n976 VSSD.n948 0.120292
R9885 VSSD.n980 VSSD.n948 0.120292
R9886 VSSD.n981 VSSD.n980 0.120292
R9887 VSSD.n982 VSSD.n981 0.120292
R9888 VSSD.n982 VSSD.n946 0.120292
R9889 VSSD.n986 VSSD.n946 0.120292
R9890 VSSD.n987 VSSD.n986 0.120292
R9891 VSSD.n988 VSSD.n987 0.120292
R9892 VSSD.n942 VSSD.n941 0.120292
R9893 VSSD.n993 VSSD.n941 0.120292
R9894 VSSD.n994 VSSD.n993 0.120292
R9895 VSSD.n995 VSSD.n994 0.120292
R9896 VSSD.n995 VSSD.n937 0.120292
R9897 VSSD.n1000 VSSD.n937 0.120292
R9898 VSSD.n1001 VSSD.n1000 0.120292
R9899 VSSD.n1002 VSSD.n1001 0.120292
R9900 VSSD.n1002 VSSD.n935 0.120292
R9901 VSSD.n1009 VSSD.n935 0.120292
R9902 VSSD.n1010 VSSD.n1009 0.120292
R9903 VSSD.n1011 VSSD.n1010 0.120292
R9904 VSSD.n1011 VSSD.n933 0.120292
R9905 VSSD.n1015 VSSD.n933 0.120292
R9906 VSSD.n1016 VSSD.n1015 0.120292
R9907 VSSD.n1017 VSSD.n1016 0.120292
R9908 VSSD.n1017 VSSD.n931 0.120292
R9909 VSSD.n1021 VSSD.n931 0.120292
R9910 VSSD.n1022 VSSD.n1021 0.120292
R9911 VSSD.n1023 VSSD.n1022 0.120292
R9912 VSSD.n927 VSSD.n926 0.120292
R9913 VSSD.n1028 VSSD.n926 0.120292
R9914 VSSD.n1029 VSSD.n1028 0.120292
R9915 VSSD.n1030 VSSD.n1029 0.120292
R9916 VSSD.n1030 VSSD.n922 0.120292
R9917 VSSD.n1035 VSSD.n922 0.120292
R9918 VSSD.n1036 VSSD.n1035 0.120292
R9919 VSSD.n1037 VSSD.n1036 0.120292
R9920 VSSD.n1037 VSSD.n920 0.120292
R9921 VSSD.n1044 VSSD.n920 0.120292
R9922 VSSD.n1045 VSSD.n1044 0.120292
R9923 VSSD.n1046 VSSD.n1045 0.120292
R9924 VSSD.n1046 VSSD.n918 0.120292
R9925 VSSD.n1050 VSSD.n918 0.120292
R9926 VSSD.n1051 VSSD.n1050 0.120292
R9927 VSSD.n1052 VSSD.n1051 0.120292
R9928 VSSD.n1052 VSSD.n916 0.120292
R9929 VSSD.n1056 VSSD.n916 0.120292
R9930 VSSD.n1057 VSSD.n1056 0.120292
R9931 VSSD.n1058 VSSD.n1057 0.120292
R9932 VSSD.n912 VSSD.n911 0.120292
R9933 VSSD.n1063 VSSD.n911 0.120292
R9934 VSSD.n1064 VSSD.n1063 0.120292
R9935 VSSD.n1065 VSSD.n1064 0.120292
R9936 VSSD.n1065 VSSD.n907 0.120292
R9937 VSSD.n1070 VSSD.n907 0.120292
R9938 VSSD.n1071 VSSD.n1070 0.120292
R9939 VSSD.n1072 VSSD.n1071 0.120292
R9940 VSSD.n1072 VSSD.n905 0.120292
R9941 VSSD.n1079 VSSD.n905 0.120292
R9942 VSSD.n1080 VSSD.n1079 0.120292
R9943 VSSD.n1081 VSSD.n1080 0.120292
R9944 VSSD.n1081 VSSD.n903 0.120292
R9945 VSSD.n1085 VSSD.n903 0.120292
R9946 VSSD.n1086 VSSD.n1085 0.120292
R9947 VSSD.n1087 VSSD.n1086 0.120292
R9948 VSSD.n1087 VSSD.n901 0.120292
R9949 VSSD.n1091 VSSD.n901 0.120292
R9950 VSSD.n1092 VSSD.n1091 0.120292
R9951 VSSD.n1093 VSSD.n1092 0.120292
R9952 VSSD.n897 VSSD.n896 0.120292
R9953 VSSD.n1098 VSSD.n896 0.120292
R9954 VSSD.n1099 VSSD.n1098 0.120292
R9955 VSSD.n1100 VSSD.n1099 0.120292
R9956 VSSD.n1100 VSSD.n892 0.120292
R9957 VSSD.n1105 VSSD.n892 0.120292
R9958 VSSD.n1106 VSSD.n1105 0.120292
R9959 VSSD.n1107 VSSD.n1106 0.120292
R9960 VSSD.n1107 VSSD.n890 0.120292
R9961 VSSD.n1114 VSSD.n890 0.120292
R9962 VSSD.n1115 VSSD.n1114 0.120292
R9963 VSSD.n1116 VSSD.n1115 0.120292
R9964 VSSD.n1116 VSSD.n888 0.120292
R9965 VSSD.n1120 VSSD.n888 0.120292
R9966 VSSD.n1121 VSSD.n1120 0.120292
R9967 VSSD.n1122 VSSD.n1121 0.120292
R9968 VSSD.n1122 VSSD.n886 0.120292
R9969 VSSD.n1126 VSSD.n886 0.120292
R9970 VSSD.n1127 VSSD.n1126 0.120292
R9971 VSSD.n1128 VSSD.n1127 0.120292
R9972 VSSD.n882 VSSD.n881 0.120292
R9973 VSSD.n1133 VSSD.n881 0.120292
R9974 VSSD.n1134 VSSD.n1133 0.120292
R9975 VSSD.n1135 VSSD.n1134 0.120292
R9976 VSSD.n1135 VSSD.n877 0.120292
R9977 VSSD.n1140 VSSD.n877 0.120292
R9978 VSSD.n1141 VSSD.n1140 0.120292
R9979 VSSD.n1142 VSSD.n1141 0.120292
R9980 VSSD.n1142 VSSD.n875 0.120292
R9981 VSSD.n1149 VSSD.n875 0.120292
R9982 VSSD.n1150 VSSD.n1149 0.120292
R9983 VSSD.n1151 VSSD.n1150 0.120292
R9984 VSSD.n1151 VSSD.n873 0.120292
R9985 VSSD.n1155 VSSD.n873 0.120292
R9986 VSSD.n1156 VSSD.n1155 0.120292
R9987 VSSD.n1157 VSSD.n1156 0.120292
R9988 VSSD.n1157 VSSD.n871 0.120292
R9989 VSSD.n1161 VSSD.n871 0.120292
R9990 VSSD.n1162 VSSD.n1161 0.120292
R9991 VSSD.n1163 VSSD.n1162 0.120292
R9992 VSSD.n867 VSSD.n866 0.120292
R9993 VSSD.n1168 VSSD.n866 0.120292
R9994 VSSD.n1169 VSSD.n1168 0.120292
R9995 VSSD.n1170 VSSD.n1169 0.120292
R9996 VSSD.n1170 VSSD.n862 0.120292
R9997 VSSD.n1175 VSSD.n862 0.120292
R9998 VSSD.n1176 VSSD.n1175 0.120292
R9999 VSSD.n1177 VSSD.n1176 0.120292
R10000 VSSD.n1177 VSSD.n860 0.120292
R10001 VSSD.n1184 VSSD.n860 0.120292
R10002 VSSD.n1185 VSSD.n1184 0.120292
R10003 VSSD.n1186 VSSD.n1185 0.120292
R10004 VSSD.n1186 VSSD.n858 0.120292
R10005 VSSD.n1190 VSSD.n858 0.120292
R10006 VSSD.n1191 VSSD.n1190 0.120292
R10007 VSSD.n1192 VSSD.n1191 0.120292
R10008 VSSD.n1192 VSSD.n856 0.120292
R10009 VSSD.n1196 VSSD.n856 0.120292
R10010 VSSD.n1197 VSSD.n1196 0.120292
R10011 VSSD.n1198 VSSD.n1197 0.120292
R10012 VSSD.n852 VSSD.n851 0.120292
R10013 VSSD.n1203 VSSD.n851 0.120292
R10014 VSSD.n1204 VSSD.n1203 0.120292
R10015 VSSD.n1205 VSSD.n1204 0.120292
R10016 VSSD.n1205 VSSD.n847 0.120292
R10017 VSSD.n1210 VSSD.n847 0.120292
R10018 VSSD.n1211 VSSD.n1210 0.120292
R10019 VSSD.n1212 VSSD.n1211 0.120292
R10020 VSSD.n1212 VSSD.n845 0.120292
R10021 VSSD.n1219 VSSD.n845 0.120292
R10022 VSSD.n1220 VSSD.n1219 0.120292
R10023 VSSD.n1221 VSSD.n1220 0.120292
R10024 VSSD.n1221 VSSD.n843 0.120292
R10025 VSSD.n1225 VSSD.n843 0.120292
R10026 VSSD.n1226 VSSD.n1225 0.120292
R10027 VSSD.n1227 VSSD.n1226 0.120292
R10028 VSSD.n1227 VSSD.n841 0.120292
R10029 VSSD.n1231 VSSD.n841 0.120292
R10030 VSSD.n1232 VSSD.n1231 0.120292
R10031 VSSD.n1233 VSSD.n1232 0.120292
R10032 VSSD.n837 VSSD.n836 0.120292
R10033 VSSD.n1238 VSSD.n836 0.120292
R10034 VSSD.n1239 VSSD.n1238 0.120292
R10035 VSSD.n1240 VSSD.n1239 0.120292
R10036 VSSD.n1240 VSSD.n832 0.120292
R10037 VSSD.n1245 VSSD.n832 0.120292
R10038 VSSD.n1246 VSSD.n1245 0.120292
R10039 VSSD.n1247 VSSD.n1246 0.120292
R10040 VSSD.n1247 VSSD.n830 0.120292
R10041 VSSD.n1254 VSSD.n830 0.120292
R10042 VSSD.n1255 VSSD.n1254 0.120292
R10043 VSSD.n1256 VSSD.n1255 0.120292
R10044 VSSD.n1256 VSSD.n828 0.120292
R10045 VSSD.n1260 VSSD.n828 0.120292
R10046 VSSD.n1261 VSSD.n1260 0.120292
R10047 VSSD.n1262 VSSD.n1261 0.120292
R10048 VSSD.n1262 VSSD.n826 0.120292
R10049 VSSD.n1266 VSSD.n826 0.120292
R10050 VSSD.n1267 VSSD.n1266 0.120292
R10051 VSSD.n1268 VSSD.n1267 0.120292
R10052 VSSD.n822 VSSD.n821 0.120292
R10053 VSSD.n1273 VSSD.n821 0.120292
R10054 VSSD.n1274 VSSD.n1273 0.120292
R10055 VSSD.n1275 VSSD.n1274 0.120292
R10056 VSSD.n1275 VSSD.n817 0.120292
R10057 VSSD.n1280 VSSD.n817 0.120292
R10058 VSSD.n1281 VSSD.n1280 0.120292
R10059 VSSD.n1282 VSSD.n1281 0.120292
R10060 VSSD.n1282 VSSD.n815 0.120292
R10061 VSSD.n1289 VSSD.n815 0.120292
R10062 VSSD.n1290 VSSD.n1289 0.120292
R10063 VSSD.n1291 VSSD.n1290 0.120292
R10064 VSSD.n1291 VSSD.n813 0.120292
R10065 VSSD.n1295 VSSD.n813 0.120292
R10066 VSSD.n1296 VSSD.n1295 0.120292
R10067 VSSD.n1297 VSSD.n1296 0.120292
R10068 VSSD.n1297 VSSD.n811 0.120292
R10069 VSSD.n811 VSSD.n808 0.120292
R10070 VSSD.n1302 VSSD.n808 0.120292
R10071 VSSD.n1303 VSSD.n1302 0.120292
R10072 VSSD.n1304 VSSD.n806 0.120292
R10073 VSSD.n1308 VSSD.n806 0.120292
R10074 VSSD.n1309 VSSD.n1308 0.120292
R10075 VSSD.n1310 VSSD.n1309 0.120292
R10076 VSSD.n1310 VSSD.n800 0.120292
R10077 VSSD.n1315 VSSD.n800 0.120292
R10078 VSSD.n1316 VSSD.n1315 0.120292
R10079 VSSD.n1316 VSSD.n795 0.120292
R10080 VSSD.n795 VSSD.n791 0.120292
R10081 VSSD.n1321 VSSD.n791 0.120292
R10082 VSSD.n1322 VSSD.n1321 0.120292
R10083 VSSD.n1446 VSSD 0.114842
R10084 VSSD.n4 VSSD 0.0981562
R10085 VSSD.n25 VSSD 0.0981562
R10086 VSSD.n46 VSSD 0.0981562
R10087 VSSD.n67 VSSD 0.0981562
R10088 VSSD.n1884 VSSD 0.0981562
R10089 VSSD.n1626 VSSD 0.0981562
R10090 VSSD.n1633 VSSD 0.0981562
R10091 VSSD.n1645 VSSD 0.0981562
R10092 VSSD.n1678 VSSD 0.0981562
R10093 VSSD.n1716 VSSD 0.0981562
R10094 VSSD.n1749 VSSD 0.0981562
R10095 VSSD.n1787 VSSD 0.0981562
R10096 VSSD VSSD.n1848 0.0968542
R10097 VSSD.n24 VSSD 0.0603958
R10098 VSSD.n45 VSSD 0.0603958
R10099 VSSD.n66 VSSD 0.0603958
R10100 VSSD.n87 VSSD 0.0603958
R10101 VSSD.n467 VSSD 0.0603958
R10102 VSSD VSSD.n432 0.0603958
R10103 VSSD VSSD.n397 0.0603958
R10104 VSSD VSSD.n362 0.0603958
R10105 VSSD VSSD.n327 0.0603958
R10106 VSSD VSSD.n292 0.0603958
R10107 VSSD.n533 VSSD 0.0603958
R10108 VSSD.n574 VSSD 0.0603958
R10109 VSSD.n760 VSSD 0.0603958
R10110 VSSD VSSD.n725 0.0603958
R10111 VSSD VSSD.n690 0.0603958
R10112 VSSD.n490 VSSD 0.0603958
R10113 VSSD.n773 VSSD 0.0603958
R10114 VSSD.n781 VSSD 0.0603958
R10115 VSSD VSSD.n1386 0.0603958
R10116 VSSD VSSD.n1586 0.0603958
R10117 VSSD VSSD.n1550 0.0603958
R10118 VSSD.n1514 VSSD 0.0603958
R10119 VSSD VSSD.n1480 0.0603958
R10120 VSSD VSSD.n1640 0.0603958
R10121 VSSD VSSD.n1676 0.0603958
R10122 VSSD.n1677 VSSD 0.0603958
R10123 VSSD VSSD.n1711 0.0603958
R10124 VSSD.n1712 VSSD 0.0603958
R10125 VSSD VSSD.n1747 0.0603958
R10126 VSSD.n1748 VSSD 0.0603958
R10127 VSSD VSSD.n1782 0.0603958
R10128 VSSD.n1783 VSSD 0.0603958
R10129 VSSD VSSD.n1818 0.0603958
R10130 VSSD VSSD.n942 0.0603958
R10131 VSSD VSSD.n927 0.0603958
R10132 VSSD VSSD.n912 0.0603958
R10133 VSSD VSSD.n897 0.0603958
R10134 VSSD VSSD.n882 0.0603958
R10135 VSSD VSSD.n867 0.0603958
R10136 VSSD VSSD.n852 0.0603958
R10137 VSSD VSSD.n837 0.0603958
R10138 VSSD VSSD.n822 0.0603958
R10139 VSSD.n1304 VSSD 0.0603958
R10140 VSSD VSSD.n1849 0.0590938
R10141 VSSD.n1620 VSSD 0.0590938
R10142 VSSD.n1641 VSSD 0.0590938
R10143 VSSD.n1849 VSSD 0.0239375
R10144 VSSD.n2011 VSSD 0.0226354
R10145 VSSD VSSD.n23 0.0226354
R10146 VSSD VSSD.n24 0.0226354
R10147 VSSD VSSD.n44 0.0226354
R10148 VSSD VSSD.n45 0.0226354
R10149 VSSD VSSD.n65 0.0226354
R10150 VSSD VSSD.n66 0.0226354
R10151 VSSD VSSD.n86 0.0226354
R10152 VSSD VSSD.n87 0.0226354
R10153 VSSD.n1850 VSSD 0.0226354
R10154 VSSD.n470 VSSD 0.0226354
R10155 VSSD.n433 VSSD 0.0226354
R10156 VSSD.n398 VSSD 0.0226354
R10157 VSSD.n363 VSSD 0.0226354
R10158 VSSD.n328 VSSD 0.0226354
R10159 VSSD.n293 VSSD 0.0226354
R10160 VSSD.n259 VSSD 0.0226354
R10161 VSSD VSSD.n532 0.0226354
R10162 VSSD.n571 VSSD 0.0226354
R10163 VSSD VSSD.n610 0.0226354
R10164 VSSD.n726 VSSD 0.0226354
R10165 VSSD.n691 VSSD 0.0226354
R10166 VSSD.n657 VSSD 0.0226354
R10167 VSSD.n493 VSSD 0.0226354
R10168 VSSD.n770 VSSD 0.0226354
R10169 VSSD VSSD.n780 0.0226354
R10170 VSSD VSSD.n786 0.0226354
R10171 VSSD.n1628 VSSD 0.0226354
R10172 VSSD.n1587 VSSD 0.0226354
R10173 VSSD.n1551 VSSD 0.0226354
R10174 VSSD VSSD.n1423 0.0226354
R10175 VSSD.n1481 VSSD 0.0226354
R10176 VSSD VSSD.n1632 0.0226354
R10177 VSSD.n1641 VSSD 0.0226354
R10178 VSSD VSSD.n1677 0.0226354
R10179 VSSD.n1712 VSSD 0.0226354
R10180 VSSD VSSD.n1748 0.0226354
R10181 VSSD.n1783 VSSD 0.0226354
R10182 VSSD.n988 VSSD 0.0226354
R10183 VSSD.n1023 VSSD 0.0226354
R10184 VSSD.n1058 VSSD 0.0226354
R10185 VSSD.n1093 VSSD 0.0226354
R10186 VSSD.n1128 VSSD 0.0226354
R10187 VSSD.n1163 VSSD 0.0226354
R10188 VSSD.n1198 VSSD 0.0226354
R10189 VSSD.n1233 VSSD 0.0226354
R10190 VSSD.n1268 VSSD 0.0226354
R10191 VSSD VSSD.n1303 0.0226354
R10192 VSSD.n1323 VSSD 0.0148229
R10193 VSSD.n1323 VSSD.n1322 0.00701042
R10194 a_5911_n5372.n3 a_5911_n5372.n2 636.953
R10195 a_5911_n5372.n1 a_5911_n5372.t5 366.856
R10196 a_5911_n5372.n2 a_5911_n5372.n0 300.2
R10197 a_5911_n5372.n2 a_5911_n5372.n1 225.036
R10198 a_5911_n5372.n1 a_5911_n5372.t4 174.056
R10199 a_5911_n5372.n0 a_5911_n5372.t3 70.0005
R10200 a_5911_n5372.t1 a_5911_n5372.n3 68.0124
R10201 a_5911_n5372.n3 a_5911_n5372.t2 63.3219
R10202 a_5911_n5372.n0 a_5911_n5372.t0 61.6672
R10203 a_5624_n5650.n5 a_5624_n5650.n4 807.871
R10204 a_5624_n5650.n0 a_5624_n5650.t3 389.183
R10205 a_5624_n5650.n1 a_5624_n5650.n0 251.167
R10206 a_5624_n5650.n1 a_5624_n5650.t2 223.571
R10207 a_5624_n5650.n3 a_5624_n5650.t8 212.081
R10208 a_5624_n5650.n2 a_5624_n5650.t7 212.081
R10209 a_5624_n5650.n4 a_5624_n5650.n3 176.576
R10210 a_5624_n5650.n0 a_5624_n5650.t5 174.891
R10211 a_5624_n5650.n3 a_5624_n5650.t6 139.78
R10212 a_5624_n5650.n2 a_5624_n5650.t4 139.78
R10213 a_5624_n5650.t0 a_5624_n5650.n5 63.3219
R10214 a_5624_n5650.n5 a_5624_n5650.t1 63.3219
R10215 a_5624_n5650.n3 a_5624_n5650.n2 61.346
R10216 a_5624_n5650.n4 a_5624_n5650.n1 37.5061
R10217 a_2155_3557.n1 a_2155_3557.t3 530.01
R10218 a_2155_3557.t0 a_2155_3557.n5 421.021
R10219 a_2155_3557.n0 a_2155_3557.t2 337.142
R10220 a_2155_3557.n3 a_2155_3557.t1 280.223
R10221 a_2155_3557.n4 a_2155_3557.t5 263.173
R10222 a_2155_3557.n4 a_2155_3557.t6 227.826
R10223 a_2155_3557.n0 a_2155_3557.t7 199.762
R10224 a_2155_3557.n2 a_2155_3557.n1 170.81
R10225 a_2155_3557.n2 a_2155_3557.n0 167.321
R10226 a_2155_3557.n5 a_2155_3557.n4 152
R10227 a_2155_3557.n1 a_2155_3557.t4 141.923
R10228 a_2155_3557.n3 a_2155_3557.n2 10.8376
R10229 a_2155_3557.n5 a_2155_3557.n3 2.50485
R10230 a_2889_3799.n3 a_2889_3799.n2 647.119
R10231 a_2889_3799.n1 a_2889_3799.t4 350.253
R10232 a_2889_3799.n2 a_2889_3799.n0 260.339
R10233 a_2889_3799.n2 a_2889_3799.n1 246.119
R10234 a_2889_3799.n1 a_2889_3799.t5 189.588
R10235 a_2889_3799.n3 a_2889_3799.t3 89.1195
R10236 a_2889_3799.n0 a_2889_3799.t2 63.3338
R10237 a_2889_3799.t0 a_2889_3799.n3 41.0422
R10238 a_2889_3799.n0 a_2889_3799.t1 31.9797
R10239 a_3236_3557.n3 a_3236_3557.n2 636.953
R10240 a_3236_3557.n1 a_3236_3557.t5 366.856
R10241 a_3236_3557.n2 a_3236_3557.n0 300.2
R10242 a_3236_3557.n2 a_3236_3557.n1 225.036
R10243 a_3236_3557.n1 a_3236_3557.t4 174.056
R10244 a_3236_3557.n0 a_3236_3557.t0 70.0005
R10245 a_3236_3557.t2 a_3236_3557.n3 68.0124
R10246 a_3236_3557.n3 a_3236_3557.t3 63.3219
R10247 a_3236_3557.n0 a_3236_3557.t1 61.6672
R10248 a_4679_n663.n0 a_4679_n663.t2 1327.82
R10249 a_4679_n663.t0 a_4679_n663.n0 194.655
R10250 a_4679_n663.n0 a_4679_n663.t1 63.3219
R10251 cdac_ctrl_0.x2.X.n31 cdac_ctrl_0.x2.X.n30 374.966
R10252 cdac_ctrl_0.x2.X.n18 cdac_ctrl_0.x2.X.t31 333.651
R10253 cdac_ctrl_0.x2.X.n16 cdac_ctrl_0.x2.X.t35 333.651
R10254 cdac_ctrl_0.x2.X.n14 cdac_ctrl_0.x2.X.t20 333.651
R10255 cdac_ctrl_0.x2.X.n12 cdac_ctrl_0.x2.X.t24 333.651
R10256 cdac_ctrl_0.x2.X.n10 cdac_ctrl_0.x2.X.t29 333.651
R10257 cdac_ctrl_0.x2.X.n8 cdac_ctrl_0.x2.X.t18 333.651
R10258 cdac_ctrl_0.x2.X.n6 cdac_ctrl_0.x2.X.t32 333.651
R10259 cdac_ctrl_0.x2.X.n4 cdac_ctrl_0.x2.X.t33 333.651
R10260 cdac_ctrl_0.x2.X.n2 cdac_ctrl_0.x2.X.t25 333.651
R10261 cdac_ctrl_0.x2.X.n1 cdac_ctrl_0.x2.X.t16 333.651
R10262 cdac_ctrl_0.x2.X.n31 cdac_ctrl_0.x2.X.n29 311.719
R10263 cdac_ctrl_0.x2.X.n32 cdac_ctrl_0.x2.X.n28 311.719
R10264 cdac_ctrl_0.x2.X.n18 cdac_ctrl_0.x2.X.t17 297.233
R10265 cdac_ctrl_0.x2.X.n16 cdac_ctrl_0.x2.X.t23 297.233
R10266 cdac_ctrl_0.x2.X.n14 cdac_ctrl_0.x2.X.t19 297.233
R10267 cdac_ctrl_0.x2.X.n12 cdac_ctrl_0.x2.X.t22 297.233
R10268 cdac_ctrl_0.x2.X.n10 cdac_ctrl_0.x2.X.t26 297.233
R10269 cdac_ctrl_0.x2.X.n8 cdac_ctrl_0.x2.X.t28 297.233
R10270 cdac_ctrl_0.x2.X.n6 cdac_ctrl_0.x2.X.t34 297.233
R10271 cdac_ctrl_0.x2.X.n4 cdac_ctrl_0.x2.X.t27 297.233
R10272 cdac_ctrl_0.x2.X.n2 cdac_ctrl_0.x2.X.t30 297.233
R10273 cdac_ctrl_0.x2.X.n1 cdac_ctrl_0.x2.X.t21 297.233
R10274 cdac_ctrl_0.x2.X.n20 cdac_ctrl_0.x2.X.n0 284.19
R10275 cdac_ctrl_0.x2.X.n24 cdac_ctrl_0.x2.X.n23 261.425
R10276 cdac_ctrl_0.x2.X.n27 cdac_ctrl_0.x2.X.n26 202.444
R10277 cdac_ctrl_0.x2.X.n25 cdac_ctrl_0.x2.X.n21 198.177
R10278 cdac_ctrl_0.x2.X.n24 cdac_ctrl_0.x2.X.n22 198.177
R10279 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n18 196.493
R10280 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n16 196.493
R10281 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n14 196.493
R10282 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n12 196.493
R10283 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n10 196.493
R10284 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n8 196.493
R10285 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n6 196.493
R10286 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n4 196.493
R10287 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n2 196.493
R10288 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n1 196.493
R10289 cdac_ctrl_0.x2.X.n25 cdac_ctrl_0.x2.X.n24 63.2476
R10290 cdac_ctrl_0.x2.X.n32 cdac_ctrl_0.x2.X.n31 63.2476
R10291 cdac_ctrl_0.x2.X.n27 cdac_ctrl_0.x2.X.n25 50.4476
R10292 cdac_ctrl_0.x2.X.n33 cdac_ctrl_0.x2.X.n32 50.4476
R10293 cdac_ctrl_0.x2.X.n3 cdac_ctrl_0.x2.X 38.2063
R10294 cdac_ctrl_0.x2.X.n3 cdac_ctrl_0.x2.X 31.159
R10295 cdac_ctrl_0.x2.X.n5 cdac_ctrl_0.x2.X 31.159
R10296 cdac_ctrl_0.x2.X.n7 cdac_ctrl_0.x2.X 31.159
R10297 cdac_ctrl_0.x2.X.n9 cdac_ctrl_0.x2.X 31.159
R10298 cdac_ctrl_0.x2.X.n11 cdac_ctrl_0.x2.X 31.159
R10299 cdac_ctrl_0.x2.X.n13 cdac_ctrl_0.x2.X 31.159
R10300 cdac_ctrl_0.x2.X.n15 cdac_ctrl_0.x2.X 31.159
R10301 cdac_ctrl_0.x2.X.n17 cdac_ctrl_0.x2.X 31.159
R10302 cdac_ctrl_0.x2.X.n19 cdac_ctrl_0.x2.X 31.159
R10303 cdac_ctrl_0.x2.X.n20 cdac_ctrl_0.x2.X.n19 28.2061
R10304 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n20 27.5288
R10305 cdac_ctrl_0.x2.X.n0 cdac_ctrl_0.x2.X.t2 26.5955
R10306 cdac_ctrl_0.x2.X.n0 cdac_ctrl_0.x2.X.t8 26.5955
R10307 cdac_ctrl_0.x2.X.n29 cdac_ctrl_0.x2.X.t7 26.5955
R10308 cdac_ctrl_0.x2.X.n29 cdac_ctrl_0.x2.X.t15 26.5955
R10309 cdac_ctrl_0.x2.X.n28 cdac_ctrl_0.x2.X.t10 26.5955
R10310 cdac_ctrl_0.x2.X.n28 cdac_ctrl_0.x2.X.t3 26.5955
R10311 cdac_ctrl_0.x2.X.n30 cdac_ctrl_0.x2.X.t1 26.5955
R10312 cdac_ctrl_0.x2.X.n30 cdac_ctrl_0.x2.X.t5 26.5955
R10313 cdac_ctrl_0.x2.X.n21 cdac_ctrl_0.x2.X.t13 24.9236
R10314 cdac_ctrl_0.x2.X.n21 cdac_ctrl_0.x2.X.t12 24.9236
R10315 cdac_ctrl_0.x2.X.n22 cdac_ctrl_0.x2.X.t0 24.9236
R10316 cdac_ctrl_0.x2.X.n22 cdac_ctrl_0.x2.X.t14 24.9236
R10317 cdac_ctrl_0.x2.X.n23 cdac_ctrl_0.x2.X.t6 24.9236
R10318 cdac_ctrl_0.x2.X.n23 cdac_ctrl_0.x2.X.t4 24.9236
R10319 cdac_ctrl_0.x2.X.n26 cdac_ctrl_0.x2.X.t11 24.9236
R10320 cdac_ctrl_0.x2.X.n26 cdac_ctrl_0.x2.X.t9 24.9236
R10321 cdac_ctrl_0.x2.X.n33 cdac_ctrl_0.x2.X 12.8005
R10322 cdac_ctrl_0.x2.X.n5 cdac_ctrl_0.x2.X.n3 7.04781
R10323 cdac_ctrl_0.x2.X.n7 cdac_ctrl_0.x2.X.n5 7.04781
R10324 cdac_ctrl_0.x2.X.n9 cdac_ctrl_0.x2.X.n7 7.04781
R10325 cdac_ctrl_0.x2.X.n11 cdac_ctrl_0.x2.X.n9 7.04781
R10326 cdac_ctrl_0.x2.X.n13 cdac_ctrl_0.x2.X.n11 7.04781
R10327 cdac_ctrl_0.x2.X.n15 cdac_ctrl_0.x2.X.n13 7.04781
R10328 cdac_ctrl_0.x2.X.n17 cdac_ctrl_0.x2.X.n15 7.04781
R10329 cdac_ctrl_0.x2.X.n19 cdac_ctrl_0.x2.X.n17 7.04781
R10330 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n27 5.77305
R10331 cdac_ctrl_0.x2.X cdac_ctrl_0.x2.X.n33 4.26717
R10332 a_8520_n9662.n1 a_8520_n9662.n0 926.024
R10333 a_8520_n9662.t1 a_8520_n9662.n1 82.0838
R10334 a_8520_n9662.n0 a_8520_n9662.t0 63.3338
R10335 a_8520_n9662.n1 a_8520_n9662.t3 63.3219
R10336 a_8520_n9662.n0 a_8520_n9662.t2 29.7268
R10337 a_n784_n1599.n22 a_n784_n1599.t2 286.348
R10338 a_n784_n1599.n24 a_n784_n1599.t4 271.051
R10339 a_n784_n1599.n1 a_n784_n1599.t12 221.72
R10340 a_n784_n1599.n18 a_n784_n1599.t17 221.72
R10341 a_n784_n1599.n2 a_n784_n1599.t15 221.72
R10342 a_n784_n1599.n12 a_n784_n1599.t20 221.72
R10343 a_n784_n1599.n10 a_n784_n1599.t18 221.72
R10344 a_n784_n1599.n4 a_n784_n1599.t6 221.72
R10345 a_n784_n1599.n6 a_n784_n1599.t21 221.72
R10346 a_n784_n1599.n5 a_n784_n1599.t19 221.72
R10347 a_n784_n1599.n25 a_n784_n1599.n24 206.055
R10348 a_n784_n1599.n22 a_n784_n1599.n21 198.177
R10349 a_n784_n1599.n8 a_n784_n1599.n7 177.601
R10350 a_n784_n1599.n9 a_n784_n1599.n8 152
R10351 a_n784_n1599.n11 a_n784_n1599.n3 152
R10352 a_n784_n1599.n14 a_n784_n1599.n13 152
R10353 a_n784_n1599.n16 a_n784_n1599.n15 152
R10354 a_n784_n1599.n17 a_n784_n1599.n0 152
R10355 a_n784_n1599.n20 a_n784_n1599.n19 152
R10356 a_n784_n1599.n1 a_n784_n1599.t7 149.421
R10357 a_n784_n1599.n18 a_n784_n1599.t9 149.421
R10358 a_n784_n1599.n2 a_n784_n1599.t8 149.421
R10359 a_n784_n1599.n12 a_n784_n1599.t13 149.421
R10360 a_n784_n1599.n10 a_n784_n1599.t10 149.421
R10361 a_n784_n1599.n4 a_n784_n1599.t16 149.421
R10362 a_n784_n1599.n6 a_n784_n1599.t14 149.421
R10363 a_n784_n1599.n5 a_n784_n1599.t11 149.421
R10364 a_n784_n1599.n6 a_n784_n1599.n5 74.9783
R10365 a_n784_n1599.n7 a_n784_n1599.n6 66.0523
R10366 a_n784_n1599.n17 a_n784_n1599.n16 60.6968
R10367 a_n784_n1599.n19 a_n784_n1599.n18 55.3412
R10368 a_n784_n1599.n13 a_n784_n1599.n2 51.7709
R10369 a_n784_n1599.n9 a_n784_n1599.n4 51.7709
R10370 a_n784_n1599.n23 a_n784_n1599.n22 48.9632
R10371 a_n784_n1599.n24 a_n784_n1599.n23 38.7339
R10372 a_n784_n1599.n12 a_n784_n1599.n11 37.4894
R10373 a_n784_n1599.n11 a_n784_n1599.n10 37.4894
R10374 a_n784_n1599.n25 a_n784_n1599.t5 26.5955
R10375 a_n784_n1599.t0 a_n784_n1599.n25 26.5955
R10376 a_n784_n1599.n20 a_n784_n1599.n0 25.6005
R10377 a_n784_n1599.n15 a_n784_n1599.n0 25.6005
R10378 a_n784_n1599.n15 a_n784_n1599.n14 25.6005
R10379 a_n784_n1599.n14 a_n784_n1599.n3 25.6005
R10380 a_n784_n1599.n8 a_n784_n1599.n3 25.6005
R10381 a_n784_n1599.n21 a_n784_n1599.t1 24.9236
R10382 a_n784_n1599.n21 a_n784_n1599.t3 24.9236
R10383 a_n784_n1599.n13 a_n784_n1599.n12 23.2079
R10384 a_n784_n1599.n10 a_n784_n1599.n9 23.2079
R10385 a_n784_n1599.n19 a_n784_n1599.n1 19.6375
R10386 a_n784_n1599.n23 a_n784_n1599.n20 18.4476
R10387 a_n784_n1599.n16 a_n784_n1599.n2 8.92643
R10388 a_n784_n1599.n7 a_n784_n1599.n4 8.92643
R10389 a_n784_n1599.n18 a_n784_n1599.n17 5.35606
R10390 out_latch_0.FINAL.n18 out_latch_0.FINAL.n17 374.966
R10391 out_latch_0.FINAL out_latch_0.FINAL.n0 311.719
R10392 out_latch_0.FINAL.n18 out_latch_0.FINAL.n16 311.719
R10393 out_latch_0.FINAL.n20 out_latch_0.FINAL.n19 311.719
R10394 out_latch_0.FINAL.n4 out_latch_0.FINAL.n3 261.425
R10395 out_latch_0.FINAL.n8 out_latch_0.FINAL.t19 256.07
R10396 out_latch_0.FINAL.n10 out_latch_0.FINAL.t17 256.07
R10397 out_latch_0.FINAL.n7 out_latch_0.FINAL.n6 202.444
R10398 out_latch_0.FINAL.n4 out_latch_0.FINAL.n2 198.177
R10399 out_latch_0.FINAL.n5 out_latch_0.FINAL.n1 198.177
R10400 out_latch_0.FINAL.n9 out_latch_0.FINAL.n8 152
R10401 out_latch_0.FINAL.n11 out_latch_0.FINAL.n10 152
R10402 out_latch_0.FINAL.n8 out_latch_0.FINAL.t18 150.03
R10403 out_latch_0.FINAL.n10 out_latch_0.FINAL.t16 150.03
R10404 out_latch_0.FINAL.n14 out_latch_0.FINAL 94.1985
R10405 out_latch_0.FINAL.n5 out_latch_0.FINAL.n4 63.2476
R10406 out_latch_0.FINAL.n20 out_latch_0.FINAL.n18 63.2476
R10407 out_latch_0.FINAL.n7 out_latch_0.FINAL.n5 50.4476
R10408 out_latch_0.FINAL.n21 out_latch_0.FINAL.n20 50.4476
R10409 out_latch_0.FINAL out_latch_0.FINAL.n14 47.336
R10410 out_latch_0.FINAL.n13 out_latch_0.FINAL.n12 32.1552
R10411 out_latch_0.FINAL.n13 out_latch_0.FINAL 29.6287
R10412 out_latch_0.FINAL.n0 out_latch_0.FINAL.t8 26.5955
R10413 out_latch_0.FINAL.n0 out_latch_0.FINAL.t10 26.5955
R10414 out_latch_0.FINAL.n16 out_latch_0.FINAL.t13 26.5955
R10415 out_latch_0.FINAL.n16 out_latch_0.FINAL.t9 26.5955
R10416 out_latch_0.FINAL.n17 out_latch_0.FINAL.t14 26.5955
R10417 out_latch_0.FINAL.n17 out_latch_0.FINAL.t12 26.5955
R10418 out_latch_0.FINAL.n19 out_latch_0.FINAL.t11 26.5955
R10419 out_latch_0.FINAL.n19 out_latch_0.FINAL.t15 26.5955
R10420 out_latch_0.FINAL.n3 out_latch_0.FINAL.t7 24.9236
R10421 out_latch_0.FINAL.n3 out_latch_0.FINAL.t5 24.9236
R10422 out_latch_0.FINAL.n2 out_latch_0.FINAL.t6 24.9236
R10423 out_latch_0.FINAL.n2 out_latch_0.FINAL.t2 24.9236
R10424 out_latch_0.FINAL.n1 out_latch_0.FINAL.t4 24.9236
R10425 out_latch_0.FINAL.n1 out_latch_0.FINAL.t0 24.9236
R10426 out_latch_0.FINAL.n6 out_latch_0.FINAL.t1 24.9236
R10427 out_latch_0.FINAL.n6 out_latch_0.FINAL.t3 24.9236
R10428 out_latch_0.FINAL.n9 out_latch_0.FINAL 16.3845
R10429 out_latch_0.FINAL.n11 out_latch_0.FINAL 16.3845
R10430 out_latch_0.FINAL.n21 out_latch_0.FINAL.n15 11.0436
R10431 out_latch_0.FINAL out_latch_0.FINAL.n9 8.23114
R10432 out_latch_0.FINAL.n15 out_latch_0.FINAL 6.02403
R10433 out_latch_0.FINAL out_latch_0.FINAL.n7 5.77305
R10434 out_latch_0.FINAL.n14 out_latch_0.FINAL 4.69099
R10435 out_latch_0.FINAL.n12 out_latch_0.FINAL.n11 4.6085
R10436 out_latch_0.FINAL.n12 out_latch_0.FINAL 4.58918
R10437 out_latch_0.FINAL out_latch_0.FINAL.n21 4.26717
R10438 out_latch_0.FINAL.n15 out_latch_0.FINAL 2.00834
R10439 out_latch_0.FINAL out_latch_0.FINAL.n13 1.5005
R10440 a_8160_n5482.n1 a_8160_n5482.t3 530.01
R10441 a_8160_n5482.t1 a_8160_n5482.n5 421.021
R10442 a_8160_n5482.n0 a_8160_n5482.t6 337.171
R10443 a_8160_n5482.n3 a_8160_n5482.t0 280.223
R10444 a_8160_n5482.n4 a_8160_n5482.t7 263.173
R10445 a_8160_n5482.n4 a_8160_n5482.t2 227.826
R10446 a_8160_n5482.n0 a_8160_n5482.t5 199.762
R10447 a_8160_n5482.n2 a_8160_n5482.n1 170.81
R10448 a_8160_n5482.n2 a_8160_n5482.n0 167.321
R10449 a_8160_n5482.n5 a_8160_n5482.n4 152
R10450 a_8160_n5482.n1 a_8160_n5482.t4 141.923
R10451 a_8160_n5482.n3 a_8160_n5482.n2 10.8376
R10452 a_8160_n5482.n5 a_8160_n5482.n3 2.50485
R10453 a_8121_n5356.t1 a_8121_n5356.n3 370.026
R10454 a_8121_n5356.n0 a_8121_n5356.t3 351.356
R10455 a_8121_n5356.n1 a_8121_n5356.t5 334.717
R10456 a_8121_n5356.n3 a_8121_n5356.t0 325.971
R10457 a_8121_n5356.n1 a_8121_n5356.t4 309.935
R10458 a_8121_n5356.n0 a_8121_n5356.t2 305.683
R10459 a_8121_n5356.n2 a_8121_n5356.n0 16.879
R10460 a_8121_n5356.n3 a_8121_n5356.n2 10.8867
R10461 a_8121_n5356.n2 a_8121_n5356.n1 9.3005
R10462 CLK.n61 CLK.t11 294.557
R10463 CLK.n58 CLK.t28 294.557
R10464 CLK.n55 CLK.t39 294.557
R10465 CLK.n52 CLK.t41 294.557
R10466 CLK.n49 CLK.t24 294.557
R10467 CLK.n46 CLK.t20 294.557
R10468 CLK.n44 CLK.t38 294.557
R10469 CLK.n41 CLK.t33 294.557
R10470 CLK.n38 CLK.t37 294.557
R10471 CLK.n35 CLK.t23 294.557
R10472 CLK.n32 CLK.t16 294.557
R10473 CLK.n30 CLK.t32 294.557
R10474 CLK.n27 CLK.t13 294.557
R10475 CLK.n8 CLK.t25 294.557
R10476 CLK.n23 CLK.t0 294.557
R10477 CLK.n20 CLK.t2 294.557
R10478 CLK.n17 CLK.t19 294.557
R10479 CLK.n14 CLK.t8 294.557
R10480 CLK.n11 CLK.t12 294.557
R10481 CLK.n5 CLK.t3 294.557
R10482 CLK.n2 CLK.t27 294.557
R10483 CLK.n0 CLK.t10 294.557
R10484 CLK.n61 CLK.t9 211.01
R10485 CLK.n58 CLK.t31 211.01
R10486 CLK.n55 CLK.t43 211.01
R10487 CLK.n52 CLK.t1 211.01
R10488 CLK.n49 CLK.t26 211.01
R10489 CLK.n46 CLK.t22 211.01
R10490 CLK.n44 CLK.t42 211.01
R10491 CLK.n41 CLK.t30 211.01
R10492 CLK.n38 CLK.t36 211.01
R10493 CLK.n35 CLK.t21 211.01
R10494 CLK.n32 CLK.t15 211.01
R10495 CLK.n30 CLK.t29 211.01
R10496 CLK.n27 CLK.t18 211.01
R10497 CLK.n8 CLK.t4 211.01
R10498 CLK.n23 CLK.t34 211.01
R10499 CLK.n20 CLK.t40 211.01
R10500 CLK.n17 CLK.t14 211.01
R10501 CLK.n14 CLK.t5 211.01
R10502 CLK.n11 CLK.t7 211.01
R10503 CLK.n5 CLK.t6 211.01
R10504 CLK.n2 CLK.t35 211.01
R10505 CLK.n0 CLK.t17 211.01
R10506 CLK CLK.n23 156.207
R10507 CLK CLK.n20 156.207
R10508 CLK CLK.n17 156.207
R10509 CLK CLK.n14 156.207
R10510 CLK CLK.n11 156.207
R10511 CLK.n62 CLK.n61 152
R10512 CLK.n59 CLK.n58 152
R10513 CLK.n56 CLK.n55 152
R10514 CLK.n53 CLK.n52 152
R10515 CLK.n50 CLK.n49 152
R10516 CLK.n47 CLK.n46 152
R10517 CLK.n45 CLK.n44 152
R10518 CLK.n42 CLK.n41 152
R10519 CLK.n39 CLK.n38 152
R10520 CLK.n36 CLK.n35 152
R10521 CLK.n33 CLK.n32 152
R10522 CLK.n31 CLK.n30 152
R10523 CLK.n28 CLK.n27 152
R10524 CLK.n9 CLK.n8 152
R10525 CLK.n6 CLK.n5 152
R10526 CLK.n3 CLK.n2 152
R10527 CLK.n1 CLK.n0 152
R10528 CLK CLK.n65 42.0599
R10529 CLK.n65 CLK.n64 39.6039
R10530 CLK.n48 CLK 21.5434
R10531 CLK.n34 CLK 21.5194
R10532 CLK.n4 CLK 18.9565
R10533 CLK.n60 CLK 16.9379
R10534 CLK.n57 CLK 16.9379
R10535 CLK.n54 CLK 16.9379
R10536 CLK.n51 CLK 16.9379
R10537 CLK.n48 CLK 16.9379
R10538 CLK.n63 CLK 16.9139
R10539 CLK.n43 CLK 16.9139
R10540 CLK.n40 CLK 16.9139
R10541 CLK.n37 CLK 16.9139
R10542 CLK.n34 CLK 16.9139
R10543 CLK.n7 CLK 14.1662
R10544 CLK.n4 CLK 14.1662
R10545 CLK.n25 CLK.n24 13.889
R10546 CLK.n29 CLK 13.8005
R10547 CLK.n10 CLK 13.8005
R10548 CLK.n22 CLK.n21 13.8005
R10549 CLK.n19 CLK.n18 13.8005
R10550 CLK.n16 CLK.n15 13.8005
R10551 CLK.n13 CLK.n12 13.8005
R10552 CLK CLK.n62 10.4234
R10553 CLK CLK.n59 10.4234
R10554 CLK CLK.n56 10.4234
R10555 CLK CLK.n53 10.4234
R10556 CLK CLK.n50 10.4234
R10557 CLK CLK.n47 10.4234
R10558 CLK CLK.n45 10.4234
R10559 CLK CLK.n42 10.4234
R10560 CLK CLK.n39 10.4234
R10561 CLK CLK.n36 10.4234
R10562 CLK CLK.n33 10.4234
R10563 CLK CLK.n31 10.4234
R10564 CLK CLK.n28 10.4234
R10565 CLK CLK.n9 10.4234
R10566 CLK CLK.n6 10.4234
R10567 CLK CLK.n3 10.4234
R10568 CLK CLK.n1 10.4234
R10569 CLK.n63 CLK.n60 7.39156
R10570 CLK.n26 CLK.n25 7.26543
R10571 CLK.n24 CLK 6.58336
R10572 CLK.n21 CLK 6.58336
R10573 CLK.n18 CLK 6.58336
R10574 CLK.n15 CLK 6.21764
R10575 CLK.n15 CLK 6.21764
R10576 CLK.n12 CLK 6.21764
R10577 CLK.n12 CLK 6.21764
R10578 CLK.n24 CLK 5.85193
R10579 CLK.n21 CLK 5.85193
R10580 CLK.n18 CLK 5.85193
R10581 CLK.n10 CLK.n7 4.80266
R10582 CLK.n16 CLK.n13 4.79078
R10583 CLK.n19 CLK.n16 4.79078
R10584 CLK.n22 CLK.n19 4.79078
R10585 CLK.n7 CLK.n4 4.79078
R10586 CLK.n29 CLK.n26 4.69678
R10587 CLK.n25 CLK.n22 4.66022
R10588 CLK.n51 CLK.n48 4.606
R10589 CLK.n54 CLK.n51 4.606
R10590 CLK.n57 CLK.n54 4.606
R10591 CLK.n37 CLK.n34 4.606
R10592 CLK.n40 CLK.n37 4.606
R10593 CLK.n43 CLK.n40 4.606
R10594 CLK.n60 CLK.n57 4.58461
R10595 CLK.n63 CLK.n43 4.58461
R10596 CLK.n62 CLK 2.01193
R10597 CLK.n59 CLK 2.01193
R10598 CLK.n56 CLK 2.01193
R10599 CLK.n53 CLK 2.01193
R10600 CLK.n50 CLK 2.01193
R10601 CLK.n47 CLK 2.01193
R10602 CLK.n45 CLK 2.01193
R10603 CLK.n42 CLK 2.01193
R10604 CLK.n39 CLK 2.01193
R10605 CLK.n36 CLK 2.01193
R10606 CLK.n33 CLK 2.01193
R10607 CLK.n31 CLK 2.01193
R10608 CLK.n28 CLK 2.01193
R10609 CLK.n9 CLK 2.01193
R10610 CLK.n6 CLK 2.01193
R10611 CLK.n3 CLK 2.01193
R10612 CLK.n1 CLK 2.01193
R10613 CLK.n65 CLK 1.82675
R10614 CLK.n64 CLK.n63 1.13282
R10615 CLK.n13 CLK 0.415639
R10616 CLK CLK.n29 0.415639
R10617 CLK.n26 CLK.n10 0.0904123
R10618 CLK.n64 CLK 0.0413654
R10619 a_855_n1331.n1 a_855_n1331.t5 530.01
R10620 a_855_n1331.t1 a_855_n1331.n5 421.021
R10621 a_855_n1331.n0 a_855_n1331.t6 337.171
R10622 a_855_n1331.n3 a_855_n1331.t0 280.223
R10623 a_855_n1331.n4 a_855_n1331.t4 263.173
R10624 a_855_n1331.n4 a_855_n1331.t2 227.826
R10625 a_855_n1331.n0 a_855_n1331.t7 199.762
R10626 a_855_n1331.n2 a_855_n1331.n1 170.81
R10627 a_855_n1331.n2 a_855_n1331.n0 167.321
R10628 a_855_n1331.n5 a_855_n1331.n4 152
R10629 a_855_n1331.n1 a_855_n1331.t3 141.923
R10630 a_855_n1331.n3 a_855_n1331.n2 10.8376
R10631 a_855_n1331.n5 a_855_n1331.n3 2.50485
R10632 a_7274_2691.n3 a_7274_2691.n0 807.871
R10633 a_7274_2691.n4 a_7274_2691.t5 389.183
R10634 a_7274_2691.n5 a_7274_2691.n4 251.167
R10635 a_7274_2691.t0 a_7274_2691.n5 223.571
R10636 a_7274_2691.n1 a_7274_2691.t7 212.081
R10637 a_7274_2691.n2 a_7274_2691.t4 212.081
R10638 a_7274_2691.n3 a_7274_2691.n2 176.576
R10639 a_7274_2691.n4 a_7274_2691.t8 174.891
R10640 a_7274_2691.n1 a_7274_2691.t3 139.78
R10641 a_7274_2691.n2 a_7274_2691.t6 139.78
R10642 a_7274_2691.n0 a_7274_2691.t1 63.3219
R10643 a_7274_2691.n0 a_7274_2691.t2 63.3219
R10644 a_7274_2691.n2 a_7274_2691.n1 61.346
R10645 a_7274_2691.n5 a_7274_2691.n3 37.7195
R10646 auto_sampling_0.x21.D.n5 auto_sampling_0.x21.D.n4 585
R10647 auto_sampling_0.x21.D.n4 auto_sampling_0.x21.D.n3 585
R10648 auto_sampling_0.x21.D.n2 auto_sampling_0.x21.D.t4 333.651
R10649 auto_sampling_0.x21.D.n2 auto_sampling_0.x21.D.t5 297.233
R10650 auto_sampling_0.x21.D auto_sampling_0.x21.D.n2 196.493
R10651 auto_sampling_0.x21.D.n1 auto_sampling_0.x21.D.n0 185
R10652 auto_sampling_0.x21.D auto_sampling_0.x21.D.n1 49.0339
R10653 auto_sampling_0.x21.D.n3 auto_sampling_0.x21.D 44.2533
R10654 auto_sampling_0.x21.D.n4 auto_sampling_0.x21.D.t2 26.5955
R10655 auto_sampling_0.x21.D.n4 auto_sampling_0.x21.D.t3 26.5955
R10656 auto_sampling_0.x21.D.n0 auto_sampling_0.x21.D.t1 24.9236
R10657 auto_sampling_0.x21.D.n0 auto_sampling_0.x21.D.t0 24.9236
R10658 auto_sampling_0.x21.D.n5 auto_sampling_0.x21.D 15.6165
R10659 auto_sampling_0.x21.D.n1 auto_sampling_0.x21.D 10.4965
R10660 auto_sampling_0.x21.D.n3 auto_sampling_0.x21.D 1.7925
R10661 auto_sampling_0.x21.D auto_sampling_0.x21.D.n5 1.7925
R10662 a_n10393_n10028.n22 a_n10393_n10028.t2 286.348
R10663 a_n10393_n10028.n24 a_n10393_n10028.t4 271.051
R10664 a_n10393_n10028.n4 a_n10393_n10028.t8 221.72
R10665 a_n10393_n10028.n5 a_n10393_n10028.t14 221.72
R10666 a_n10393_n10028.n3 a_n10393_n10028.t16 221.72
R10667 a_n10393_n10028.n9 a_n10393_n10028.t9 221.72
R10668 a_n10393_n10028.n11 a_n10393_n10028.t13 221.72
R10669 a_n10393_n10028.n1 a_n10393_n10028.t21 221.72
R10670 a_n10393_n10028.n17 a_n10393_n10028.t7 221.72
R10671 a_n10393_n10028.n18 a_n10393_n10028.t11 221.72
R10672 a_n10393_n10028.n25 a_n10393_n10028.n24 206.055
R10673 a_n10393_n10028.n22 a_n10393_n10028.n21 198.177
R10674 a_n10393_n10028.n7 a_n10393_n10028.n6 177.601
R10675 a_n10393_n10028.n20 a_n10393_n10028.n19 152
R10676 a_n10393_n10028.n16 a_n10393_n10028.n0 152
R10677 a_n10393_n10028.n15 a_n10393_n10028.n14 152
R10678 a_n10393_n10028.n13 a_n10393_n10028.n12 152
R10679 a_n10393_n10028.n10 a_n10393_n10028.n2 152
R10680 a_n10393_n10028.n8 a_n10393_n10028.n7 152
R10681 a_n10393_n10028.n4 a_n10393_n10028.t17 149.421
R10682 a_n10393_n10028.n5 a_n10393_n10028.t15 149.421
R10683 a_n10393_n10028.n3 a_n10393_n10028.t19 149.421
R10684 a_n10393_n10028.n9 a_n10393_n10028.t18 149.421
R10685 a_n10393_n10028.n11 a_n10393_n10028.t6 149.421
R10686 a_n10393_n10028.n1 a_n10393_n10028.t20 149.421
R10687 a_n10393_n10028.n17 a_n10393_n10028.t12 149.421
R10688 a_n10393_n10028.n18 a_n10393_n10028.t10 149.421
R10689 a_n10393_n10028.n5 a_n10393_n10028.n4 74.9783
R10690 a_n10393_n10028.n6 a_n10393_n10028.n5 66.0523
R10691 a_n10393_n10028.n16 a_n10393_n10028.n15 60.6968
R10692 a_n10393_n10028.n19 a_n10393_n10028.n17 55.3412
R10693 a_n10393_n10028.n8 a_n10393_n10028.n3 51.7709
R10694 a_n10393_n10028.n12 a_n10393_n10028.n1 51.7709
R10695 a_n10393_n10028.n23 a_n10393_n10028.n22 48.9632
R10696 a_n10393_n10028.n24 a_n10393_n10028.n23 38.7339
R10697 a_n10393_n10028.n10 a_n10393_n10028.n9 37.4894
R10698 a_n10393_n10028.n11 a_n10393_n10028.n10 37.4894
R10699 a_n10393_n10028.n25 a_n10393_n10028.t5 26.5955
R10700 a_n10393_n10028.t0 a_n10393_n10028.n25 26.5955
R10701 a_n10393_n10028.n7 a_n10393_n10028.n2 25.6005
R10702 a_n10393_n10028.n13 a_n10393_n10028.n2 25.6005
R10703 a_n10393_n10028.n14 a_n10393_n10028.n13 25.6005
R10704 a_n10393_n10028.n14 a_n10393_n10028.n0 25.6005
R10705 a_n10393_n10028.n20 a_n10393_n10028.n0 25.6005
R10706 a_n10393_n10028.n21 a_n10393_n10028.t1 24.9236
R10707 a_n10393_n10028.n21 a_n10393_n10028.t3 24.9236
R10708 a_n10393_n10028.n9 a_n10393_n10028.n8 23.2079
R10709 a_n10393_n10028.n12 a_n10393_n10028.n11 23.2079
R10710 a_n10393_n10028.n19 a_n10393_n10028.n18 19.6375
R10711 a_n10393_n10028.n23 a_n10393_n10028.n20 18.4476
R10712 a_n10393_n10028.n6 a_n10393_n10028.n3 8.92643
R10713 a_n10393_n10028.n15 a_n10393_n10028.n1 8.92643
R10714 a_n10393_n10028.n17 a_n10393_n10028.n16 5.35606
R10715 a_6333_n9484.t0 a_6333_n9484.n3 370.026
R10716 a_6333_n9484.n0 a_6333_n9484.t4 351.356
R10717 a_6333_n9484.n1 a_6333_n9484.t2 334.717
R10718 a_6333_n9484.n3 a_6333_n9484.t1 325.971
R10719 a_6333_n9484.n1 a_6333_n9484.t5 309.935
R10720 a_6333_n9484.n0 a_6333_n9484.t3 305.683
R10721 a_6333_n9484.n2 a_6333_n9484.n0 16.879
R10722 a_6333_n9484.n3 a_6333_n9484.n2 10.8867
R10723 a_6333_n9484.n2 a_6333_n9484.n1 9.3005
R10724 a_6683_n9484.n3 a_6683_n9484.n2 674.338
R10725 a_6683_n9484.n1 a_6683_n9484.t5 332.58
R10726 a_6683_n9484.n2 a_6683_n9484.n0 284.012
R10727 a_6683_n9484.n2 a_6683_n9484.n1 253.648
R10728 a_6683_n9484.n1 a_6683_n9484.t4 168.701
R10729 a_6683_n9484.n3 a_6683_n9484.t3 96.1553
R10730 a_6683_n9484.t0 a_6683_n9484.n3 65.6672
R10731 a_6683_n9484.n0 a_6683_n9484.t2 65.0005
R10732 a_6683_n9484.n0 a_6683_n9484.t1 45.0005
R10733 a_6779_n9484.t0 a_6779_n9484.t1 198.571
R10734 a_n8773_n9484.n3 a_n8773_n9484.n2 674.338
R10735 a_n8773_n9484.n1 a_n8773_n9484.t4 332.58
R10736 a_n8773_n9484.n2 a_n8773_n9484.n0 284.012
R10737 a_n8773_n9484.n2 a_n8773_n9484.n1 253.648
R10738 a_n8773_n9484.n1 a_n8773_n9484.t5 168.701
R10739 a_n8773_n9484.n3 a_n8773_n9484.t3 96.1553
R10740 a_n8773_n9484.t1 a_n8773_n9484.n3 65.6672
R10741 a_n8773_n9484.n0 a_n8773_n9484.t0 65.0005
R10742 a_n8773_n9484.n0 a_n8773_n9484.t2 45.0005
R10743 a_n8555_n9242.n3 a_n8555_n9242.n2 647.119
R10744 a_n8555_n9242.n1 a_n8555_n9242.t5 350.253
R10745 a_n8555_n9242.n2 a_n8555_n9242.n0 260.339
R10746 a_n8555_n9242.n2 a_n8555_n9242.n1 246.119
R10747 a_n8555_n9242.n1 a_n8555_n9242.t4 189.588
R10748 a_n8555_n9242.n3 a_n8555_n9242.t0 89.1195
R10749 a_n8555_n9242.n0 a_n8555_n9242.t1 63.3338
R10750 a_n8555_n9242.t3 a_n8555_n9242.n3 41.0422
R10751 a_n8555_n9242.n0 a_n8555_n9242.t2 31.9797
R10752 a_4452_n5387.n3 a_4452_n5387.n2 674.338
R10753 a_4452_n5387.n1 a_4452_n5387.t4 332.58
R10754 a_4452_n5387.n2 a_4452_n5387.n0 284.012
R10755 a_4452_n5387.n2 a_4452_n5387.n1 253.648
R10756 a_4452_n5387.n1 a_4452_n5387.t5 168.701
R10757 a_4452_n5387.n3 a_4452_n5387.t3 96.1553
R10758 a_4452_n5387.t1 a_4452_n5387.n3 65.6672
R10759 a_4452_n5387.n0 a_4452_n5387.t2 65.0005
R10760 a_4452_n5387.n0 a_4452_n5387.t0 45.0005
R10761 a_4383_n5258.n3 a_4383_n5258.n2 647.119
R10762 a_4383_n5258.n1 a_4383_n5258.t4 350.253
R10763 a_4383_n5258.n2 a_4383_n5258.n0 260.339
R10764 a_4383_n5258.n2 a_4383_n5258.n1 246.119
R10765 a_4383_n5258.n1 a_4383_n5258.t5 189.588
R10766 a_4383_n5258.n3 a_4383_n5258.t3 89.1195
R10767 a_4383_n5258.n0 a_4383_n5258.t0 63.3338
R10768 a_4383_n5258.t2 a_4383_n5258.n3 41.0422
R10769 a_4383_n5258.n0 a_4383_n5258.t1 31.9797
R10770 a_2451_n5258.n3 a_2451_n5258.n2 647.119
R10771 a_2451_n5258.n1 a_2451_n5258.t4 350.253
R10772 a_2451_n5258.n2 a_2451_n5258.n0 260.339
R10773 a_2451_n5258.n2 a_2451_n5258.n1 246.119
R10774 a_2451_n5258.n1 a_2451_n5258.t5 189.588
R10775 a_2451_n5258.n3 a_2451_n5258.t1 89.1195
R10776 a_2451_n5258.n0 a_2451_n5258.t3 63.3338
R10777 a_2451_n5258.t0 a_2451_n5258.n3 41.0422
R10778 a_2451_n5258.n0 a_2451_n5258.t2 31.9797
R10779 a_2758_n5624.t0 a_2758_n5624.t1 60.0005
R10780 a_2830_n5624.t0 a_2830_n5624.t1 198.571
R10781 a_4713_n4702.n3 a_4713_n4702.n2 636.953
R10782 a_4713_n4702.n1 a_4713_n4702.t5 366.856
R10783 a_4713_n4702.n2 a_4713_n4702.n0 300.2
R10784 a_4713_n4702.n2 a_4713_n4702.n1 225.036
R10785 a_4713_n4702.n1 a_4713_n4702.t4 174.056
R10786 a_4713_n4702.n0 a_4713_n4702.t3 70.0005
R10787 a_4713_n4702.t1 a_4713_n4702.n3 68.0124
R10788 a_4713_n4702.n3 a_4713_n4702.t2 63.3219
R10789 a_4713_n4702.n0 a_4713_n4702.t0 61.6672
R10790 a_4888_n4776.n5 a_4888_n4776.n4 807.871
R10791 a_4888_n4776.n2 a_4888_n4776.t8 389.183
R10792 a_4888_n4776.n3 a_4888_n4776.n2 251.167
R10793 a_4888_n4776.n3 a_4888_n4776.t2 223.571
R10794 a_4888_n4776.n0 a_4888_n4776.t3 212.081
R10795 a_4888_n4776.n1 a_4888_n4776.t4 212.081
R10796 a_4888_n4776.n4 a_4888_n4776.n1 176.576
R10797 a_4888_n4776.n2 a_4888_n4776.t5 174.891
R10798 a_4888_n4776.n0 a_4888_n4776.t6 139.78
R10799 a_4888_n4776.n1 a_4888_n4776.t7 139.78
R10800 a_4888_n4776.n5 a_4888_n4776.t1 63.3219
R10801 a_4888_n4776.t0 a_4888_n4776.n5 63.3219
R10802 a_4888_n4776.n1 a_4888_n4776.n0 61.346
R10803 a_4888_n4776.n4 a_4888_n4776.n3 37.7195
R10804 a_n1395_n10022.t0 a_n1395_n10022.n3 370.026
R10805 a_n1395_n10022.n0 a_n1395_n10022.t2 351.356
R10806 a_n1395_n10022.n1 a_n1395_n10022.t3 334.717
R10807 a_n1395_n10022.n3 a_n1395_n10022.t1 325.971
R10808 a_n1395_n10022.n1 a_n1395_n10022.t5 309.935
R10809 a_n1395_n10022.n0 a_n1395_n10022.t4 305.683
R10810 a_n1395_n10022.n2 a_n1395_n10022.n0 16.879
R10811 a_n1395_n10022.n3 a_n1395_n10022.n2 10.8867
R10812 a_n1395_n10022.n2 a_n1395_n10022.n1 9.3005
R10813 a_n827_n10054.n3 a_n827_n10054.n2 647.119
R10814 a_n827_n10054.n1 a_n827_n10054.t4 350.253
R10815 a_n827_n10054.n2 a_n827_n10054.n0 260.339
R10816 a_n827_n10054.n2 a_n827_n10054.n1 246.119
R10817 a_n827_n10054.n1 a_n827_n10054.t5 189.588
R10818 a_n827_n10054.n3 a_n827_n10054.t1 89.1195
R10819 a_n827_n10054.n0 a_n827_n10054.t0 63.3338
R10820 a_n827_n10054.t2 a_n827_n10054.n3 41.0422
R10821 a_n827_n10054.n0 a_n827_n10054.t3 31.9797
R10822 a_n480_n9650.n3 a_n480_n9650.n2 636.953
R10823 a_n480_n9650.n1 a_n480_n9650.t4 366.856
R10824 a_n480_n9650.n2 a_n480_n9650.n0 300.2
R10825 a_n480_n9650.n2 a_n480_n9650.n1 225.036
R10826 a_n480_n9650.n1 a_n480_n9650.t5 174.056
R10827 a_n480_n9650.n0 a_n480_n9650.t0 70.0005
R10828 a_n480_n9650.n3 a_n480_n9650.t2 68.0124
R10829 a_n480_n9650.t1 a_n480_n9650.n3 63.3219
R10830 a_n480_n9650.n0 a_n480_n9650.t3 61.6672
R10831 a_n172_n5650.n3 a_n172_n5650.n0 807.871
R10832 a_n172_n5650.n4 a_n172_n5650.t6 389.183
R10833 a_n172_n5650.n5 a_n172_n5650.n4 251.167
R10834 a_n172_n5650.t0 a_n172_n5650.n5 223.571
R10835 a_n172_n5650.n2 a_n172_n5650.t7 212.081
R10836 a_n172_n5650.n1 a_n172_n5650.t3 212.081
R10837 a_n172_n5650.n3 a_n172_n5650.n2 176.576
R10838 a_n172_n5650.n4 a_n172_n5650.t5 174.891
R10839 a_n172_n5650.n2 a_n172_n5650.t4 139.78
R10840 a_n172_n5650.n1 a_n172_n5650.t8 139.78
R10841 a_n172_n5650.n0 a_n172_n5650.t2 63.3219
R10842 a_n172_n5650.n0 a_n172_n5650.t1 63.3219
R10843 a_n172_n5650.n2 a_n172_n5650.n1 61.346
R10844 a_n172_n5650.n5 a_n172_n5650.n3 37.5061
R10845 DOUT[0].n3 DOUT[0].n2 585
R10846 DOUT[0].n4 DOUT[0].n3 585
R10847 DOUT[0].n1 DOUT[0].n0 185
R10848 DOUT[0] DOUT[0].n1 49.0339
R10849 DOUT[0].n3 DOUT[0].t2 26.5955
R10850 DOUT[0].n3 DOUT[0].t3 26.5955
R10851 DOUT[0].n0 DOUT[0].t1 24.9236
R10852 DOUT[0].n0 DOUT[0].t0 24.9236
R10853 DOUT[0].n5 DOUT[0] 23.8854
R10854 DOUT[0].n5 DOUT[0].n4 20.576
R10855 DOUT[0].n2 DOUT[0] 15.6165
R10856 DOUT[0].n1 DOUT[0] 10.4965
R10857 DOUT[0].n4 DOUT[0] 1.7925
R10858 DOUT[0].n2 DOUT[0] 1.7925
R10859 DOUT[0] DOUT[0].n5 0.00285
R10860 a_n454_2691.n5 a_n454_2691.n4 807.871
R10861 a_n454_2691.n2 a_n454_2691.t4 389.183
R10862 a_n454_2691.n3 a_n454_2691.n2 251.167
R10863 a_n454_2691.n3 a_n454_2691.t2 223.571
R10864 a_n454_2691.n0 a_n454_2691.t7 212.081
R10865 a_n454_2691.n1 a_n454_2691.t6 212.081
R10866 a_n454_2691.n4 a_n454_2691.n1 176.576
R10867 a_n454_2691.n2 a_n454_2691.t5 174.891
R10868 a_n454_2691.n0 a_n454_2691.t3 139.78
R10869 a_n454_2691.n1 a_n454_2691.t8 139.78
R10870 a_n454_2691.n5 a_n454_2691.t1 63.3219
R10871 a_n454_2691.t0 a_n454_2691.n5 63.3219
R10872 a_n454_2691.n1 a_n454_2691.n0 61.346
R10873 a_n454_2691.n4 a_n454_2691.n3 37.7195
R10874 auto_sampling_0.x22.A.n9 auto_sampling_0.x22.A.n8 585
R10875 auto_sampling_0.x22.A.n8 auto_sampling_0.x22.A.n7 585
R10876 auto_sampling_0.x22.A.n2 auto_sampling_0.x22.A.t9 333.651
R10877 auto_sampling_0.x22.A.n2 auto_sampling_0.x22.A.t6 297.233
R10878 auto_sampling_0.x22.A.n3 auto_sampling_0.x22.A.t5 212.081
R10879 auto_sampling_0.x22.A.n4 auto_sampling_0.x22.A.t7 212.081
R10880 auto_sampling_0.x22.A auto_sampling_0.x22.A.n2 196.493
R10881 auto_sampling_0.x22.A.n1 auto_sampling_0.x22.A.n0 185
R10882 auto_sampling_0.x22.A.n5 auto_sampling_0.x22.A.n4 184.721
R10883 auto_sampling_0.x22.A.n3 auto_sampling_0.x22.A.t8 139.78
R10884 auto_sampling_0.x22.A.n4 auto_sampling_0.x22.A.t4 139.78
R10885 auto_sampling_0.x22.A.n4 auto_sampling_0.x22.A.n3 61.346
R10886 auto_sampling_0.x22.A auto_sampling_0.x22.A.n1 49.0339
R10887 auto_sampling_0.x22.A.n6 auto_sampling_0.x22.A 32.3715
R10888 auto_sampling_0.x22.A.n6 auto_sampling_0.x22.A.n5 27.2303
R10889 auto_sampling_0.x22.A.n8 auto_sampling_0.x22.A.t2 26.5955
R10890 auto_sampling_0.x22.A.n8 auto_sampling_0.x22.A.t3 26.5955
R10891 auto_sampling_0.x22.A.n0 auto_sampling_0.x22.A.t1 24.9236
R10892 auto_sampling_0.x22.A.n0 auto_sampling_0.x22.A.t0 24.9236
R10893 auto_sampling_0.x22.A.n9 auto_sampling_0.x22.A 15.6165
R10894 auto_sampling_0.x22.A.n7 auto_sampling_0.x22.A.n6 11.8605
R10895 auto_sampling_0.x22.A.n1 auto_sampling_0.x22.A 10.4965
R10896 auto_sampling_0.x22.A.n5 auto_sampling_0.x22.A 4.3525
R10897 auto_sampling_0.x22.A.n7 auto_sampling_0.x22.A 1.7925
R10898 auto_sampling_0.x22.A auto_sampling_0.x22.A.n9 1.7925
R10899 a_n66_n5074.t1 a_n66_n5074.n3 370.026
R10900 a_n66_n5074.n0 a_n66_n5074.t5 351.356
R10901 a_n66_n5074.n1 a_n66_n5074.t3 334.717
R10902 a_n66_n5074.n3 a_n66_n5074.t0 325.971
R10903 a_n66_n5074.n1 a_n66_n5074.t4 309.935
R10904 a_n66_n5074.n0 a_n66_n5074.t2 305.683
R10905 a_n66_n5074.n2 a_n66_n5074.n0 16.879
R10906 a_n66_n5074.n3 a_n66_n5074.n2 10.8867
R10907 a_n66_n5074.n2 a_n66_n5074.n1 9.3005
R10908 a_849_n4702.n3 a_849_n4702.n2 636.953
R10909 a_849_n4702.n1 a_849_n4702.t5 366.856
R10910 a_849_n4702.n2 a_849_n4702.n0 300.2
R10911 a_849_n4702.n2 a_849_n4702.n1 225.036
R10912 a_849_n4702.n1 a_849_n4702.t4 174.056
R10913 a_849_n4702.n0 a_849_n4702.t1 70.0005
R10914 a_849_n4702.n3 a_849_n4702.t2 68.0124
R10915 a_849_n4702.t0 a_849_n4702.n3 63.3219
R10916 a_849_n4702.n0 a_849_n4702.t3 61.6672
R10917 a_1011_n5080.t0 a_1011_n5080.t1 126.644
R10918 a_371_n9484.n1 a_371_n9484.t2 530.01
R10919 a_371_n9484.t0 a_371_n9484.n5 421.021
R10920 a_371_n9484.n0 a_371_n9484.t5 337.142
R10921 a_371_n9484.n3 a_371_n9484.t1 280.223
R10922 a_371_n9484.n4 a_371_n9484.t4 263.173
R10923 a_371_n9484.n4 a_371_n9484.t7 227.826
R10924 a_371_n9484.n0 a_371_n9484.t6 199.762
R10925 a_371_n9484.n2 a_371_n9484.n1 170.81
R10926 a_371_n9484.n2 a_371_n9484.n0 167.321
R10927 a_371_n9484.n5 a_371_n9484.n4 152
R10928 a_371_n9484.n1 a_371_n9484.t3 141.923
R10929 a_371_n9484.n3 a_371_n9484.n2 10.8376
R10930 a_371_n9484.n5 a_371_n9484.n3 2.50485
R10931 a_887_n9484.n3 a_887_n9484.n2 674.338
R10932 a_887_n9484.n1 a_887_n9484.t4 332.58
R10933 a_887_n9484.n2 a_887_n9484.n0 284.012
R10934 a_887_n9484.n2 a_887_n9484.n1 253.648
R10935 a_887_n9484.n1 a_887_n9484.t5 168.701
R10936 a_887_n9484.t0 a_887_n9484.n3 96.1553
R10937 a_887_n9484.n3 a_887_n9484.t2 65.6672
R10938 a_887_n9484.n0 a_887_n9484.t1 65.0005
R10939 a_887_n9484.n0 a_887_n9484.t3 45.0005
R10940 a_995_n9118.n0 a_995_n9118.t1 1327.82
R10941 a_995_n9118.t0 a_995_n9118.n0 194.655
R10942 a_995_n9118.n0 a_995_n9118.t2 63.3219
R10943 a_n1543_3557.t1 a_n1543_3557.n3 370.026
R10944 a_n1543_3557.n0 a_n1543_3557.t4 351.356
R10945 a_n1543_3557.n1 a_n1543_3557.t3 334.717
R10946 a_n1543_3557.n3 a_n1543_3557.t0 325.971
R10947 a_n1543_3557.n1 a_n1543_3557.t2 309.935
R10948 a_n1543_3557.n0 a_n1543_3557.t5 305.683
R10949 a_n1543_3557.n2 a_n1543_3557.n0 16.879
R10950 a_n1543_3557.n3 a_n1543_3557.n2 10.8867
R10951 a_n1543_3557.n2 a_n1543_3557.n1 9.3005
R10952 a_n1288_3557.n1 a_n1288_3557.n0 926.024
R10953 a_n1288_3557.t0 a_n1288_3557.n1 82.0838
R10954 a_n1288_3557.n0 a_n1288_3557.t1 63.3338
R10955 a_n1288_3557.n1 a_n1288_3557.t3 63.3219
R10956 a_n1288_3557.n0 a_n1288_3557.t2 29.7268
R10957 a_n305_n9510.n5 a_n305_n9510.n4 807.871
R10958 a_n305_n9510.n2 a_n305_n9510.t4 389.183
R10959 a_n305_n9510.n3 a_n305_n9510.n2 251.167
R10960 a_n305_n9510.n3 a_n305_n9510.t1 223.571
R10961 a_n305_n9510.n0 a_n305_n9510.t8 212.081
R10962 a_n305_n9510.n1 a_n305_n9510.t6 212.081
R10963 a_n305_n9510.n4 a_n305_n9510.n1 176.576
R10964 a_n305_n9510.n2 a_n305_n9510.t3 174.891
R10965 a_n305_n9510.n0 a_n305_n9510.t7 139.78
R10966 a_n305_n9510.n1 a_n305_n9510.t5 139.78
R10967 a_n305_n9510.t0 a_n305_n9510.n5 63.3219
R10968 a_n305_n9510.n5 a_n305_n9510.t2 63.3219
R10969 a_n305_n9510.n1 a_n305_n9510.n0 61.346
R10970 a_n305_n9510.n4 a_n305_n9510.n3 37.7195
R10971 a_n371_n9484.t1 a_n371_n9484.t0 94.7268
R10972 a_n2869_n10028.n0 a_n2869_n10028.t2 1327.82
R10973 a_n2869_n10028.t0 a_n2869_n10028.n0 194.655
R10974 a_n2869_n10028.n0 a_n2869_n10028.t1 63.3219
R10975 a_n8665_n9118.n0 a_n8665_n9118.t2 1327.82
R10976 a_n8665_n9118.t0 a_n8665_n9118.n0 194.655
R10977 a_n8665_n9118.n0 a_n8665_n9118.t1 63.3219
R10978 a_1626_n1029.t0 a_1626_n1029.t1 87.1434
R10979 a_2320_2717.t1 a_2320_2717.n3 370.026
R10980 a_2320_2717.n0 a_2320_2717.t3 351.356
R10981 a_2320_2717.n1 a_2320_2717.t5 334.717
R10982 a_2320_2717.n3 a_2320_2717.t0 325.971
R10983 a_2320_2717.n1 a_2320_2717.t4 309.935
R10984 a_2320_2717.n0 a_2320_2717.t2 305.683
R10985 a_2320_2717.n2 a_2320_2717.n0 16.879
R10986 a_2320_2717.n3 a_2320_2717.n2 10.8867
R10987 a_2320_2717.n2 a_2320_2717.n1 9.3005
R10988 a_3235_2717.n3 a_3235_2717.n2 636.953
R10989 a_3235_2717.n1 a_3235_2717.t4 366.856
R10990 a_3235_2717.n2 a_3235_2717.n0 300.2
R10991 a_3235_2717.n2 a_3235_2717.n1 225.036
R10992 a_3235_2717.n1 a_3235_2717.t5 174.056
R10993 a_3235_2717.n0 a_3235_2717.t0 70.0005
R10994 a_3235_2717.n3 a_3235_2717.t3 68.0124
R10995 a_3235_2717.t1 a_3235_2717.n3 63.3219
R10996 a_3235_2717.n0 a_3235_2717.t2 61.6672
R10997 a_3397_3083.t0 a_3397_3083.t1 126.644
R10998 EN.n208 EN.t78 408.63
R10999 EN.n197 EN.t23 408.63
R11000 EN.n186 EN.t56 408.63
R11001 EN.n175 EN.t88 408.63
R11002 EN.n164 EN.t58 408.63
R11003 EN.n153 EN.t51 408.63
R11004 EN.n103 EN.t35 408.63
R11005 EN.n146 EN.t65 408.63
R11006 EN.n137 EN.t75 408.63
R11007 EN.n128 EN.t38 408.63
R11008 EN.n119 EN.t4 408.63
R11009 EN.n111 EN.t10 408.63
R11010 EN.n89 EN.t72 408.63
R11011 EN.n79 EN.t46 408.63
R11012 EN.n48 EN.t31 408.63
R11013 EN.n57 EN.t29 408.63
R11014 EN.n67 EN.t0 408.63
R11015 EN.n38 EN.t48 408.63
R11016 EN.n29 EN.t52 408.63
R11017 EN.n19 EN.t17 408.63
R11018 EN.n9 EN.t86 408.63
R11019 EN.n0 EN.t89 408.63
R11020 EN.n211 EN.t11 347.577
R11021 EN.n200 EN.t62 347.577
R11022 EN.n189 EN.t32 347.577
R11023 EN.n178 EN.t20 347.577
R11024 EN.n167 EN.t59 347.577
R11025 EN.n156 EN.t26 347.577
R11026 EN.n100 EN.t7 347.577
R11027 EN.n143 EN.t43 347.577
R11028 EN.n134 EN.t2 347.577
R11029 EN.n125 EN.t39 347.577
R11030 EN.n116 EN.t47 347.577
R11031 EN.n108 EN.t44 347.577
R11032 EN.n92 EN.t28 347.577
R11033 EN.n82 EN.t36 347.577
R11034 EN.n51 EN.t63 347.577
R11035 EN.n60 EN.t30 347.577
R11036 EN.n70 EN.t1 347.577
R11037 EN.n41 EN.t6 347.577
R11038 EN.n32 EN.t87 347.577
R11039 EN.n22 EN.t5 347.577
R11040 EN.n12 EN.t84 347.577
R11041 EN.n3 EN.t69 347.577
R11042 EN.n220 EN.t54 333.651
R11043 EN.n220 EN.t64 297.233
R11044 EN.n221 EN.n220 196.493
R11045 EN.n211 EN.t61 193.337
R11046 EN.n200 EN.t16 193.337
R11047 EN.n189 EN.t81 193.337
R11048 EN.n178 EN.t73 193.337
R11049 EN.n167 EN.t14 193.337
R11050 EN.n156 EN.t79 193.337
R11051 EN.n100 EN.t85 193.337
R11052 EN.n143 EN.t22 193.337
R11053 EN.n134 EN.t82 193.337
R11054 EN.n125 EN.t18 193.337
R11055 EN.n116 EN.t27 193.337
R11056 EN.n108 EN.t24 193.337
R11057 EN.n92 EN.t9 193.337
R11058 EN.n82 EN.t15 193.337
R11059 EN.n51 EN.t12 193.337
R11060 EN.n60 EN.t76 193.337
R11061 EN.n70 EN.t49 193.337
R11062 EN.n41 EN.t55 193.337
R11063 EN.n32 EN.t40 193.337
R11064 EN.n22 EN.t83 193.337
R11065 EN.n12 EN.t70 193.337
R11066 EN.n3 EN.t50 193.337
R11067 EN EN.n48 165.201
R11068 EN EN.n57 165.201
R11069 EN EN.n67 165.201
R11070 EN EN.n38 165.201
R11071 EN EN.n29 165.201
R11072 EN.n209 EN.n208 165.072
R11073 EN.n198 EN.n197 165.072
R11074 EN.n187 EN.n186 165.072
R11075 EN.n176 EN.n175 165.072
R11076 EN.n165 EN.n164 165.072
R11077 EN.n154 EN.n153 165.072
R11078 EN.n104 EN.n103 165.072
R11079 EN.n147 EN.n146 165.072
R11080 EN.n138 EN.n137 165.072
R11081 EN.n129 EN.n128 165.072
R11082 EN.n120 EN.n119 165.072
R11083 EN.n112 EN.n111 165.072
R11084 EN.n90 EN.n89 165.072
R11085 EN.n80 EN.n79 165.072
R11086 EN.n20 EN.n19 165.072
R11087 EN.n10 EN.n9 165.072
R11088 EN.n1 EN.n0 165.072
R11089 EN.n212 EN.n211 152
R11090 EN.n201 EN.n200 152
R11091 EN.n190 EN.n189 152
R11092 EN.n179 EN.n178 152
R11093 EN.n168 EN.n167 152
R11094 EN.n157 EN.n156 152
R11095 EN.n101 EN.n100 152
R11096 EN.n144 EN.n143 152
R11097 EN.n135 EN.n134 152
R11098 EN.n126 EN.n125 152
R11099 EN.n117 EN.n116 152
R11100 EN.n109 EN.n108 152
R11101 EN.n93 EN.n92 152
R11102 EN.n83 EN.n82 152
R11103 EN.n52 EN.n51 152
R11104 EN.n61 EN.n60 152
R11105 EN.n71 EN.n70 152
R11106 EN.n42 EN.n41 152
R11107 EN.n33 EN.n32 152
R11108 EN.n23 EN.n22 152
R11109 EN.n13 EN.n12 152
R11110 EN.n4 EN.n3 152
R11111 EN.n208 EN.t74 132.282
R11112 EN.n197 EN.t33 132.282
R11113 EN.n186 EN.t60 132.282
R11114 EN.n175 EN.t3 132.282
R11115 EN.n164 EN.t67 132.282
R11116 EN.n153 EN.t57 132.282
R11117 EN.n103 EN.t68 132.282
R11118 EN.n146 EN.t77 132.282
R11119 EN.n137 EN.t13 132.282
R11120 EN.n128 EN.t71 132.282
R11121 EN.n119 EN.t42 132.282
R11122 EN.n111 EN.t37 132.282
R11123 EN.n89 EN.t8 132.282
R11124 EN.n79 EN.t80 132.282
R11125 EN.n48 EN.t21 132.282
R11126 EN.n57 EN.t19 132.282
R11127 EN.n67 EN.t66 132.282
R11128 EN.n38 EN.t41 132.282
R11129 EN.n29 EN.t45 132.282
R11130 EN.n19 EN.t53 132.282
R11131 EN.n9 EN.t25 132.282
R11132 EN.n0 EN.t34 132.282
R11133 EN EN.n222 42.8643
R11134 EN.n219 EN.n218 40.5582
R11135 EN EN.n221 36.3403
R11136 EN.n222 EN 35.9948
R11137 EN EN.n207 14.0185
R11138 EN EN.n196 14.0185
R11139 EN EN.n185 14.0185
R11140 EN EN.n174 14.0185
R11141 EN EN.n163 14.0185
R11142 EN EN.n152 14.0185
R11143 EN EN.n99 14.0185
R11144 EN EN.n142 14.0185
R11145 EN EN.n133 14.0185
R11146 EN EN.n124 14.0185
R11147 EN EN.n115 14.0185
R11148 EN EN.n107 14.0185
R11149 EN.n97 EN 13.8362
R11150 EN.n87 EN 13.8362
R11151 EN.n27 EN 13.8362
R11152 EN.n17 EN 13.8362
R11153 EN.n8 EN 13.8362
R11154 EN.n52 EN.n50 12.0681
R11155 EN.n61 EN.n59 12.0681
R11156 EN.n71 EN.n69 12.0681
R11157 EN.n42 EN.n40 12.0681
R11158 EN.n33 EN.n31 12.0681
R11159 EN.n54 EN.n53 9.86717
R11160 EN.n63 EN.n62 9.86717
R11161 EN.n73 EN.n72 9.86717
R11162 EN.n44 EN.n43 9.86717
R11163 EN.n35 EN.n34 9.86717
R11164 EN EN.n102 9.38671
R11165 EN EN.n145 9.38671
R11166 EN EN.n136 9.38671
R11167 EN EN.n127 9.38671
R11168 EN EN.n118 9.38671
R11169 EN EN.n110 9.38671
R11170 EN.n214 EN.n213 9.3005
R11171 EN.n216 EN.n207 9.3005
R11172 EN.n203 EN.n202 9.3005
R11173 EN.n205 EN.n196 9.3005
R11174 EN.n192 EN.n191 9.3005
R11175 EN.n194 EN.n185 9.3005
R11176 EN.n181 EN.n180 9.3005
R11177 EN.n183 EN.n174 9.3005
R11178 EN.n170 EN.n169 9.3005
R11179 EN.n172 EN.n163 9.3005
R11180 EN.n159 EN.n158 9.3005
R11181 EN.n161 EN.n152 9.3005
R11182 EN.n106 EN.n99 9.3005
R11183 EN.n149 EN.n142 9.3005
R11184 EN.n140 EN.n133 9.3005
R11185 EN.n131 EN.n124 9.3005
R11186 EN.n122 EN.n115 9.3005
R11187 EN.n114 EN.n107 9.3005
R11188 EN.n95 EN.n94 9.3005
R11189 EN.n85 EN.n84 9.3005
R11190 EN.n55 EN.n54 9.3005
R11191 EN.n64 EN.n63 9.3005
R11192 EN.n74 EN.n73 9.3005
R11193 EN.n45 EN.n44 9.3005
R11194 EN.n36 EN.n35 9.3005
R11195 EN.n25 EN.n24 9.3005
R11196 EN.n15 EN.n14 9.3005
R11197 EN.n6 EN.n5 9.3005
R11198 EN.n66 EN.n56 9.14473
R11199 EN.n47 EN.n37 9.14473
R11200 EN.n18 EN.n8 9.14473
R11201 EN.n123 EN.n114 9.106
R11202 EN.n53 EN.n52 8.82212
R11203 EN.n62 EN.n61 8.82212
R11204 EN.n72 EN.n71 8.82212
R11205 EN.n43 EN.n42 8.82212
R11206 EN.n34 EN.n33 8.82212
R11207 EN.n78 EN.n77 7.40722
R11208 EN.n162 EN.n151 7.28699
R11209 EN.n212 EN 4.67077
R11210 EN.n201 EN 4.67077
R11211 EN.n190 EN 4.67077
R11212 EN.n179 EN 4.67077
R11213 EN.n168 EN 4.67077
R11214 EN.n157 EN 4.67077
R11215 EN.n101 EN 4.67077
R11216 EN.n144 EN 4.67077
R11217 EN.n135 EN 4.67077
R11218 EN.n126 EN 4.67077
R11219 EN.n117 EN 4.67077
R11220 EN.n109 EN 4.67077
R11221 EN.n93 EN 4.67077
R11222 EN.n83 EN 4.67077
R11223 EN.n23 EN 4.67077
R11224 EN.n13 EN 4.67077
R11225 EN.n4 EN 4.67077
R11226 EN.n218 EN.n217 4.647
R11227 EN.n76 EN.n66 4.64473
R11228 EN.n28 EN.n18 4.64473
R11229 EN.n98 EN.n88 4.64473
R11230 EN.n132 EN.n123 4.606
R11231 EN.n141 EN.n132 4.606
R11232 EN.n150 EN.n141 4.606
R11233 EN.n184 EN.n173 4.606
R11234 EN.n195 EN.n184 4.606
R11235 EN.n206 EN.n195 4.606
R11236 EN.n217 EN.n206 4.606
R11237 EN.n151 EN.n150 4.58461
R11238 EN.n173 EN.n162 4.58461
R11239 EN.n207 EN 4.53383
R11240 EN.n196 EN 4.53383
R11241 EN.n185 EN 4.53383
R11242 EN.n174 EN 4.53383
R11243 EN.n163 EN 4.53383
R11244 EN.n152 EN 4.53383
R11245 EN.n99 EN 4.53383
R11246 EN.n142 EN 4.53383
R11247 EN.n133 EN 4.53383
R11248 EN.n124 EN 4.53383
R11249 EN.n115 EN 4.53383
R11250 EN.n107 EN 4.53383
R11251 EN.n54 EN 4.53383
R11252 EN.n63 EN 4.53383
R11253 EN.n73 EN 4.53383
R11254 EN.n44 EN 4.53383
R11255 EN.n35 EN 4.53383
R11256 EN.n123 EN.n122 4.5005
R11257 EN.n132 EN.n131 4.5005
R11258 EN.n141 EN.n140 4.5005
R11259 EN.n150 EN.n149 4.5005
R11260 EN.n151 EN.n106 4.5005
R11261 EN.n162 EN.n161 4.5005
R11262 EN.n173 EN.n172 4.5005
R11263 EN.n184 EN.n183 4.5005
R11264 EN.n195 EN.n194 4.5005
R11265 EN.n206 EN.n205 4.5005
R11266 EN.n217 EN.n216 4.5005
R11267 EN.n76 EN.n75 4.5005
R11268 EN.n66 EN.n65 4.5005
R11269 EN.n47 EN.n46 4.5005
R11270 EN.n18 EN.n17 4.5005
R11271 EN.n28 EN.n27 4.5005
R11272 EN.n88 EN.n87 4.5005
R11273 EN.n98 EN.n97 4.5005
R11274 EN EN.n98 4.39593
R11275 EN.n222 EN.n219 4.33925
R11276 EN.n88 EN.n78 4.15135
R11277 EN.n213 EN 2.94104
R11278 EN.n202 EN 2.94104
R11279 EN.n191 EN 2.94104
R11280 EN.n180 EN 2.94104
R11281 EN.n169 EN 2.94104
R11282 EN.n158 EN 2.94104
R11283 EN.n102 EN 2.94104
R11284 EN.n145 EN 2.94104
R11285 EN.n136 EN 2.94104
R11286 EN.n127 EN 2.94104
R11287 EN.n118 EN 2.94104
R11288 EN.n110 EN 2.94104
R11289 EN.n94 EN 2.94104
R11290 EN.n84 EN 2.94104
R11291 EN.n24 EN 2.94104
R11292 EN.n14 EN 2.94104
R11293 EN.n5 EN 2.94104
R11294 EN.n213 EN.n212 2.76807
R11295 EN.n202 EN.n201 2.76807
R11296 EN.n191 EN.n190 2.76807
R11297 EN.n180 EN.n179 2.76807
R11298 EN.n169 EN.n168 2.76807
R11299 EN.n158 EN.n157 2.76807
R11300 EN.n102 EN.n101 2.76807
R11301 EN.n145 EN.n144 2.76807
R11302 EN.n136 EN.n135 2.76807
R11303 EN.n127 EN.n126 2.76807
R11304 EN.n118 EN.n117 2.76807
R11305 EN.n110 EN.n109 2.76807
R11306 EN.n94 EN.n93 2.76807
R11307 EN.n84 EN.n83 2.76807
R11308 EN.n24 EN.n23 2.76807
R11309 EN.n14 EN.n13 2.76807
R11310 EN.n5 EN.n4 2.76807
R11311 EN.n77 EN.n47 2.55338
R11312 EN EN.n210 2.36657
R11313 EN EN.n199 2.36657
R11314 EN EN.n188 2.36657
R11315 EN EN.n177 2.36657
R11316 EN EN.n166 2.36657
R11317 EN EN.n155 2.36657
R11318 EN EN.n105 2.36657
R11319 EN EN.n148 2.36657
R11320 EN EN.n139 2.36657
R11321 EN EN.n130 2.36657
R11322 EN EN.n121 2.36657
R11323 EN EN.n113 2.36657
R11324 EN EN.n91 2.36657
R11325 EN EN.n81 2.36657
R11326 EN.n49 EN 2.36657
R11327 EN.n58 EN 2.36657
R11328 EN.n68 EN 2.36657
R11329 EN.n39 EN 2.36657
R11330 EN.n30 EN 2.36657
R11331 EN EN.n21 2.36657
R11332 EN EN.n11 2.36657
R11333 EN EN.n2 2.36657
R11334 EN.n219 EN 2.12425
R11335 EN.n77 EN.n76 2.04377
R11336 EN.n53 EN 1.73023
R11337 EN.n62 EN 1.73023
R11338 EN.n72 EN 1.73023
R11339 EN.n43 EN 1.73023
R11340 EN.n34 EN 1.73023
R11341 EN.n210 EN 0.580857
R11342 EN.n199 EN 0.580857
R11343 EN.n188 EN 0.580857
R11344 EN.n177 EN 0.580857
R11345 EN.n166 EN 0.580857
R11346 EN.n155 EN 0.580857
R11347 EN.n105 EN 0.580857
R11348 EN.n148 EN 0.580857
R11349 EN.n139 EN 0.580857
R11350 EN.n130 EN 0.580857
R11351 EN.n121 EN 0.580857
R11352 EN.n113 EN 0.580857
R11353 EN.n91 EN 0.580857
R11354 EN.n81 EN 0.580857
R11355 EN.n21 EN 0.580857
R11356 EN.n11 EN 0.580857
R11357 EN.n2 EN 0.580857
R11358 EN.n49 EN 0.527286
R11359 EN.n58 EN 0.527286
R11360 EN.n68 EN 0.527286
R11361 EN.n39 EN 0.527286
R11362 EN.n30 EN 0.527286
R11363 EN.n78 EN.n28 0.478275
R11364 EN.n221 EN 0.24431
R11365 EN.n209 EN 0.225552
R11366 EN.n198 EN 0.225552
R11367 EN.n187 EN 0.225552
R11368 EN.n176 EN 0.225552
R11369 EN.n165 EN 0.225552
R11370 EN.n154 EN 0.225552
R11371 EN.n104 EN 0.225552
R11372 EN.n147 EN 0.225552
R11373 EN.n138 EN 0.225552
R11374 EN.n129 EN 0.225552
R11375 EN.n120 EN 0.225552
R11376 EN.n112 EN 0.225552
R11377 EN.n90 EN 0.225552
R11378 EN.n80 EN 0.225552
R11379 EN.n20 EN 0.225552
R11380 EN.n10 EN 0.225552
R11381 EN.n1 EN 0.225552
R11382 EN.n106 EN 0.203203
R11383 EN.n149 EN 0.203203
R11384 EN.n140 EN 0.203203
R11385 EN.n131 EN 0.203203
R11386 EN.n122 EN 0.203203
R11387 EN.n114 EN 0.203203
R11388 EN.n215 EN 0.139923
R11389 EN.n204 EN 0.139923
R11390 EN.n193 EN 0.139923
R11391 EN.n182 EN 0.139923
R11392 EN.n171 EN 0.139923
R11393 EN.n160 EN 0.139923
R11394 EN.n96 EN 0.139923
R11395 EN.n86 EN 0.139923
R11396 EN.n26 EN 0.139923
R11397 EN.n16 EN 0.139923
R11398 EN.n7 EN 0.139923
R11399 EN.n210 EN.n209 0.128681
R11400 EN.n199 EN.n198 0.128681
R11401 EN.n188 EN.n187 0.128681
R11402 EN.n177 EN.n176 0.128681
R11403 EN.n166 EN.n165 0.128681
R11404 EN.n155 EN.n154 0.128681
R11405 EN.n105 EN.n104 0.128681
R11406 EN.n148 EN.n147 0.128681
R11407 EN.n139 EN.n138 0.128681
R11408 EN.n130 EN.n129 0.128681
R11409 EN.n121 EN.n120 0.128681
R11410 EN.n113 EN.n112 0.128681
R11411 EN.n91 EN.n90 0.128681
R11412 EN.n81 EN.n80 0.128681
R11413 EN.n21 EN.n20 0.128681
R11414 EN.n11 EN.n10 0.128681
R11415 EN.n2 EN.n1 0.128681
R11416 EN.n56 EN 0.0726154
R11417 EN.n65 EN 0.0726154
R11418 EN.n75 EN 0.0726154
R11419 EN.n46 EN 0.0726154
R11420 EN.n37 EN 0.0726154
R11421 EN.n216 EN 0.0702115
R11422 EN.n205 EN 0.0702115
R11423 EN.n194 EN 0.0702115
R11424 EN.n183 EN 0.0702115
R11425 EN.n172 EN 0.0702115
R11426 EN.n161 EN 0.0702115
R11427 EN.n55 EN 0.0702115
R11428 EN.n64 EN 0.0702115
R11429 EN.n74 EN 0.0702115
R11430 EN.n45 EN 0.0702115
R11431 EN.n36 EN 0.0702115
R11432 EN.n97 EN 0.0678077
R11433 EN.n87 EN 0.0678077
R11434 EN.n27 EN 0.0678077
R11435 EN.n17 EN 0.0678077
R11436 EN.n8 EN 0.0678077
R11437 EN.n106 EN 0.0664091
R11438 EN.n149 EN 0.0664091
R11439 EN.n140 EN 0.0664091
R11440 EN.n131 EN 0.0664091
R11441 EN.n122 EN 0.0664091
R11442 EN.n114 EN 0.0664091
R11443 EN.n214 EN 0.03675
R11444 EN.n203 EN 0.03675
R11445 EN.n192 EN 0.03675
R11446 EN.n181 EN 0.03675
R11447 EN.n170 EN 0.03675
R11448 EN.n159 EN 0.03675
R11449 EN.n95 EN 0.03675
R11450 EN.n85 EN 0.03675
R11451 EN.n50 EN.n49 0.03675
R11452 EN.n59 EN.n58 0.03675
R11453 EN.n69 EN.n68 0.03675
R11454 EN.n40 EN.n39 0.03675
R11455 EN.n31 EN.n30 0.03675
R11456 EN.n25 EN 0.03675
R11457 EN.n15 EN 0.03675
R11458 EN.n6 EN 0.03675
R11459 EN.n50 EN 0.0366675
R11460 EN.n59 EN 0.0366675
R11461 EN.n69 EN 0.0366675
R11462 EN.n40 EN 0.0366675
R11463 EN.n31 EN 0.0366675
R11464 EN.n96 EN.n95 0.036656
R11465 EN.n86 EN.n85 0.036656
R11466 EN.n26 EN.n25 0.036656
R11467 EN.n16 EN.n15 0.036656
R11468 EN.n7 EN.n6 0.036656
R11469 EN.n215 EN.n214 0.0365577
R11470 EN.n204 EN.n203 0.0365577
R11471 EN.n193 EN.n192 0.0365577
R11472 EN.n182 EN.n181 0.0365577
R11473 EN.n171 EN.n170 0.0365577
R11474 EN.n160 EN.n159 0.0365577
R11475 EN.n218 EN 0.0293462
R11476 EN EN.n215 0.00530769
R11477 EN EN.n204 0.00530769
R11478 EN EN.n193 0.00530769
R11479 EN EN.n182 0.00530769
R11480 EN EN.n171 0.00530769
R11481 EN EN.n160 0.00530769
R11482 EN EN.n96 0.00530769
R11483 EN EN.n86 0.00530769
R11484 EN EN.n26 0.00530769
R11485 EN EN.n16 0.00530769
R11486 EN EN.n7 0.00530769
R11487 EN.n56 EN.n55 0.00290385
R11488 EN.n65 EN.n64 0.00290385
R11489 EN.n75 EN.n74 0.00290385
R11490 EN.n46 EN.n45 0.00290385
R11491 EN.n37 EN.n36 0.00290385
R11492 a_4597_n5258.t0 a_4597_n5258.n0 1327.82
R11493 a_4597_n5258.n0 a_4597_n5258.t2 194.655
R11494 a_4597_n5258.n0 a_4597_n5258.t1 63.3219
R11495 a_8583_n1331.n1 a_8583_n1331.t5 530.01
R11496 a_8583_n1331.t1 a_8583_n1331.n5 421.021
R11497 a_8583_n1331.n0 a_8583_n1331.t6 337.171
R11498 a_8583_n1331.n3 a_8583_n1331.t0 280.223
R11499 a_8583_n1331.n4 a_8583_n1331.t4 263.173
R11500 a_8583_n1331.n4 a_8583_n1331.t2 227.826
R11501 a_8583_n1331.n0 a_8583_n1331.t7 199.762
R11502 a_8583_n1331.n2 a_8583_n1331.n1 170.81
R11503 a_8583_n1331.n2 a_8583_n1331.n0 167.321
R11504 a_8583_n1331.n5 a_8583_n1331.n4 152
R11505 a_8583_n1331.n1 a_8583_n1331.t3 141.923
R11506 a_8583_n1331.n3 a_8583_n1331.n2 10.8376
R11507 a_8583_n1331.n5 a_8583_n1331.n3 2.50485
R11508 a_8544_n1457.t1 a_8544_n1457.n3 370.026
R11509 a_8544_n1457.n0 a_8544_n1457.t4 351.356
R11510 a_8544_n1457.n1 a_8544_n1457.t5 334.717
R11511 a_8544_n1457.n3 a_8544_n1457.t0 325.971
R11512 a_8544_n1457.n1 a_8544_n1457.t3 309.935
R11513 a_8544_n1457.n0 a_8544_n1457.t2 305.683
R11514 a_8544_n1457.n2 a_8544_n1457.n0 16.879
R11515 a_8544_n1457.n3 a_8544_n1457.n2 10.8867
R11516 a_8544_n1457.n2 a_8544_n1457.n1 9.3005
R11517 a_1479_3531.n5 a_1479_3531.n4 807.871
R11518 a_1479_3531.n2 a_1479_3531.t7 389.183
R11519 a_1479_3531.n3 a_1479_3531.n2 251.167
R11520 a_1479_3531.n3 a_1479_3531.t2 223.571
R11521 a_1479_3531.n0 a_1479_3531.t4 212.081
R11522 a_1479_3531.n1 a_1479_3531.t5 212.081
R11523 a_1479_3531.n4 a_1479_3531.n1 176.576
R11524 a_1479_3531.n2 a_1479_3531.t3 174.891
R11525 a_1479_3531.n0 a_1479_3531.t6 139.78
R11526 a_1479_3531.n1 a_1479_3531.t8 139.78
R11527 a_1479_3531.n5 a_1479_3531.t1 63.3219
R11528 a_1479_3531.t0 a_1479_3531.n5 63.3219
R11529 a_1479_3531.n1 a_1479_3531.n0 61.346
R11530 a_1479_3531.n4 a_1479_3531.n3 37.7195
R11531 a_1413_3557.t0 a_1413_3557.t1 94.7268
R11532 a_5311_n1055.n5 a_5311_n1055.n4 807.871
R11533 a_5311_n1055.n2 a_5311_n1055.t3 389.183
R11534 a_5311_n1055.n3 a_5311_n1055.n2 251.167
R11535 a_5311_n1055.n3 a_5311_n1055.t1 223.571
R11536 a_5311_n1055.n0 a_5311_n1055.t4 212.081
R11537 a_5311_n1055.n1 a_5311_n1055.t6 212.081
R11538 a_5311_n1055.n4 a_5311_n1055.n1 176.576
R11539 a_5311_n1055.n2 a_5311_n1055.t5 174.891
R11540 a_5311_n1055.n0 a_5311_n1055.t7 139.78
R11541 a_5311_n1055.n1 a_5311_n1055.t8 139.78
R11542 a_5311_n1055.t0 a_5311_n1055.n5 63.3219
R11543 a_5311_n1055.n5 a_5311_n1055.t2 63.3219
R11544 a_5311_n1055.n1 a_5311_n1055.n0 61.346
R11545 a_5311_n1055.n4 a_5311_n1055.n3 37.7195
R11546 a_8099_n10022.n1 a_8099_n10022.t3 530.01
R11547 a_8099_n10022.t0 a_8099_n10022.n5 421.021
R11548 a_8099_n10022.n0 a_8099_n10022.t6 337.142
R11549 a_8099_n10022.n3 a_8099_n10022.t1 280.223
R11550 a_8099_n10022.n4 a_8099_n10022.t5 263.173
R11551 a_8099_n10022.n4 a_8099_n10022.t4 227.826
R11552 a_8099_n10022.n0 a_8099_n10022.t7 199.762
R11553 a_8099_n10022.n2 a_8099_n10022.n1 170.81
R11554 a_8099_n10022.n2 a_8099_n10022.n0 167.321
R11555 a_8099_n10022.n5 a_8099_n10022.n4 152
R11556 a_8099_n10022.n1 a_8099_n10022.t2 141.923
R11557 a_8099_n10022.n3 a_8099_n10022.n2 10.8376
R11558 a_8099_n10022.n5 a_8099_n10022.n3 2.50485
R11559 a_8615_n9650.n3 a_8615_n9650.n2 674.338
R11560 a_8615_n9650.n1 a_8615_n9650.t4 332.58
R11561 a_8615_n9650.n2 a_8615_n9650.n0 284.012
R11562 a_8615_n9650.n2 a_8615_n9650.n1 253.648
R11563 a_8615_n9650.n1 a_8615_n9650.t5 168.701
R11564 a_8615_n9650.t0 a_8615_n9650.n3 96.1553
R11565 a_8615_n9650.n3 a_8615_n9650.t3 65.6672
R11566 a_8615_n9650.n0 a_8615_n9650.t1 65.0005
R11567 a_8615_n9650.n0 a_8615_n9650.t2 45.0005
R11568 a_8077_n5258.t0 a_8077_n5258.t1 126.644
R11569 a_7843_n5372.n3 a_7843_n5372.n2 636.953
R11570 a_7843_n5372.n1 a_7843_n5372.t4 366.856
R11571 a_7843_n5372.n2 a_7843_n5372.n0 300.2
R11572 a_7843_n5372.n2 a_7843_n5372.n1 225.036
R11573 a_7843_n5372.n1 a_7843_n5372.t5 174.056
R11574 a_7843_n5372.n0 a_7843_n5372.t1 70.0005
R11575 a_7843_n5372.n3 a_7843_n5372.t2 68.0124
R11576 a_7843_n5372.t0 a_7843_n5372.n3 63.3219
R11577 a_7843_n5372.n0 a_7843_n5372.t3 61.6672
R11578 a_n975_3799.n3 a_n975_3799.n2 647.119
R11579 a_n975_3799.n1 a_n975_3799.t5 350.253
R11580 a_n975_3799.n2 a_n975_3799.n0 260.339
R11581 a_n975_3799.n2 a_n975_3799.n1 246.119
R11582 a_n975_3799.n1 a_n975_3799.t4 189.588
R11583 a_n975_3799.n3 a_n975_3799.t1 89.1195
R11584 a_n975_3799.n0 a_n975_3799.t0 63.3338
R11585 a_n975_3799.t3 a_n975_3799.n3 41.0422
R11586 a_n975_3799.n0 a_n975_3799.t2 31.9797
R11587 a_5564_n5074.n1 a_5564_n5074.t5 530.01
R11588 a_5564_n5074.t1 a_5564_n5074.n5 421.021
R11589 a_5564_n5074.n0 a_5564_n5074.t7 337.142
R11590 a_5564_n5074.n3 a_5564_n5074.t0 280.223
R11591 a_5564_n5074.n4 a_5564_n5074.t6 263.173
R11592 a_5564_n5074.n4 a_5564_n5074.t3 227.826
R11593 a_5564_n5074.n0 a_5564_n5074.t2 199.762
R11594 a_5564_n5074.n2 a_5564_n5074.n1 170.81
R11595 a_5564_n5074.n2 a_5564_n5074.n0 167.321
R11596 a_5564_n5074.n5 a_5564_n5074.n4 152
R11597 a_5564_n5074.n1 a_5564_n5074.t4 141.923
R11598 a_5564_n5074.n3 a_5564_n5074.n2 10.8376
R11599 a_5564_n5074.n5 a_5564_n5074.n3 2.50485
R11600 a_6645_n4702.n3 a_6645_n4702.n2 636.953
R11601 a_6645_n4702.n1 a_6645_n4702.t4 366.856
R11602 a_6645_n4702.n2 a_6645_n4702.n0 300.2
R11603 a_6645_n4702.n2 a_6645_n4702.n1 225.036
R11604 a_6645_n4702.n1 a_6645_n4702.t5 174.056
R11605 a_6645_n4702.n0 a_6645_n4702.t2 70.0005
R11606 a_6645_n4702.t0 a_6645_n4702.n3 68.0124
R11607 a_6645_n4702.n3 a_6645_n4702.t3 63.3219
R11608 a_6645_n4702.n0 a_6645_n4702.t1 61.6672
R11609 a_6754_n4702.n0 a_6754_n4702.t0 68.3338
R11610 a_6754_n4702.n0 a_6754_n4702.t1 26.3935
R11611 a_6754_n4702.n1 a_6754_n4702.n0 14.4005
R11612 a_9175_n1055.n5 a_9175_n1055.n4 807.871
R11613 a_9175_n1055.n2 a_9175_n1055.t4 389.183
R11614 a_9175_n1055.n3 a_9175_n1055.n2 251.167
R11615 a_9175_n1055.n3 a_9175_n1055.t2 223.571
R11616 a_9175_n1055.n0 a_9175_n1055.t6 212.081
R11617 a_9175_n1055.n1 a_9175_n1055.t3 212.081
R11618 a_9175_n1055.n4 a_9175_n1055.n1 176.576
R11619 a_9175_n1055.n2 a_9175_n1055.t8 174.891
R11620 a_9175_n1055.n0 a_9175_n1055.t7 139.78
R11621 a_9175_n1055.n1 a_9175_n1055.t5 139.78
R11622 a_9175_n1055.t0 a_9175_n1055.n5 63.3219
R11623 a_9175_n1055.n5 a_9175_n1055.t1 63.3219
R11624 a_9175_n1055.n1 a_9175_n1055.n0 61.346
R11625 a_9175_n1055.n4 a_9175_n1055.n3 37.7195
R11626 CF[5].n10 CF[5].n9 585
R11627 CF[5].n11 CF[5].n10 585
R11628 CF[5].n6 CF[5].t9 332.312
R11629 CF[5].n6 CF[5].t5 295.627
R11630 CF[5].n3 CF[5].t6 294.557
R11631 CF[5].n0 CF[5].t7 294.557
R11632 CF[5].n3 CF[5].t4 211.01
R11633 CF[5].n0 CF[5].t8 211.01
R11634 CF[5] CF[5].n6 196.004
R11635 CF[5].n8 CF[5].n7 185
R11636 CF[5].n4 CF[5].n3 153.097
R11637 CF[5].n1 CF[5].n0 152
R11638 CF[5] CF[5].n13 53.5834
R11639 CF[5] CF[5].n8 49.0339
R11640 CF[5].n10 CF[5].t2 26.5955
R11641 CF[5].n10 CF[5].t3 26.5955
R11642 CF[5].n7 CF[5].t0 24.9236
R11643 CF[5].n7 CF[5].t1 24.9236
R11644 CF[5].n12 CF[5].n11 16.4548
R11645 CF[5].n9 CF[5] 15.6165
R11646 CF[5].n13 CF[5] 15.2722
R11647 CF[5].n5 CF[5].n2 14.9321
R11648 CF[5].n5 CF[5].n4 13.9063
R11649 CF[5].n8 CF[5] 10.4965
R11650 CF[5].n2 CF[5] 9.32621
R11651 CF[5].n13 CF[5] 6.05175
R11652 CF[5].n12 CF[5] 3.11923
R11653 CF[5].n4 CF[5] 3.10907
R11654 CF[5].n1 CF[5] 2.01193
R11655 CF[5].n11 CF[5] 1.7925
R11656 CF[5].n9 CF[5] 1.7925
R11657 CF[5].n2 CF[5].n1 1.09764
R11658 CF[5] CF[5].n5 0.843172
R11659 CF[5] CF[5].n12 0.778096
R11660 a_7950_2717.n1 a_7950_2717.t3 530.01
R11661 a_7950_2717.t1 a_7950_2717.n5 421.021
R11662 a_7950_2717.n0 a_7950_2717.t7 337.142
R11663 a_7950_2717.n3 a_7950_2717.t0 280.223
R11664 a_7950_2717.n4 a_7950_2717.t5 263.173
R11665 a_7950_2717.n4 a_7950_2717.t4 227.826
R11666 a_7950_2717.n0 a_7950_2717.t6 199.762
R11667 a_7950_2717.n2 a_7950_2717.n1 170.81
R11668 a_7950_2717.n2 a_7950_2717.n0 167.321
R11669 a_7950_2717.n5 a_7950_2717.n4 152
R11670 a_7950_2717.n1 a_7950_2717.t2 141.923
R11671 a_7950_2717.n3 a_7950_2717.n2 10.8376
R11672 a_7950_2717.n5 a_7950_2717.n3 2.50485
R11673 a_8371_2717.n1 a_8371_2717.n0 926.024
R11674 a_8371_2717.t1 a_8371_2717.n1 82.0838
R11675 a_8371_2717.n0 a_8371_2717.t0 63.3338
R11676 a_8371_2717.n1 a_8371_2717.t3 63.3219
R11677 a_8371_2717.n0 a_8371_2717.t2 29.7268
R11678 a_8466_2717.n3 a_8466_2717.n2 674.338
R11679 a_8466_2717.n1 a_8466_2717.t4 332.58
R11680 a_8466_2717.n2 a_8466_2717.n0 284.012
R11681 a_8466_2717.n2 a_8466_2717.n1 253.648
R11682 a_8466_2717.n1 a_8466_2717.t5 168.701
R11683 a_8466_2717.t0 a_8466_2717.n3 96.1553
R11684 a_8466_2717.n3 a_8466_2717.t2 65.6672
R11685 a_8466_2717.n0 a_8466_2717.t1 65.0005
R11686 a_8466_2717.n0 a_8466_2717.t3 45.0005
R11687 CF[4].n9 CF[4].n8 585
R11688 CF[4].n10 CF[4].n9 585
R11689 CF[4].n12 CF[4].t5 332.312
R11690 CF[4].n12 CF[4].t6 295.627
R11691 CF[4].n3 CF[4].t8 294.557
R11692 CF[4].n0 CF[4].t7 294.557
R11693 CF[4].n3 CF[4].t4 211.01
R11694 CF[4].n0 CF[4].t9 211.01
R11695 CF[4] CF[4].n12 196.004
R11696 CF[4].n7 CF[4].n6 185
R11697 CF[4].n4 CF[4].n3 153.097
R11698 CF[4].n1 CF[4].n0 152
R11699 CF[4] CF[4].n7 57.7379
R11700 CF[4] CF[4].n15 55.7291
R11701 CF[4].n13 CF[4] 37.1376
R11702 CF[4].n9 CF[4].t2 26.5955
R11703 CF[4].n9 CF[4].t3 26.5955
R11704 CF[4].n6 CF[4].t0 24.9236
R11705 CF[4].n6 CF[4].t1 24.9236
R11706 CF[4].n15 CF[4].n14 19.926
R11707 CF[4].n5 CF[4].n2 14.9321
R11708 CF[4].n13 CF[4].n11 14.7472
R11709 CF[4].n5 CF[4].n4 13.9063
R11710 CF[4].n8 CF[4] 10.4965
R11711 CF[4].n10 CF[4] 10.4965
R11712 CF[4].n2 CF[4] 9.32621
R11713 CF[4].n15 CF[4] 8.1005
R11714 CF[4].n8 CF[4] 6.9125
R11715 CF[4].n11 CF[4] 4.3525
R11716 CF[4].n4 CF[4] 3.10907
R11717 CF[4].n11 CF[4].n10 2.5605
R11718 CF[4].n1 CF[4] 2.01193
R11719 CF[4].n7 CF[4] 1.7925
R11720 CF[4].n2 CF[4].n1 1.09764
R11721 CF[4].n14 CF[4].n13 0.865885
R11722 CF[4] CF[4].n5 0.856103
R11723 CF[4].n14 CF[4] 0.0341538
R11724 a_n1561_n10022.n1 a_n1561_n10022.t3 530.01
R11725 a_n1561_n10022.t1 a_n1561_n10022.n5 421.021
R11726 a_n1561_n10022.n0 a_n1561_n10022.t5 337.142
R11727 a_n1561_n10022.n3 a_n1561_n10022.t0 280.223
R11728 a_n1561_n10022.n4 a_n1561_n10022.t4 263.173
R11729 a_n1561_n10022.n4 a_n1561_n10022.t7 227.826
R11730 a_n1561_n10022.n0 a_n1561_n10022.t6 199.762
R11731 a_n1561_n10022.n2 a_n1561_n10022.n1 170.81
R11732 a_n1561_n10022.n2 a_n1561_n10022.n0 167.321
R11733 a_n1561_n10022.n5 a_n1561_n10022.n4 152
R11734 a_n1561_n10022.n1 a_n1561_n10022.t2 141.923
R11735 a_n1561_n10022.n3 a_n1561_n10022.n2 10.8376
R11736 a_n1561_n10022.n5 a_n1561_n10022.n3 2.50485
R11737 CF[8].n11 CF[8].n10 585
R11738 CF[8].n12 CF[8].n11 585
R11739 CF[8].n6 CF[8].t6 333.651
R11740 CF[8].n6 CF[8].t7 297.233
R11741 CF[8].n3 CF[8].t4 294.557
R11742 CF[8].n0 CF[8].t9 294.557
R11743 CF[8].n3 CF[8].t8 211.01
R11744 CF[8].n0 CF[8].t5 211.01
R11745 CF[8].n7 CF[8].n6 196.493
R11746 CF[8].n9 CF[8].n8 185
R11747 CF[8].n4 CF[8].n3 153.097
R11748 CF[8].n1 CF[8].n0 152
R11749 CF[8] CF[8].n9 49.0339
R11750 CF[8] CF[8].n14 41.5204
R11751 CF[8].n13 CF[8].n7 35.37
R11752 CF[8].n14 CF[8] 30.8106
R11753 CF[8].n11 CF[8].t0 26.5955
R11754 CF[8].n11 CF[8].t2 26.5955
R11755 CF[8].n8 CF[8].t1 24.9236
R11756 CF[8].n8 CF[8].t3 24.9236
R11757 CF[8].n13 CF[8].n12 17.2879
R11758 CF[8].n10 CF[8] 15.6165
R11759 CF[8].n5 CF[8].n2 14.9321
R11760 CF[8].n5 CF[8].n4 13.9063
R11761 CF[8].n9 CF[8] 10.4965
R11762 CF[8].n2 CF[8] 9.32621
R11763 CF[8].n14 CF[8] 5.613
R11764 CF[8].n4 CF[8] 3.10907
R11765 CF[8].n1 CF[8] 2.01193
R11766 CF[8].n12 CF[8] 1.7925
R11767 CF[8].n10 CF[8] 1.7925
R11768 CF[8].n2 CF[8].n1 1.09764
R11769 CF[8] CF[8].n5 0.843172
R11770 CF[8] CF[8].n13 0.740885
R11771 CF[8].n7 CF[8] 0.24431
R11772 a_6167_n10022.n1 a_6167_n10022.t5 530.01
R11773 a_6167_n10022.t1 a_6167_n10022.n5 421.021
R11774 a_6167_n10022.n0 a_6167_n10022.t7 337.142
R11775 a_6167_n10022.n3 a_6167_n10022.t0 280.223
R11776 a_6167_n10022.n4 a_6167_n10022.t6 263.173
R11777 a_6167_n10022.n4 a_6167_n10022.t4 227.826
R11778 a_6167_n10022.n0 a_6167_n10022.t2 199.762
R11779 a_6167_n10022.n2 a_6167_n10022.n1 170.81
R11780 a_6167_n10022.n2 a_6167_n10022.n0 167.321
R11781 a_6167_n10022.n5 a_6167_n10022.n4 152
R11782 a_6167_n10022.n1 a_6167_n10022.t3 141.923
R11783 a_6167_n10022.n3 a_6167_n10022.n2 10.8376
R11784 a_6167_n10022.n5 a_6167_n10022.n3 2.50485
R11785 a_6047_n1599.n4 a_6047_n1599.n1 807.871
R11786 a_6047_n1599.n0 a_6047_n1599.t4 389.183
R11787 a_6047_n1599.n5 a_6047_n1599.n0 251.167
R11788 a_6047_n1599.t0 a_6047_n1599.n5 223.571
R11789 a_6047_n1599.n3 a_6047_n1599.t8 212.081
R11790 a_6047_n1599.n2 a_6047_n1599.t3 212.081
R11791 a_6047_n1599.n4 a_6047_n1599.n3 176.576
R11792 a_6047_n1599.n0 a_6047_n1599.t7 174.891
R11793 a_6047_n1599.n3 a_6047_n1599.t5 139.78
R11794 a_6047_n1599.n2 a_6047_n1599.t6 139.78
R11795 a_6047_n1599.n1 a_6047_n1599.t2 63.3219
R11796 a_6047_n1599.n1 a_6047_n1599.t1 63.3219
R11797 a_6047_n1599.n3 a_6047_n1599.n2 61.346
R11798 a_6047_n1599.n5 a_6047_n1599.n4 37.5061
R11799 CF[3].n9 CF[3].n8 585
R11800 CF[3].n10 CF[3].n9 585
R11801 CF[3].n12 CF[3].t5 332.312
R11802 CF[3].n12 CF[3].t8 295.627
R11803 CF[3].n3 CF[3].t7 294.557
R11804 CF[3].n0 CF[3].t9 294.557
R11805 CF[3].n3 CF[3].t6 211.01
R11806 CF[3].n0 CF[3].t4 211.01
R11807 CF[3] CF[3].n12 196.004
R11808 CF[3].n7 CF[3].n6 185
R11809 CF[3].n4 CF[3].n3 153.097
R11810 CF[3].n1 CF[3].n0 152
R11811 CF[3] CF[3].n14 59.706
R11812 CF[3] CF[3].n7 57.7379
R11813 CF[3].n13 CF[3] 37.1376
R11814 CF[3].n9 CF[3].t2 26.5955
R11815 CF[3].n9 CF[3].t3 26.5955
R11816 CF[3].n6 CF[3].t1 24.9236
R11817 CF[3].n6 CF[3].t0 24.9236
R11818 CF[3].n14 CF[3] 24.3539
R11819 CF[3].n5 CF[3].n2 14.9321
R11820 CF[3].n13 CF[3].n11 14.7279
R11821 CF[3].n5 CF[3].n4 13.9063
R11822 CF[3].n8 CF[3] 10.4965
R11823 CF[3].n10 CF[3] 10.4965
R11824 CF[3].n2 CF[3] 9.32621
R11825 CF[3].n14 CF[3] 8.258
R11826 CF[3].n8 CF[3] 6.9125
R11827 CF[3].n11 CF[3] 4.3525
R11828 CF[3].n4 CF[3] 3.10907
R11829 CF[3].n11 CF[3].n10 2.5605
R11830 CF[3].n1 CF[3] 2.01193
R11831 CF[3].n7 CF[3] 1.7925
R11832 CF[3].n2 CF[3].n1 1.09764
R11833 CF[3] CF[3].n13 0.904346
R11834 CF[3] CF[3].n5 0.847483
R11835 a_4751_n9484.n3 a_4751_n9484.n2 674.338
R11836 a_4751_n9484.n1 a_4751_n9484.t4 332.58
R11837 a_4751_n9484.n2 a_4751_n9484.n0 284.012
R11838 a_4751_n9484.n2 a_4751_n9484.n1 253.648
R11839 a_4751_n9484.n1 a_4751_n9484.t5 168.701
R11840 a_4751_n9484.t0 a_4751_n9484.n3 96.1553
R11841 a_4751_n9484.n3 a_4751_n9484.t2 65.6672
R11842 a_4751_n9484.n0 a_4751_n9484.t1 65.0005
R11843 a_4751_n9484.n0 a_4751_n9484.t3 45.0005
R11844 a_4969_n9242.n3 a_4969_n9242.n2 647.119
R11845 a_4969_n9242.n1 a_4969_n9242.t5 350.253
R11846 a_4969_n9242.n2 a_4969_n9242.n0 260.339
R11847 a_4969_n9242.n2 a_4969_n9242.n1 246.119
R11848 a_4969_n9242.n1 a_4969_n9242.t4 189.588
R11849 a_4969_n9242.n3 a_4969_n9242.t2 89.1195
R11850 a_4969_n9242.n0 a_4969_n9242.t3 63.3338
R11851 a_4969_n9242.t1 a_4969_n9242.n3 41.0422
R11852 a_4969_n9242.n0 a_4969_n9242.t0 31.9797
R11853 a_502_n5106.n3 a_502_n5106.n2 647.119
R11854 a_502_n5106.n1 a_502_n5106.t5 350.253
R11855 a_502_n5106.n2 a_502_n5106.n0 260.339
R11856 a_502_n5106.n2 a_502_n5106.n1 246.119
R11857 a_502_n5106.n1 a_502_n5106.t4 189.588
R11858 a_502_n5106.n3 a_502_n5106.t1 89.1195
R11859 a_502_n5106.n0 a_502_n5106.t0 63.3338
R11860 a_502_n5106.t2 a_502_n5106.n3 41.0422
R11861 a_502_n5106.n0 a_502_n5106.t3 31.9797
R11862 a_392_n5080.t0 a_392_n5080.n0 1327.82
R11863 a_392_n5080.n0 a_392_n5080.t1 194.655
R11864 a_392_n5080.n0 a_392_n5080.t2 63.3219
R11865 a_1447_n1055.n5 a_1447_n1055.n4 807.871
R11866 a_1447_n1055.n2 a_1447_n1055.t7 389.183
R11867 a_1447_n1055.n3 a_1447_n1055.n2 251.167
R11868 a_1447_n1055.n3 a_1447_n1055.t1 223.571
R11869 a_1447_n1055.n0 a_1447_n1055.t8 212.081
R11870 a_1447_n1055.n1 a_1447_n1055.t6 212.081
R11871 a_1447_n1055.n4 a_1447_n1055.n1 176.576
R11872 a_1447_n1055.n2 a_1447_n1055.t3 174.891
R11873 a_1447_n1055.n0 a_1447_n1055.t5 139.78
R11874 a_1447_n1055.n1 a_1447_n1055.t4 139.78
R11875 a_1447_n1055.t0 a_1447_n1055.n5 63.3219
R11876 a_1447_n1055.n5 a_1447_n1055.t2 63.3219
R11877 a_1447_n1055.n1 a_1447_n1055.n0 61.346
R11878 a_1447_n1055.n4 a_1447_n1055.n3 37.7195
R11879 a_1381_n1029.t0 a_1381_n1029.t1 94.7268
R11880 a_1024_n4776.n4 a_1024_n4776.n1 807.871
R11881 a_1024_n4776.n0 a_1024_n4776.t3 389.183
R11882 a_1024_n4776.n5 a_1024_n4776.n0 251.167
R11883 a_1024_n4776.t0 a_1024_n4776.n5 223.571
R11884 a_1024_n4776.n2 a_1024_n4776.t7 212.081
R11885 a_1024_n4776.n3 a_1024_n4776.t6 212.081
R11886 a_1024_n4776.n4 a_1024_n4776.n3 176.576
R11887 a_1024_n4776.n0 a_1024_n4776.t4 174.891
R11888 a_1024_n4776.n2 a_1024_n4776.t5 139.78
R11889 a_1024_n4776.n3 a_1024_n4776.t8 139.78
R11890 a_1024_n4776.n1 a_1024_n4776.t1 63.3219
R11891 a_1024_n4776.n1 a_1024_n4776.t2 63.3219
R11892 a_1024_n4776.n3 a_1024_n4776.n2 61.346
R11893 a_1024_n4776.n5 a_1024_n4776.n4 37.7195
R11894 a_n937_n10028.n0 a_n937_n10028.t2 1327.82
R11895 a_n937_n10028.t0 a_n937_n10028.n0 194.655
R11896 a_n937_n10028.n0 a_n937_n10028.t1 63.3219
R11897 a_4235_n10022.n1 a_4235_n10022.t5 530.01
R11898 a_4235_n10022.t1 a_4235_n10022.n5 421.021
R11899 a_4235_n10022.n0 a_4235_n10022.t3 337.142
R11900 a_4235_n10022.n3 a_4235_n10022.t0 280.223
R11901 a_4235_n10022.n4 a_4235_n10022.t7 263.173
R11902 a_4235_n10022.n4 a_4235_n10022.t4 227.826
R11903 a_4235_n10022.n0 a_4235_n10022.t2 199.762
R11904 a_4235_n10022.n2 a_4235_n10022.n1 170.81
R11905 a_4235_n10022.n2 a_4235_n10022.n0 167.321
R11906 a_4235_n10022.n5 a_4235_n10022.n4 152
R11907 a_4235_n10022.n1 a_4235_n10022.t6 141.923
R11908 a_4235_n10022.n3 a_4235_n10022.n2 10.8376
R11909 a_4235_n10022.n5 a_4235_n10022.n3 2.50485
R11910 a_5316_n9650.n3 a_5316_n9650.n2 636.953
R11911 a_5316_n9650.n1 a_5316_n9650.t5 366.856
R11912 a_5316_n9650.n2 a_5316_n9650.n0 300.2
R11913 a_5316_n9650.n2 a_5316_n9650.n1 225.036
R11914 a_5316_n9650.n1 a_5316_n9650.t4 174.056
R11915 a_5316_n9650.n0 a_5316_n9650.t2 70.0005
R11916 a_5316_n9650.t1 a_5316_n9650.n3 68.0124
R11917 a_5316_n9650.n3 a_5316_n9650.t3 63.3219
R11918 a_5316_n9650.n0 a_5316_n9650.t0 61.6672
R11919 a_5425_n9650.n0 a_5425_n9650.t0 68.3338
R11920 a_5425_n9650.n0 a_5425_n9650.t1 26.3935
R11921 a_5425_n9650.n1 a_5425_n9650.n0 14.4005
R11922 a_6189_n5356.t0 a_6189_n5356.n3 370.026
R11923 a_6189_n5356.n0 a_6189_n5356.t5 351.356
R11924 a_6189_n5356.n1 a_6189_n5356.t4 334.717
R11925 a_6189_n5356.n3 a_6189_n5356.t1 325.971
R11926 a_6189_n5356.n1 a_6189_n5356.t2 309.935
R11927 a_6189_n5356.n0 a_6189_n5356.t3 305.683
R11928 a_6189_n5356.n2 a_6189_n5356.n0 16.879
R11929 a_6189_n5356.n3 a_6189_n5356.n2 10.8867
R11930 a_6189_n5356.n2 a_6189_n5356.n1 9.3005
R11931 a_6384_n5387.n3 a_6384_n5387.n2 674.338
R11932 a_6384_n5387.n1 a_6384_n5387.t4 332.58
R11933 a_6384_n5387.n2 a_6384_n5387.n0 284.012
R11934 a_6384_n5387.n2 a_6384_n5387.n1 253.648
R11935 a_6384_n5387.n1 a_6384_n5387.t5 168.701
R11936 a_6384_n5387.n3 a_6384_n5387.t3 96.1553
R11937 a_6384_n5387.t1 a_6384_n5387.n3 65.6672
R11938 a_6384_n5387.n0 a_6384_n5387.t2 65.0005
R11939 a_6384_n5387.n0 a_6384_n5387.t0 45.0005
R11940 a_6947_n5258.n1 a_6947_n5258.n0 926.024
R11941 a_6947_n5258.t0 a_6947_n5258.n1 82.0838
R11942 a_6947_n5258.n0 a_6947_n5258.t1 63.3338
R11943 a_6947_n5258.n1 a_6947_n5258.t2 63.3219
R11944 a_6947_n5258.n0 a_6947_n5258.t3 29.7268
R11945 a_n1097_3557.t1 a_n1097_3557.t0 198.571
R11946 a_2671_3557.n3 a_2671_3557.n2 674.338
R11947 a_2671_3557.n1 a_2671_3557.t4 332.58
R11948 a_2671_3557.n2 a_2671_3557.n0 284.012
R11949 a_2671_3557.n2 a_2671_3557.n1 253.648
R11950 a_2671_3557.n1 a_2671_3557.t5 168.701
R11951 a_2671_3557.t0 a_2671_3557.n3 96.1553
R11952 a_2671_3557.n3 a_2671_3557.t2 65.6672
R11953 a_2671_3557.n0 a_2671_3557.t1 65.0005
R11954 a_2671_3557.n0 a_2671_3557.t3 45.0005
R11955 a_3692_n5650.n5 a_3692_n5650.n4 807.871
R11956 a_3692_n5650.n0 a_3692_n5650.t3 389.183
R11957 a_3692_n5650.n1 a_3692_n5650.n0 251.167
R11958 a_3692_n5650.n1 a_3692_n5650.t1 223.571
R11959 a_3692_n5650.n3 a_3692_n5650.t8 212.081
R11960 a_3692_n5650.n2 a_3692_n5650.t6 212.081
R11961 a_3692_n5650.n4 a_3692_n5650.n3 176.576
R11962 a_3692_n5650.n0 a_3692_n5650.t7 174.891
R11963 a_3692_n5650.n3 a_3692_n5650.t5 139.78
R11964 a_3692_n5650.n2 a_3692_n5650.t4 139.78
R11965 a_3692_n5650.t0 a_3692_n5650.n5 63.3219
R11966 a_3692_n5650.n5 a_3692_n5650.t2 63.3219
R11967 a_3692_n5650.n3 a_3692_n5650.n2 61.346
R11968 a_3692_n5650.n4 a_3692_n5650.n1 37.5061
R11969 CF[9].n11 CF[9].n10 585
R11970 CF[9].n12 CF[9].n11 585
R11971 CF[9].n6 CF[9].t6 333.651
R11972 CF[9].n6 CF[9].t8 297.233
R11973 CF[9].n3 CF[9].t4 294.557
R11974 CF[9].n0 CF[9].t5 294.557
R11975 CF[9].n3 CF[9].t9 211.01
R11976 CF[9].n0 CF[9].t7 211.01
R11977 CF[9].n7 CF[9].n6 196.493
R11978 CF[9].n9 CF[9].n8 185
R11979 CF[9].n4 CF[9].n3 153.097
R11980 CF[9].n1 CF[9].n0 152
R11981 CF[9] CF[9].n9 49.0339
R11982 CF[9] CF[9].n14 37.5283
R11983 CF[9].n14 CF[9] 36.2072
R11984 CF[9].n13 CF[9].n7 35.37
R11985 CF[9].n11 CF[9].t2 26.5955
R11986 CF[9].n11 CF[9].t3 26.5955
R11987 CF[9].n8 CF[9].t0 24.9236
R11988 CF[9].n8 CF[9].t1 24.9236
R11989 CF[9].n13 CF[9].n12 17.3072
R11990 CF[9].n10 CF[9] 15.6165
R11991 CF[9].n5 CF[9].n2 14.9321
R11992 CF[9].n5 CF[9].n4 13.9063
R11993 CF[9].n9 CF[9] 10.4965
R11994 CF[9].n2 CF[9] 9.32621
R11995 CF[9].n14 CF[9] 5.46175
R11996 CF[9].n4 CF[9] 3.10907
R11997 CF[9].n1 CF[9] 2.01193
R11998 CF[9].n12 CF[9] 1.7925
R11999 CF[9].n10 CF[9] 1.7925
R12000 CF[9].n2 CF[9].n1 1.09764
R12001 CF[9] CF[9].n5 0.847483
R12002 CF[9] CF[9].n13 0.745692
R12003 CF[9].n7 CF[9] 0.24431
R12004 a_n628_3557.n3 a_n628_3557.n2 636.953
R12005 a_n628_3557.n1 a_n628_3557.t4 366.856
R12006 a_n628_3557.n2 a_n628_3557.n0 300.2
R12007 a_n628_3557.n2 a_n628_3557.n1 225.036
R12008 a_n628_3557.n1 a_n628_3557.t5 174.056
R12009 a_n628_3557.n0 a_n628_3557.t1 70.0005
R12010 a_n628_3557.n3 a_n628_3557.t3 68.0124
R12011 a_n628_3557.t0 a_n628_3557.n3 63.3219
R12012 a_n628_3557.n0 a_n628_3557.t2 61.6672
R12013 a_8577_n4702.n3 a_8577_n4702.n2 636.953
R12014 a_8577_n4702.n1 a_8577_n4702.t4 366.856
R12015 a_8577_n4702.n2 a_8577_n4702.n0 300.2
R12016 a_8577_n4702.n2 a_8577_n4702.n1 225.036
R12017 a_8577_n4702.n1 a_8577_n4702.t5 174.056
R12018 a_8577_n4702.n0 a_8577_n4702.t3 70.0005
R12019 a_8577_n4702.t1 a_8577_n4702.n3 68.0124
R12020 a_8577_n4702.n3 a_8577_n4702.t2 63.3219
R12021 a_8577_n4702.n0 a_8577_n4702.t0 61.6672
R12022 a_8931_n4714.t0 a_8931_n4714.t1 87.1434
R12023 a_8752_n4776.n5 a_8752_n4776.n4 807.871
R12024 a_8752_n4776.n2 a_8752_n4776.t3 389.183
R12025 a_8752_n4776.n3 a_8752_n4776.n2 251.167
R12026 a_8752_n4776.n3 a_8752_n4776.t2 223.571
R12027 a_8752_n4776.n0 a_8752_n4776.t7 212.081
R12028 a_8752_n4776.n1 a_8752_n4776.t8 212.081
R12029 a_8752_n4776.n4 a_8752_n4776.n1 176.576
R12030 a_8752_n4776.n2 a_8752_n4776.t5 174.891
R12031 a_8752_n4776.n0 a_8752_n4776.t4 139.78
R12032 a_8752_n4776.n1 a_8752_n4776.t6 139.78
R12033 a_8752_n4776.n5 a_8752_n4776.t1 63.3219
R12034 a_8752_n4776.t0 a_8752_n4776.n5 63.3219
R12035 a_8752_n4776.n1 a_8752_n4776.n0 61.346
R12036 a_8752_n4776.n4 a_8752_n4776.n3 37.7195
R12037 SWP[4].n0 SWP[4].t4 332.312
R12038 SWP[4].n0 SWP[4].t5 295.627
R12039 SWP[4].n4 SWP[4].n3 289.096
R12040 SWP[4] SWP[4].n0 196.004
R12041 SWP[4].n6 SWP[4].n5 185
R12042 SWP[4] SWP[4].n6 49.0339
R12043 SWP[4].n1 SWP[4] 41.1196
R12044 SWP[4].n2 SWP[4] 40.0305
R12045 SWP[4].n3 SWP[4].t2 26.5955
R12046 SWP[4].n3 SWP[4].t3 26.5955
R12047 SWP[4].n5 SWP[4].t0 24.9236
R12048 SWP[4].n5 SWP[4].t1 24.9236
R12049 SWP[4] SWP[4].n2 16.8044
R12050 SWP[4] SWP[4].n7 14.6049
R12051 SWP[4].n7 SWP[4] 13.0565
R12052 SWP[4].n2 SWP[4].n1 12.3917
R12053 SWP[4].n6 SWP[4] 10.4965
R12054 SWP[4] SWP[4].n4 9.48653
R12055 SWP[4].n4 SWP[4] 7.7181
R12056 SWP[4].n7 SWP[4] 4.3525
R12057 SWP[4].n1 SWP[4] 0.0034375
R12058 a_5015_n5258.n1 a_5015_n5258.n0 926.024
R12059 a_5015_n5258.n0 a_5015_n5258.t2 82.0838
R12060 a_5015_n5258.n1 a_5015_n5258.t3 63.3338
R12061 a_5015_n5258.n0 a_5015_n5258.t1 63.3219
R12062 a_5015_n5258.t0 a_5015_n5258.n1 29.7268
R12063 a_5343_3531.n5 a_5343_3531.n4 807.871
R12064 a_5343_3531.n2 a_5343_3531.t3 389.183
R12065 a_5343_3531.n3 a_5343_3531.n2 251.167
R12066 a_5343_3531.n3 a_5343_3531.t2 223.571
R12067 a_5343_3531.n0 a_5343_3531.t4 212.081
R12068 a_5343_3531.n1 a_5343_3531.t8 212.081
R12069 a_5343_3531.n4 a_5343_3531.n1 176.576
R12070 a_5343_3531.n2 a_5343_3531.t5 174.891
R12071 a_5343_3531.n0 a_5343_3531.t7 139.78
R12072 a_5343_3531.n1 a_5343_3531.t6 139.78
R12073 a_5343_3531.n5 a_5343_3531.t1 63.3219
R12074 a_5343_3531.t0 a_5343_3531.n5 63.3219
R12075 a_5343_3531.n1 a_5343_3531.n0 61.346
R12076 a_5343_3531.n4 a_5343_3531.n3 37.7195
R12077 auto_sampling_0.x24.A.n5 auto_sampling_0.x24.A.n4 244.069
R12078 auto_sampling_0.x24.A.n2 auto_sampling_0.x24.A.n0 236.589
R12079 auto_sampling_0.x24.A.n9 auto_sampling_0.x24.A.t13 212.081
R12080 auto_sampling_0.x24.A.n11 auto_sampling_0.x24.A.t17 212.081
R12081 auto_sampling_0.x24.A.n8 auto_sampling_0.x24.A.t21 212.081
R12082 auto_sampling_0.x24.A.n16 auto_sampling_0.x24.A.t11 212.081
R12083 auto_sampling_0.x24.A.n7 auto_sampling_0.x24.A.t23 212.081
R12084 auto_sampling_0.x24.A.n21 auto_sampling_0.x24.A.t18 212.081
R12085 auto_sampling_0.x24.A.n23 auto_sampling_0.x24.A.t9 212.081
R12086 auto_sampling_0.x24.A.n24 auto_sampling_0.x24.A.t15 212.081
R12087 auto_sampling_0.x24.A.n5 auto_sampling_0.x24.A.n3 204.892
R12088 auto_sampling_0.x24.A.n2 auto_sampling_0.x24.A.n1 200.321
R12089 auto_sampling_0.x24.A auto_sampling_0.x24.A.n25 163.264
R12090 auto_sampling_0.x24.A.n22 auto_sampling_0.x24.A.n6 152
R12091 auto_sampling_0.x24.A.n20 auto_sampling_0.x24.A.n19 152
R12092 auto_sampling_0.x24.A.n18 auto_sampling_0.x24.A.n17 152
R12093 auto_sampling_0.x24.A.n15 auto_sampling_0.x24.A.n14 152
R12094 auto_sampling_0.x24.A.n13 auto_sampling_0.x24.A.n12 152
R12095 auto_sampling_0.x24.A.n10 auto_sampling_0.x24.A 152
R12096 auto_sampling_0.x24.A.n9 auto_sampling_0.x24.A.t20 139.78
R12097 auto_sampling_0.x24.A.n11 auto_sampling_0.x24.A.t8 139.78
R12098 auto_sampling_0.x24.A.n8 auto_sampling_0.x24.A.t12 139.78
R12099 auto_sampling_0.x24.A.n16 auto_sampling_0.x24.A.t19 139.78
R12100 auto_sampling_0.x24.A.n7 auto_sampling_0.x24.A.t14 139.78
R12101 auto_sampling_0.x24.A.n21 auto_sampling_0.x24.A.t10 139.78
R12102 auto_sampling_0.x24.A.n23 auto_sampling_0.x24.A.t16 139.78
R12103 auto_sampling_0.x24.A.n24 auto_sampling_0.x24.A.t22 139.78
R12104 auto_sampling_0.x24.A.n10 auto_sampling_0.x24.A.n9 30.6732
R12105 auto_sampling_0.x24.A.n11 auto_sampling_0.x24.A.n10 30.6732
R12106 auto_sampling_0.x24.A.n12 auto_sampling_0.x24.A.n11 30.6732
R12107 auto_sampling_0.x24.A.n12 auto_sampling_0.x24.A.n8 30.6732
R12108 auto_sampling_0.x24.A.n15 auto_sampling_0.x24.A.n8 30.6732
R12109 auto_sampling_0.x24.A.n16 auto_sampling_0.x24.A.n15 30.6732
R12110 auto_sampling_0.x24.A.n17 auto_sampling_0.x24.A.n16 30.6732
R12111 auto_sampling_0.x24.A.n17 auto_sampling_0.x24.A.n7 30.6732
R12112 auto_sampling_0.x24.A.n20 auto_sampling_0.x24.A.n7 30.6732
R12113 auto_sampling_0.x24.A.n21 auto_sampling_0.x24.A.n20 30.6732
R12114 auto_sampling_0.x24.A.n22 auto_sampling_0.x24.A.n21 30.6732
R12115 auto_sampling_0.x24.A.n23 auto_sampling_0.x24.A.n22 30.6732
R12116 auto_sampling_0.x24.A.n25 auto_sampling_0.x24.A.n23 30.6732
R12117 auto_sampling_0.x24.A.n25 auto_sampling_0.x24.A.n24 30.6732
R12118 auto_sampling_0.x24.A.n4 auto_sampling_0.x24.A.t6 26.5955
R12119 auto_sampling_0.x24.A.n4 auto_sampling_0.x24.A.t5 26.5955
R12120 auto_sampling_0.x24.A.n3 auto_sampling_0.x24.A.t1 26.5955
R12121 auto_sampling_0.x24.A.n3 auto_sampling_0.x24.A.t3 26.5955
R12122 auto_sampling_0.x24.A.n0 auto_sampling_0.x24.A.t2 24.9236
R12123 auto_sampling_0.x24.A.n0 auto_sampling_0.x24.A.t0 24.9236
R12124 auto_sampling_0.x24.A.n1 auto_sampling_0.x24.A.t4 24.9236
R12125 auto_sampling_0.x24.A.n1 auto_sampling_0.x24.A.t7 24.9236
R12126 auto_sampling_0.x24.A.n13 auto_sampling_0.x24.A 21.5045
R12127 auto_sampling_0.x24.A.n27 auto_sampling_0.x24.A.n26 19.5596
R12128 auto_sampling_0.x24.A.n14 auto_sampling_0.x24.A 19.4565
R12129 auto_sampling_0.x24.A auto_sampling_0.x24.A.n5 18.4569
R12130 auto_sampling_0.x24.A.n18 auto_sampling_0.x24.A 17.4085
R12131 auto_sampling_0.x24.A.n19 auto_sampling_0.x24.A 15.3605
R12132 auto_sampling_0.x24.A.n28 auto_sampling_0.x24.A 14.008
R12133 auto_sampling_0.x24.A auto_sampling_0.x24.A.n6 13.3125
R12134 auto_sampling_0.x24.A.n27 auto_sampling_0.x24.A 12.3175
R12135 auto_sampling_0.x24.A.n28 auto_sampling_0.x24.A.n2 12.0894
R12136 auto_sampling_0.x24.A.n19 auto_sampling_0.x24.A 8.1925
R12137 auto_sampling_0.x24.A auto_sampling_0.x24.A.n18 6.1445
R12138 auto_sampling_0.x24.A.n26 auto_sampling_0.x24.A.n6 5.8885
R12139 auto_sampling_0.x24.A.n26 auto_sampling_0.x24.A 4.3525
R12140 auto_sampling_0.x24.A auto_sampling_0.x24.A.n27 4.10616
R12141 auto_sampling_0.x24.A.n14 auto_sampling_0.x24.A 4.0965
R12142 auto_sampling_0.x24.A auto_sampling_0.x24.A.n28 2.41559
R12143 auto_sampling_0.x24.A auto_sampling_0.x24.A.n13 2.0485
R12144 a_2888_2959.n3 a_2888_2959.n2 647.119
R12145 a_2888_2959.n1 a_2888_2959.t5 350.253
R12146 a_2888_2959.n2 a_2888_2959.n0 260.339
R12147 a_2888_2959.n2 a_2888_2959.n1 246.119
R12148 a_2888_2959.n1 a_2888_2959.t4 189.588
R12149 a_2888_2959.n3 a_2888_2959.t3 89.1195
R12150 a_2888_2959.n0 a_2888_2959.t0 63.3338
R12151 a_2888_2959.t2 a_2888_2959.n3 41.0422
R12152 a_2888_2959.n0 a_2888_2959.t1 31.9797
R12153 a_2778_3083.t0 a_2778_3083.n0 1327.82
R12154 a_2778_3083.n0 a_2778_3083.t2 194.655
R12155 a_2778_3083.n0 a_2778_3083.t1 63.3219
R12156 a_n8868_n9662.n1 a_n8868_n9662.n0 926.024
R12157 a_n8868_n9662.t1 a_n8868_n9662.n1 82.0838
R12158 a_n8868_n9662.n0 a_n8868_n9662.t0 63.3338
R12159 a_n8868_n9662.n1 a_n8868_n9662.t3 63.3219
R12160 a_n8868_n9662.n0 a_n8868_n9662.t2 29.7268
R12161 DOUT[5].n3 DOUT[5].n2 585
R12162 DOUT[5].n4 DOUT[5].n3 585
R12163 DOUT[5].n1 DOUT[5].n0 185
R12164 DOUT[5] DOUT[5].n1 57.7379
R12165 DOUT[5].n3 DOUT[5].t3 26.5955
R12166 DOUT[5].n3 DOUT[5].t2 26.5955
R12167 DOUT[5].n0 DOUT[5].t1 24.9236
R12168 DOUT[5].n0 DOUT[5].t0 24.9236
R12169 DOUT[5] DOUT[5].n5 17.8877
R12170 DOUT[5].n2 DOUT[5] 10.4965
R12171 DOUT[5].n4 DOUT[5] 10.4965
R12172 DOUT[5].n2 DOUT[5] 6.9125
R12173 DOUT[5].n5 DOUT[5] 4.3525
R12174 DOUT[5].n5 DOUT[5].n4 2.5605
R12175 DOUT[5].n1 DOUT[5] 1.7925
R12176 a_5987_n1029.n1 a_5987_n1029.t6 530.01
R12177 a_5987_n1029.t1 a_5987_n1029.n5 421.021
R12178 a_5987_n1029.n0 a_5987_n1029.t2 337.142
R12179 a_5987_n1029.n3 a_5987_n1029.t0 280.223
R12180 a_5987_n1029.n4 a_5987_n1029.t4 263.173
R12181 a_5987_n1029.n4 a_5987_n1029.t7 227.826
R12182 a_5987_n1029.n0 a_5987_n1029.t3 199.762
R12183 a_5987_n1029.n2 a_5987_n1029.n1 170.81
R12184 a_5987_n1029.n2 a_5987_n1029.n0 167.321
R12185 a_5987_n1029.n5 a_5987_n1029.n4 152
R12186 a_5987_n1029.n1 a_5987_n1029.t5 141.923
R12187 a_5987_n1029.n3 a_5987_n1029.n2 10.8376
R12188 a_5987_n1029.n5 a_5987_n1029.n3 2.50485
R12189 a_6721_n787.n3 a_6721_n787.n2 647.119
R12190 a_6721_n787.n1 a_6721_n787.t5 350.253
R12191 a_6721_n787.n2 a_6721_n787.n0 260.339
R12192 a_6721_n787.n2 a_6721_n787.n1 246.119
R12193 a_6721_n787.n1 a_6721_n787.t4 189.588
R12194 a_6721_n787.n3 a_6721_n787.t3 89.1195
R12195 a_6721_n787.n0 a_6721_n787.t2 63.3338
R12196 a_6721_n787.t1 a_6721_n787.n3 41.0422
R12197 a_6721_n787.n0 a_6721_n787.t0 31.9797
R12198 a_9206_2691.n5 a_9206_2691.n4 807.871
R12199 a_9206_2691.n2 a_9206_2691.t5 389.183
R12200 a_9206_2691.n3 a_9206_2691.n2 251.167
R12201 a_9206_2691.n3 a_9206_2691.t1 223.571
R12202 a_9206_2691.n0 a_9206_2691.t7 212.081
R12203 a_9206_2691.n1 a_9206_2691.t3 212.081
R12204 a_9206_2691.n4 a_9206_2691.n1 176.576
R12205 a_9206_2691.n2 a_9206_2691.t4 174.891
R12206 a_9206_2691.n0 a_9206_2691.t8 139.78
R12207 a_9206_2691.n1 a_9206_2691.t6 139.78
R12208 a_9206_2691.n5 a_9206_2691.t2 63.3219
R12209 a_9206_2691.t0 a_9206_2691.n5 63.3219
R12210 a_9206_2691.n1 a_9206_2691.n0 61.346
R12211 a_9206_2691.n4 a_9206_2691.n3 37.7195
R12212 auto_sampling_0.x21.Q.n4 auto_sampling_0.x21.Q.t4 333.651
R12213 auto_sampling_0.x21.Q.n4 auto_sampling_0.x21.Q.t5 297.233
R12214 auto_sampling_0.x21.Q.n3 auto_sampling_0.x21.Q.n2 289.096
R12215 auto_sampling_0.x21.Q auto_sampling_0.x21.Q.n4 194.062
R12216 auto_sampling_0.x21.Q.n1 auto_sampling_0.x21.Q.n0 185
R12217 auto_sampling_0.x21.Q.n5 auto_sampling_0.x21.Q 69.9921
R12218 auto_sampling_0.x21.Q auto_sampling_0.x21.Q.n1 49.0339
R12219 auto_sampling_0.x21.Q.n2 auto_sampling_0.x21.Q.t2 26.5955
R12220 auto_sampling_0.x21.Q.n2 auto_sampling_0.x21.Q.t3 26.5955
R12221 auto_sampling_0.x21.Q.n0 auto_sampling_0.x21.Q.t0 24.9236
R12222 auto_sampling_0.x21.Q.n0 auto_sampling_0.x21.Q.t1 24.9236
R12223 auto_sampling_0.x21.Q.n5 auto_sampling_0.x21.Q 13.0565
R12224 auto_sampling_0.x21.Q.n1 auto_sampling_0.x21.Q 10.4965
R12225 auto_sampling_0.x21.Q auto_sampling_0.x21.Q.n3 9.48653
R12226 auto_sampling_0.x21.Q.n3 auto_sampling_0.x21.Q 7.7181
R12227 auto_sampling_0.x21.Q auto_sampling_0.x21.Q.n5 4.3525
R12228 a_4864_2717.t0 a_4864_2717.t1 60.0005
R12229 a_815_n663.n0 a_815_n663.t2 1327.82
R12230 a_815_n663.t0 a_815_n663.n0 194.655
R12231 a_815_n663.n0 a_815_n663.t1 63.3219
R12232 auto_sampling_0.x5.D.n5 auto_sampling_0.x5.D.n4 585
R12233 auto_sampling_0.x5.D.n4 auto_sampling_0.x5.D.n3 585
R12234 auto_sampling_0.x5.D.n2 auto_sampling_0.x5.D.t5 333.651
R12235 auto_sampling_0.x5.D.n2 auto_sampling_0.x5.D.t4 297.233
R12236 auto_sampling_0.x5.D auto_sampling_0.x5.D.n2 196.493
R12237 auto_sampling_0.x5.D.n1 auto_sampling_0.x5.D.n0 185
R12238 auto_sampling_0.x5.D auto_sampling_0.x5.D.n1 49.0339
R12239 auto_sampling_0.x5.D.n3 auto_sampling_0.x5.D 44.2533
R12240 auto_sampling_0.x5.D.n4 auto_sampling_0.x5.D.t3 26.5955
R12241 auto_sampling_0.x5.D.n4 auto_sampling_0.x5.D.t2 26.5955
R12242 auto_sampling_0.x5.D.n0 auto_sampling_0.x5.D.t0 24.9236
R12243 auto_sampling_0.x5.D.n0 auto_sampling_0.x5.D.t1 24.9236
R12244 auto_sampling_0.x5.D.n5 auto_sampling_0.x5.D 15.6165
R12245 auto_sampling_0.x5.D.n1 auto_sampling_0.x5.D 10.4965
R12246 auto_sampling_0.x5.D.n3 auto_sampling_0.x5.D 1.7925
R12247 auto_sampling_0.x5.D auto_sampling_0.x5.D.n5 1.7925
R12248 a_6440_3557.n1 a_6440_3557.n0 926.024
R12249 a_6440_3557.t1 a_6440_3557.n1 82.0838
R12250 a_6440_3557.n0 a_6440_3557.t0 63.3338
R12251 a_6440_3557.n1 a_6440_3557.t3 63.3219
R12252 a_6440_3557.n0 a_6440_3557.t2 29.7268
R12253 a_n7357_n9484.n1 a_n7357_n9484.t3 530.01
R12254 a_n7357_n9484.t0 a_n7357_n9484.n5 421.021
R12255 a_n7357_n9484.n0 a_n7357_n9484.t4 337.142
R12256 a_n7357_n9484.n3 a_n7357_n9484.t1 280.223
R12257 a_n7357_n9484.n4 a_n7357_n9484.t6 263.173
R12258 a_n7357_n9484.n4 a_n7357_n9484.t7 227.826
R12259 a_n7357_n9484.n0 a_n7357_n9484.t5 199.762
R12260 a_n7357_n9484.n2 a_n7357_n9484.n1 170.81
R12261 a_n7357_n9484.n2 a_n7357_n9484.n0 167.321
R12262 a_n7357_n9484.n5 a_n7357_n9484.n4 152
R12263 a_n7357_n9484.n1 a_n7357_n9484.t2 141.923
R12264 a_n7357_n9484.n3 a_n7357_n9484.n2 10.8376
R12265 a_n7357_n9484.n5 a_n7357_n9484.n3 2.50485
R12266 a_n6936_n9484.n1 a_n6936_n9484.n0 926.024
R12267 a_n6936_n9484.t0 a_n6936_n9484.n1 82.0838
R12268 a_n6936_n9484.n0 a_n6936_n9484.t1 63.3338
R12269 a_n6936_n9484.n1 a_n6936_n9484.t2 63.3219
R12270 a_n6936_n9484.n0 a_n6936_n9484.t3 29.7268
R12271 a_n6841_n9484.n3 a_n6841_n9484.n2 674.338
R12272 a_n6841_n9484.n1 a_n6841_n9484.t4 332.58
R12273 a_n6841_n9484.n2 a_n6841_n9484.n0 284.012
R12274 a_n6841_n9484.n2 a_n6841_n9484.n1 253.648
R12275 a_n6841_n9484.n1 a_n6841_n9484.t5 168.701
R12276 a_n6841_n9484.n3 a_n6841_n9484.t1 96.1553
R12277 a_n6841_n9484.t0 a_n6841_n9484.n3 65.6672
R12278 a_n6841_n9484.n0 a_n6841_n9484.t2 65.0005
R12279 a_n6841_n9484.n0 a_n6841_n9484.t3 45.0005
R12280 a_8012_n4702.n3 a_8012_n4702.n2 674.338
R12281 a_8012_n4702.n1 a_8012_n4702.t5 332.58
R12282 a_8012_n4702.n2 a_8012_n4702.n0 284.012
R12283 a_8012_n4702.n2 a_8012_n4702.n1 253.648
R12284 a_8012_n4702.n1 a_8012_n4702.t4 168.701
R12285 a_8012_n4702.t0 a_8012_n4702.n3 96.1553
R12286 a_8012_n4702.n3 a_8012_n4702.t3 65.6672
R12287 a_8012_n4702.n0 a_8012_n4702.t2 65.0005
R12288 a_8012_n4702.n0 a_8012_n4702.t1 45.0005
R12289 a_8230_n5106.n3 a_8230_n5106.n2 647.119
R12290 a_8230_n5106.n1 a_8230_n5106.t4 350.253
R12291 a_8230_n5106.n2 a_8230_n5106.n0 260.339
R12292 a_8230_n5106.n2 a_8230_n5106.n1 246.119
R12293 a_8230_n5106.n1 a_8230_n5106.t5 189.588
R12294 a_8230_n5106.n3 a_8230_n5106.t0 89.1195
R12295 a_8230_n5106.n0 a_8230_n5106.t1 63.3338
R12296 a_8230_n5106.t3 a_8230_n5106.n3 41.0422
R12297 a_8230_n5106.n0 a_8230_n5106.t2 31.9797
R12298 a_2505_n1207.t0 a_2505_n1207.t1 87.1434
R12299 a_4969_n10054.n3 a_4969_n10054.n2 647.119
R12300 a_4969_n10054.n1 a_4969_n10054.t5 350.253
R12301 a_4969_n10054.n2 a_4969_n10054.n0 260.339
R12302 a_4969_n10054.n2 a_4969_n10054.n1 246.119
R12303 a_4969_n10054.n1 a_4969_n10054.t4 189.588
R12304 a_4969_n10054.n3 a_4969_n10054.t0 89.1195
R12305 a_4969_n10054.n0 a_4969_n10054.t2 63.3338
R12306 a_4969_n10054.t1 a_4969_n10054.n3 41.0422
R12307 a_4969_n10054.n0 a_4969_n10054.t3 31.9797
R12308 a_4859_n10028.n0 a_4859_n10028.t2 1327.82
R12309 a_4859_n10028.t0 a_4859_n10028.n0 194.655
R12310 a_4859_n10028.n0 a_4859_n10028.t1 63.3219
R12311 a_n6733_n9118.n0 a_n6733_n9118.t1 1327.82
R12312 a_n6733_n9118.t0 a_n6733_n9118.n0 194.655
R12313 a_n6733_n9118.n0 a_n6733_n9118.t2 63.3219
R12314 a_2364_n5482.n1 a_2364_n5482.t2 530.01
R12315 a_2364_n5482.t0 a_2364_n5482.n5 421.021
R12316 a_2364_n5482.n0 a_2364_n5482.t3 337.171
R12317 a_2364_n5482.n3 a_2364_n5482.t1 280.223
R12318 a_2364_n5482.n4 a_2364_n5482.t5 263.173
R12319 a_2364_n5482.n4 a_2364_n5482.t6 227.826
R12320 a_2364_n5482.n0 a_2364_n5482.t4 199.762
R12321 a_2364_n5482.n2 a_2364_n5482.n1 170.81
R12322 a_2364_n5482.n2 a_2364_n5482.n0 167.321
R12323 a_2364_n5482.n5 a_2364_n5482.n4 152
R12324 a_2364_n5482.n1 a_2364_n5482.t7 141.923
R12325 a_2364_n5482.n3 a_2364_n5482.n2 10.8376
R12326 a_2364_n5482.n5 a_2364_n5482.n3 2.50485
R12327 a_2665_n5258.t0 a_2665_n5258.n0 1327.82
R12328 a_2665_n5258.n0 a_2665_n5258.t2 194.655
R12329 a_2665_n5258.n0 a_2665_n5258.t1 63.3219
R12330 a_2520_n5387.n3 a_2520_n5387.n2 674.338
R12331 a_2520_n5387.n1 a_2520_n5387.t4 332.58
R12332 a_2520_n5387.n2 a_2520_n5387.n0 284.012
R12333 a_2520_n5387.n2 a_2520_n5387.n1 253.648
R12334 a_2520_n5387.n1 a_2520_n5387.t5 168.701
R12335 a_2520_n5387.t1 a_2520_n5387.n3 96.1553
R12336 a_2520_n5387.n3 a_2520_n5387.t3 65.6672
R12337 a_2520_n5387.n0 a_2520_n5387.t0 65.0005
R12338 a_2520_n5387.n0 a_2520_n5387.t2 45.0005
R12339 a_n2759_n10054.n3 a_n2759_n10054.n2 647.119
R12340 a_n2759_n10054.n1 a_n2759_n10054.t4 350.253
R12341 a_n2759_n10054.n2 a_n2759_n10054.n0 260.339
R12342 a_n2759_n10054.n2 a_n2759_n10054.n1 246.119
R12343 a_n2759_n10054.n1 a_n2759_n10054.t5 189.588
R12344 a_n2759_n10054.n3 a_n2759_n10054.t2 89.1195
R12345 a_n2759_n10054.n0 a_n2759_n10054.t3 63.3338
R12346 a_n2759_n10054.t1 a_n2759_n10054.n3 41.0422
R12347 a_n2759_n10054.n0 a_n2759_n10054.t0 31.9797
R12348 a_n2881_n9650.t1 a_n2881_n9650.t0 198.571
R12349 a_n7357_n10022.n1 a_n7357_n10022.t5 530.01
R12350 a_n7357_n10022.t1 a_n7357_n10022.n5 421.021
R12351 a_n7357_n10022.n0 a_n7357_n10022.t4 337.142
R12352 a_n7357_n10022.n3 a_n7357_n10022.t0 280.223
R12353 a_n7357_n10022.n4 a_n7357_n10022.t7 263.173
R12354 a_n7357_n10022.n4 a_n7357_n10022.t3 227.826
R12355 a_n7357_n10022.n0 a_n7357_n10022.t2 199.762
R12356 a_n7357_n10022.n2 a_n7357_n10022.n1 170.81
R12357 a_n7357_n10022.n2 a_n7357_n10022.n0 167.321
R12358 a_n7357_n10022.n5 a_n7357_n10022.n4 152
R12359 a_n7357_n10022.n1 a_n7357_n10022.t6 141.923
R12360 a_n7357_n10022.n3 a_n7357_n10022.n2 10.8376
R12361 a_n7357_n10022.n5 a_n7357_n10022.n3 2.50485
R12362 a_n6276_n9650.n3 a_n6276_n9650.n2 636.953
R12363 a_n6276_n9650.n1 a_n6276_n9650.t5 366.856
R12364 a_n6276_n9650.n2 a_n6276_n9650.n0 300.2
R12365 a_n6276_n9650.n2 a_n6276_n9650.n1 225.036
R12366 a_n6276_n9650.n1 a_n6276_n9650.t4 174.056
R12367 a_n6276_n9650.n0 a_n6276_n9650.t0 70.0005
R12368 a_n6276_n9650.n3 a_n6276_n9650.t2 68.0124
R12369 a_n6276_n9650.t1 a_n6276_n9650.n3 63.3219
R12370 a_n6276_n9650.n0 a_n6276_n9650.t3 61.6672
R12371 a_n6167_n9650.n0 a_n6167_n9650.t1 68.3338
R12372 a_n6167_n9650.n0 a_n6167_n9650.t0 26.3935
R12373 a_n6167_n9650.n1 a_n6167_n9650.n0 14.4005
R12374 a_6901_n10054.n3 a_6901_n10054.n2 647.119
R12375 a_6901_n10054.n1 a_6901_n10054.t4 350.253
R12376 a_6901_n10054.n2 a_6901_n10054.n0 260.339
R12377 a_6901_n10054.n2 a_6901_n10054.n1 246.119
R12378 a_6901_n10054.n1 a_6901_n10054.t5 189.588
R12379 a_6901_n10054.n3 a_6901_n10054.t0 89.1195
R12380 a_6901_n10054.n0 a_6901_n10054.t1 63.3338
R12381 a_6901_n10054.t3 a_6901_n10054.n3 41.0422
R12382 a_6901_n10054.n0 a_6901_n10054.t2 31.9797
R12383 a_6779_n9650.t0 a_6779_n9650.t1 198.571
R12384 a_6945_n9662.t0 a_6945_n9662.t1 60.0005
R12385 a_2434_n5106.n3 a_2434_n5106.n2 647.119
R12386 a_2434_n5106.n1 a_2434_n5106.t4 350.253
R12387 a_2434_n5106.n2 a_2434_n5106.n0 260.339
R12388 a_2434_n5106.n2 a_2434_n5106.n1 246.119
R12389 a_2434_n5106.n1 a_2434_n5106.t5 189.588
R12390 a_2434_n5106.n3 a_2434_n5106.t2 89.1195
R12391 a_2434_n5106.n0 a_2434_n5106.t1 63.3338
R12392 a_2434_n5106.t3 a_2434_n5106.n3 41.0422
R12393 a_2434_n5106.n0 a_2434_n5106.t0 31.9797
R12394 a_2312_n4702.t0 a_2312_n4702.t1 198.571
R12395 a_2478_n4714.t0 a_2478_n4714.t1 60.0005
R12396 a_n6101_n9724.n4 a_n6101_n9724.n1 807.871
R12397 a_n6101_n9724.n0 a_n6101_n9724.t4 389.183
R12398 a_n6101_n9724.n5 a_n6101_n9724.n0 251.167
R12399 a_n6101_n9724.t0 a_n6101_n9724.n5 223.571
R12400 a_n6101_n9724.n2 a_n6101_n9724.t7 212.081
R12401 a_n6101_n9724.n3 a_n6101_n9724.t5 212.081
R12402 a_n6101_n9724.n4 a_n6101_n9724.n3 176.576
R12403 a_n6101_n9724.n0 a_n6101_n9724.t6 174.891
R12404 a_n6101_n9724.n2 a_n6101_n9724.t3 139.78
R12405 a_n6101_n9724.n3 a_n6101_n9724.t8 139.78
R12406 a_n6101_n9724.n1 a_n6101_n9724.t1 63.3219
R12407 a_n6101_n9724.n1 a_n6101_n9724.t2 63.3219
R12408 a_n6101_n9724.n3 a_n6101_n9724.n2 61.346
R12409 a_n6101_n9724.n5 a_n6101_n9724.n4 37.7195
R12410 SWN[1].n4 SWN[1].n3 585
R12411 SWN[1].n3 SWN[1].n2 585
R12412 SWN[1].n1 SWN[1].n0 185
R12413 SWN[1].n5 SWN[1].n1 53.3859
R12414 SWN[1].n3 SWN[1].t2 26.5955
R12415 SWN[1].n3 SWN[1].t3 26.5955
R12416 SWN[1].n0 SWN[1].t1 24.9236
R12417 SWN[1].n0 SWN[1].t0 24.9236
R12418 SWN[1] SWN[1].n5 14.676
R12419 SWN[1] SWN[1].n4 10.4965
R12420 SWN[1].n2 SWN[1] 10.4965
R12421 SWN[1].n4 SWN[1] 6.9125
R12422 SWN[1].n2 SWN[1] 6.9125
R12423 SWN[1].n5 SWN[1] 4.3525
R12424 SWN[1].n1 SWN[1] 1.7925
R12425 a_4221_n1029.t1 a_4221_n1029.n3 370.026
R12426 a_4221_n1029.n0 a_4221_n1029.t5 351.356
R12427 a_4221_n1029.n1 a_4221_n1029.t2 334.717
R12428 a_4221_n1029.n3 a_4221_n1029.t0 325.971
R12429 a_4221_n1029.n1 a_4221_n1029.t3 309.935
R12430 a_4221_n1029.n0 a_4221_n1029.t4 305.683
R12431 a_4221_n1029.n2 a_4221_n1029.n0 16.879
R12432 a_4221_n1029.n3 a_4221_n1029.n2 10.8867
R12433 a_4221_n1029.n2 a_4221_n1029.n1 9.3005
R12434 a_4571_n1029.n3 a_4571_n1029.n2 674.338
R12435 a_4571_n1029.n1 a_4571_n1029.t5 332.58
R12436 a_4571_n1029.n2 a_4571_n1029.n0 284.012
R12437 a_4571_n1029.n2 a_4571_n1029.n1 253.648
R12438 a_4571_n1029.n1 a_4571_n1029.t4 168.701
R12439 a_4571_n1029.n3 a_4571_n1029.t3 96.1553
R12440 a_4571_n1029.t0 a_4571_n1029.n3 65.6672
R12441 a_4571_n1029.n0 a_4571_n1029.t2 65.0005
R12442 a_4571_n1029.n0 a_4571_n1029.t1 45.0005
R12443 a_4667_n1029.t1 a_4667_n1029.t0 198.571
R12444 a_8099_n9484.n1 a_8099_n9484.t7 530.01
R12445 a_8099_n9484.t1 a_8099_n9484.n5 421.021
R12446 a_8099_n9484.n0 a_8099_n9484.t2 337.142
R12447 a_8099_n9484.n3 a_8099_n9484.t0 280.223
R12448 a_8099_n9484.n4 a_8099_n9484.t5 263.173
R12449 a_8099_n9484.n4 a_8099_n9484.t6 227.826
R12450 a_8099_n9484.n0 a_8099_n9484.t3 199.762
R12451 a_8099_n9484.n2 a_8099_n9484.n1 170.81
R12452 a_8099_n9484.n2 a_8099_n9484.n0 167.321
R12453 a_8099_n9484.n5 a_8099_n9484.n4 152
R12454 a_8099_n9484.n1 a_8099_n9484.t4 141.923
R12455 a_8099_n9484.n3 a_8099_n9484.n2 10.8376
R12456 a_8099_n9484.n5 a_8099_n9484.n3 2.50485
R12457 a_8833_n9242.n3 a_8833_n9242.n2 647.119
R12458 a_8833_n9242.n1 a_8833_n9242.t5 350.253
R12459 a_8833_n9242.n2 a_8833_n9242.n0 260.339
R12460 a_8833_n9242.n2 a_8833_n9242.n1 246.119
R12461 a_8833_n9242.n1 a_8833_n9242.t4 189.588
R12462 a_8833_n9242.n3 a_8833_n9242.t1 89.1195
R12463 a_8833_n9242.n0 a_8833_n9242.t0 63.3338
R12464 a_8833_n9242.t3 a_8833_n9242.n3 41.0422
R12465 a_8833_n9242.n0 a_8833_n9242.t2 31.9797
R12466 a_9180_n9484.n3 a_9180_n9484.n2 636.953
R12467 a_9180_n9484.n1 a_9180_n9484.t4 366.856
R12468 a_9180_n9484.n2 a_9180_n9484.n0 300.2
R12469 a_9180_n9484.n2 a_9180_n9484.n1 225.036
R12470 a_9180_n9484.n1 a_9180_n9484.t5 174.056
R12471 a_9180_n9484.n0 a_9180_n9484.t0 70.0005
R12472 a_9180_n9484.t1 a_9180_n9484.n3 68.0124
R12473 a_9180_n9484.n3 a_9180_n9484.t3 63.3219
R12474 a_9180_n9484.n0 a_9180_n9484.t2 61.6672
R12475 a_n4691_n9242.n3 a_n4691_n9242.n2 647.119
R12476 a_n4691_n9242.n1 a_n4691_n9242.t5 350.253
R12477 a_n4691_n9242.n2 a_n4691_n9242.n0 260.339
R12478 a_n4691_n9242.n2 a_n4691_n9242.n1 246.119
R12479 a_n4691_n9242.n1 a_n4691_n9242.t4 189.588
R12480 a_n4691_n9242.n3 a_n4691_n9242.t3 89.1195
R12481 a_n4691_n9242.n0 a_n4691_n9242.t0 63.3338
R12482 a_n4691_n9242.t1 a_n4691_n9242.n3 41.0422
R12483 a_n4691_n9242.n0 a_n4691_n9242.t2 31.9797
R12484 a_n4801_n9118.n0 a_n4801_n9118.t2 1327.82
R12485 a_n4801_n9118.n0 a_n4801_n9118.t1 194.655
R12486 a_n4801_n9118.t0 a_n4801_n9118.n0 63.3219
R12487 a_9661_n5596.t0 a_9661_n5596.t1 77.1434
R12488 a_9487_n5472.n2 a_9487_n5472.n0 672.948
R12489 a_9487_n5472.t0 a_9487_n5472.n2 314.563
R12490 a_9487_n5472.n1 a_9487_n5472.t4 236.18
R12491 a_9487_n5472.n1 a_9487_n5472.t3 163.881
R12492 a_9487_n5472.n2 a_9487_n5472.n1 152
R12493 a_9487_n5472.n0 a_9487_n5472.t1 63.3219
R12494 a_9487_n5472.n0 a_9487_n5472.t2 63.3219
R12495 a_3379_n1055.n5 a_3379_n1055.n4 807.871
R12496 a_3379_n1055.n2 a_3379_n1055.t6 389.183
R12497 a_3379_n1055.n3 a_3379_n1055.n2 251.167
R12498 a_3379_n1055.n3 a_3379_n1055.t1 223.571
R12499 a_3379_n1055.n0 a_3379_n1055.t7 212.081
R12500 a_3379_n1055.n1 a_3379_n1055.t4 212.081
R12501 a_3379_n1055.n4 a_3379_n1055.n1 176.576
R12502 a_3379_n1055.n2 a_3379_n1055.t8 174.891
R12503 a_3379_n1055.n0 a_3379_n1055.t3 139.78
R12504 a_3379_n1055.n1 a_3379_n1055.t5 139.78
R12505 a_3379_n1055.t0 a_3379_n1055.n5 63.3219
R12506 a_3379_n1055.n5 a_3379_n1055.t2 63.3219
R12507 a_3379_n1055.n1 a_3379_n1055.n0 61.346
R12508 a_3379_n1055.n4 a_3379_n1055.n3 37.7195
R12509 a_6334_n1441.n3 a_6334_n1441.n2 636.953
R12510 a_6334_n1441.n1 a_6334_n1441.t5 366.856
R12511 a_6334_n1441.n2 a_6334_n1441.n0 300.2
R12512 a_6334_n1441.n2 a_6334_n1441.n1 225.036
R12513 a_6334_n1441.n1 a_6334_n1441.t4 174.056
R12514 a_6334_n1441.n0 a_6334_n1441.t2 70.0005
R12515 a_6334_n1441.t0 a_6334_n1441.n3 68.0124
R12516 a_6334_n1441.n3 a_6334_n1441.t1 63.3219
R12517 a_6334_n1441.n0 a_6334_n1441.t3 61.6672
R12518 SWP[8].n0 SWP[8].t5 332.312
R12519 SWP[8].n0 SWP[8].t4 295.627
R12520 SWP[8].n4 SWP[8].n3 289.096
R12521 SWP[8] SWP[8].n0 196.004
R12522 SWP[8].n6 SWP[8].n5 185
R12523 SWP[8] SWP[8].n6 49.0339
R12524 SWP[8].n1 SWP[8] 41.1194
R12525 SWP[8].n2 SWP[8] 30.6188
R12526 SWP[8].n3 SWP[8].t3 26.5955
R12527 SWP[8].n3 SWP[8].t1 26.5955
R12528 SWP[8].n5 SWP[8].t2 24.9236
R12529 SWP[8].n5 SWP[8].t0 24.9236
R12530 SWP[8] SWP[8].n7 14.6049
R12531 SWP[8].n2 SWP[8].n1 13.4647
R12532 SWP[8].n7 SWP[8] 13.0565
R12533 SWP[8].n6 SWP[8] 10.4965
R12534 SWP[8] SWP[8].n4 9.48653
R12535 SWP[8].n4 SWP[8] 7.7181
R12536 SWP[8] SWP[8].n2 7.36911
R12537 SWP[8].n7 SWP[8] 4.3525
R12538 SWP[8].n1 SWP[8] 0.00285
R12539 a_8879_n5258.n1 a_8879_n5258.n0 926.024
R12540 a_8879_n5258.n0 a_8879_n5258.t2 82.0838
R12541 a_8879_n5258.n1 a_8879_n5258.t3 63.3338
R12542 a_8879_n5258.n0 a_8879_n5258.t1 63.3219
R12543 a_8879_n5258.t0 a_8879_n5258.n1 29.7268
R12544 a_7100_3557.n3 a_7100_3557.n2 636.953
R12545 a_7100_3557.n1 a_7100_3557.t4 366.856
R12546 a_7100_3557.n2 a_7100_3557.n0 300.2
R12547 a_7100_3557.n2 a_7100_3557.n1 225.036
R12548 a_7100_3557.n1 a_7100_3557.t5 174.056
R12549 a_7100_3557.n0 a_7100_3557.t2 70.0005
R12550 a_7100_3557.n3 a_7100_3557.t3 68.0124
R12551 a_7100_3557.t1 a_7100_3557.n3 63.3219
R12552 a_7100_3557.n0 a_7100_3557.t0 61.6672
R12553 a_7454_3557.t0 a_7454_3557.t1 87.1434
R12554 a_7275_3531.n5 a_7275_3531.n4 807.871
R12555 a_7275_3531.n2 a_7275_3531.t5 389.183
R12556 a_7275_3531.n3 a_7275_3531.n2 251.167
R12557 a_7275_3531.n3 a_7275_3531.t1 223.571
R12558 a_7275_3531.n0 a_7275_3531.t6 212.081
R12559 a_7275_3531.n1 a_7275_3531.t4 212.081
R12560 a_7275_3531.n4 a_7275_3531.n1 176.576
R12561 a_7275_3531.n2 a_7275_3531.t8 174.891
R12562 a_7275_3531.n0 a_7275_3531.t3 139.78
R12563 a_7275_3531.n1 a_7275_3531.t7 139.78
R12564 a_7275_3531.n5 a_7275_3531.t2 63.3219
R12565 a_7275_3531.t0 a_7275_3531.n5 63.3219
R12566 a_7275_3531.n1 a_7275_3531.n0 61.346
R12567 a_7275_3531.n4 a_7275_3531.n3 37.7195
R12568 a_5298_n663.t0 a_5298_n663.t1 126.644
R12569 a_n2237_n9510.n3 a_n2237_n9510.n0 807.871
R12570 a_n2237_n9510.n4 a_n2237_n9510.t3 389.183
R12571 a_n2237_n9510.n5 a_n2237_n9510.n4 251.167
R12572 a_n2237_n9510.t0 a_n2237_n9510.n5 223.571
R12573 a_n2237_n9510.n1 a_n2237_n9510.t7 212.081
R12574 a_n2237_n9510.n2 a_n2237_n9510.t5 212.081
R12575 a_n2237_n9510.n3 a_n2237_n9510.n2 176.576
R12576 a_n2237_n9510.n4 a_n2237_n9510.t8 174.891
R12577 a_n2237_n9510.n1 a_n2237_n9510.t6 139.78
R12578 a_n2237_n9510.n2 a_n2237_n9510.t4 139.78
R12579 a_n2237_n9510.n0 a_n2237_n9510.t1 63.3219
R12580 a_n2237_n9510.n0 a_n2237_n9510.t2 63.3219
R12581 a_n2237_n9510.n2 a_n2237_n9510.n1 61.346
R12582 a_n2237_n9510.n5 a_n2237_n9510.n3 37.7195
R12583 a_n2250_n9118.t0 a_n2250_n9118.t1 126.644
R12584 a_3411_3531.n5 a_3411_3531.n4 807.871
R12585 a_3411_3531.n2 a_3411_3531.t4 389.183
R12586 a_3411_3531.n3 a_3411_3531.n2 251.167
R12587 a_3411_3531.n3 a_3411_3531.t1 223.571
R12588 a_3411_3531.n0 a_3411_3531.t6 212.081
R12589 a_3411_3531.n1 a_3411_3531.t8 212.081
R12590 a_3411_3531.n4 a_3411_3531.n1 176.576
R12591 a_3411_3531.n2 a_3411_3531.t7 174.891
R12592 a_3411_3531.n0 a_3411_3531.t3 139.78
R12593 a_3411_3531.n1 a_3411_3531.t5 139.78
R12594 a_3411_3531.n5 a_3411_3531.t2 63.3219
R12595 a_3411_3531.t0 a_3411_3531.n5 63.3219
R12596 a_3411_3531.n1 a_3411_3531.n0 61.346
R12597 a_3411_3531.n4 a_3411_3531.n3 37.7195
R12598 auto_sampling_0.x3.D.n5 auto_sampling_0.x3.D.n4 585
R12599 auto_sampling_0.x3.D.n4 auto_sampling_0.x3.D.n3 585
R12600 auto_sampling_0.x3.D.n2 auto_sampling_0.x3.D.t5 333.651
R12601 auto_sampling_0.x3.D.n2 auto_sampling_0.x3.D.t4 297.233
R12602 auto_sampling_0.x3.D auto_sampling_0.x3.D.n2 196.493
R12603 auto_sampling_0.x3.D.n1 auto_sampling_0.x3.D.n0 185
R12604 auto_sampling_0.x3.D auto_sampling_0.x3.D.n1 49.0339
R12605 auto_sampling_0.x3.D.n3 auto_sampling_0.x3.D 44.2533
R12606 auto_sampling_0.x3.D.n4 auto_sampling_0.x3.D.t3 26.5955
R12607 auto_sampling_0.x3.D.n4 auto_sampling_0.x3.D.t2 26.5955
R12608 auto_sampling_0.x3.D.n0 auto_sampling_0.x3.D.t1 24.9236
R12609 auto_sampling_0.x3.D.n0 auto_sampling_0.x3.D.t0 24.9236
R12610 auto_sampling_0.x3.D.n5 auto_sampling_0.x3.D 15.6165
R12611 auto_sampling_0.x3.D.n1 auto_sampling_0.x3.D 10.4965
R12612 auto_sampling_0.x3.D.n3 auto_sampling_0.x3.D 1.7925
R12613 auto_sampling_0.x3.D auto_sampling_0.x3.D.n5 1.7925
R12614 a_5730_n5074.t1 a_5730_n5074.n3 370.026
R12615 a_5730_n5074.n0 a_5730_n5074.t2 351.356
R12616 a_5730_n5074.n1 a_5730_n5074.t4 334.717
R12617 a_5730_n5074.n3 a_5730_n5074.t0 325.971
R12618 a_5730_n5074.n1 a_5730_n5074.t5 309.935
R12619 a_5730_n5074.n0 a_5730_n5074.t3 305.683
R12620 a_5730_n5074.n2 a_5730_n5074.n0 16.879
R12621 a_5730_n5074.n3 a_5730_n5074.n2 10.8867
R12622 a_5730_n5074.n2 a_5730_n5074.n1 9.3005
R12623 a_6298_n5106.n3 a_6298_n5106.n2 647.119
R12624 a_6298_n5106.n1 a_6298_n5106.t5 350.253
R12625 a_6298_n5106.n2 a_6298_n5106.n0 260.339
R12626 a_6298_n5106.n2 a_6298_n5106.n1 246.119
R12627 a_6298_n5106.n1 a_6298_n5106.t4 189.588
R12628 a_6298_n5106.n3 a_6298_n5106.t0 89.1195
R12629 a_6298_n5106.n0 a_6298_n5106.t2 63.3338
R12630 a_6298_n5106.t3 a_6298_n5106.n3 41.0422
R12631 a_6298_n5106.n0 a_6298_n5106.t1 31.9797
R12632 a_816_n1457.t1 a_816_n1457.n3 370.026
R12633 a_816_n1457.n0 a_816_n1457.t4 351.356
R12634 a_816_n1457.n1 a_816_n1457.t5 334.717
R12635 a_816_n1457.n3 a_816_n1457.t0 325.971
R12636 a_816_n1457.n1 a_816_n1457.t3 309.935
R12637 a_816_n1457.n0 a_816_n1457.t2 305.683
R12638 a_816_n1457.n2 a_816_n1457.n0 16.879
R12639 a_816_n1457.n3 a_816_n1457.n2 10.8867
R12640 a_816_n1457.n2 a_816_n1457.n1 9.3005
R12641 a_n5259_n9484.t0 a_n5259_n9484.n3 370.026
R12642 a_n5259_n9484.n0 a_n5259_n9484.t4 351.356
R12643 a_n5259_n9484.n1 a_n5259_n9484.t3 334.717
R12644 a_n5259_n9484.n3 a_n5259_n9484.t1 325.971
R12645 a_n5259_n9484.n1 a_n5259_n9484.t5 309.935
R12646 a_n5259_n9484.n0 a_n5259_n9484.t2 305.683
R12647 a_n5259_n9484.n2 a_n5259_n9484.n0 16.879
R12648 a_n5259_n9484.n3 a_n5259_n9484.n2 10.8867
R12649 a_n5259_n9484.n2 a_n5259_n9484.n1 9.3005
R12650 a_n4344_n9484.n3 a_n4344_n9484.n2 636.953
R12651 a_n4344_n9484.n1 a_n4344_n9484.t5 366.856
R12652 a_n4344_n9484.n2 a_n4344_n9484.n0 300.2
R12653 a_n4344_n9484.n2 a_n4344_n9484.n1 225.036
R12654 a_n4344_n9484.n1 a_n4344_n9484.t4 174.056
R12655 a_n4344_n9484.n0 a_n4344_n9484.t0 70.0005
R12656 a_n4344_n9484.n3 a_n4344_n9484.t3 68.0124
R12657 a_n4344_n9484.t1 a_n4344_n9484.n3 63.3219
R12658 a_n4344_n9484.n0 a_n4344_n9484.t2 61.6672
R12659 a_n4182_n9118.t0 a_n4182_n9118.t1 126.644
R12660 a_4235_n9484.n1 a_4235_n9484.t5 530.01
R12661 a_4235_n9484.t1 a_4235_n9484.n5 421.021
R12662 a_4235_n9484.n0 a_4235_n9484.t3 337.142
R12663 a_4235_n9484.n3 a_4235_n9484.t0 280.223
R12664 a_4235_n9484.n4 a_4235_n9484.t6 263.173
R12665 a_4235_n9484.n4 a_4235_n9484.t2 227.826
R12666 a_4235_n9484.n0 a_4235_n9484.t4 199.762
R12667 a_4235_n9484.n2 a_4235_n9484.n1 170.81
R12668 a_4235_n9484.n2 a_4235_n9484.n0 167.321
R12669 a_4235_n9484.n5 a_4235_n9484.n4 152
R12670 a_4235_n9484.n1 a_4235_n9484.t7 141.923
R12671 a_4235_n9484.n3 a_4235_n9484.n2 10.8376
R12672 a_4235_n9484.n5 a_4235_n9484.n3 2.50485
R12673 a_4401_n9484.t1 a_4401_n9484.n3 370.026
R12674 a_4401_n9484.n0 a_4401_n9484.t4 351.356
R12675 a_4401_n9484.n1 a_4401_n9484.t3 334.717
R12676 a_4401_n9484.n3 a_4401_n9484.t0 325.971
R12677 a_4401_n9484.n1 a_4401_n9484.t2 309.935
R12678 a_4401_n9484.n0 a_4401_n9484.t5 305.683
R12679 a_4401_n9484.n2 a_4401_n9484.n0 16.879
R12680 a_4401_n9484.n3 a_4401_n9484.n2 10.8867
R12681 a_4401_n9484.n2 a_4401_n9484.n1 9.3005
R12682 a_6019_3557.n1 a_6019_3557.t5 530.01
R12683 a_6019_3557.t1 a_6019_3557.n5 421.021
R12684 a_6019_3557.n0 a_6019_3557.t2 337.142
R12685 a_6019_3557.n3 a_6019_3557.t0 280.223
R12686 a_6019_3557.n4 a_6019_3557.t6 263.173
R12687 a_6019_3557.n4 a_6019_3557.t7 227.826
R12688 a_6019_3557.n0 a_6019_3557.t3 199.762
R12689 a_6019_3557.n2 a_6019_3557.n1 170.81
R12690 a_6019_3557.n2 a_6019_3557.n0 167.321
R12691 a_6019_3557.n5 a_6019_3557.n4 152
R12692 a_6019_3557.n1 a_6019_3557.t4 141.923
R12693 a_6019_3557.n3 a_6019_3557.n2 10.8376
R12694 a_6019_3557.n5 a_6019_3557.n3 2.50485
R12695 a_6753_3799.n3 a_6753_3799.n2 647.119
R12696 a_6753_3799.n1 a_6753_3799.t5 350.253
R12697 a_6753_3799.n2 a_6753_3799.n0 260.339
R12698 a_6753_3799.n2 a_6753_3799.n1 246.119
R12699 a_6753_3799.n1 a_6753_3799.t4 189.588
R12700 a_6753_3799.n3 a_6753_3799.t2 89.1195
R12701 a_6753_3799.n0 a_6753_3799.t1 63.3338
R12702 a_6753_3799.t3 a_6753_3799.n3 41.0422
R12703 a_6753_3799.n0 a_6753_3799.t0 31.9797
R12704 a_847_3923.t0 a_847_3923.n0 1327.82
R12705 a_847_3923.n0 a_847_3923.t2 194.655
R12706 a_847_3923.n0 a_847_3923.t1 63.3219
R12707 a_6651_n1331.n1 a_6651_n1331.t6 530.01
R12708 a_6651_n1331.t1 a_6651_n1331.n5 421.021
R12709 a_6651_n1331.n0 a_6651_n1331.t2 337.171
R12710 a_6651_n1331.n3 a_6651_n1331.t0 280.223
R12711 a_6651_n1331.n4 a_6651_n1331.t4 263.173
R12712 a_6651_n1331.n4 a_6651_n1331.t3 227.826
R12713 a_6651_n1331.n0 a_6651_n1331.t7 199.762
R12714 a_6651_n1331.n2 a_6651_n1331.n1 170.81
R12715 a_6651_n1331.n2 a_6651_n1331.n0 167.321
R12716 a_6651_n1331.n5 a_6651_n1331.n4 152
R12717 a_6651_n1331.n1 a_6651_n1331.t5 141.923
R12718 a_6651_n1331.n3 a_6651_n1331.n2 10.8376
R12719 a_6651_n1331.n5 a_6651_n1331.n3 2.50485
R12720 a_6738_n1573.n3 a_6738_n1573.n2 647.119
R12721 a_6738_n1573.n1 a_6738_n1573.t4 350.253
R12722 a_6738_n1573.n2 a_6738_n1573.n0 260.339
R12723 a_6738_n1573.n2 a_6738_n1573.n1 246.119
R12724 a_6738_n1573.n1 a_6738_n1573.t5 189.588
R12725 a_6738_n1573.n3 a_6738_n1573.t0 89.1195
R12726 a_6738_n1573.n0 a_6738_n1573.t2 63.3338
R12727 a_6738_n1573.t3 a_6738_n1573.n3 41.0422
R12728 a_6738_n1573.n0 a_6738_n1573.t1 31.9797
R12729 a_4680_n1457.t1 a_4680_n1457.n3 370.026
R12730 a_4680_n1457.n0 a_4680_n1457.t2 351.356
R12731 a_4680_n1457.n1 a_4680_n1457.t5 334.717
R12732 a_4680_n1457.n3 a_4680_n1457.t0 325.971
R12733 a_4680_n1457.n1 a_4680_n1457.t3 309.935
R12734 a_4680_n1457.n0 a_4680_n1457.t4 305.683
R12735 a_4680_n1457.n2 a_4680_n1457.n0 16.879
R12736 a_4680_n1457.n3 a_4680_n1457.n2 10.8867
R12737 a_4680_n1457.n2 a_4680_n1457.n1 9.3005
R12738 a_4402_n1441.n3 a_4402_n1441.n2 636.953
R12739 a_4402_n1441.n1 a_4402_n1441.t4 366.856
R12740 a_4402_n1441.n2 a_4402_n1441.n0 300.2
R12741 a_4402_n1441.n2 a_4402_n1441.n1 225.036
R12742 a_4402_n1441.n1 a_4402_n1441.t5 174.056
R12743 a_4402_n1441.n0 a_4402_n1441.t1 70.0005
R12744 a_4402_n1441.t0 a_4402_n1441.n3 68.0124
R12745 a_4402_n1441.n3 a_4402_n1441.t2 63.3219
R12746 a_4402_n1441.n0 a_4402_n1441.t3 61.6672
R12747 a_4806_n1573.n3 a_4806_n1573.n2 647.119
R12748 a_4806_n1573.n1 a_4806_n1573.t5 350.253
R12749 a_4806_n1573.n2 a_4806_n1573.n0 260.339
R12750 a_4806_n1573.n2 a_4806_n1573.n1 246.119
R12751 a_4806_n1573.n1 a_4806_n1573.t4 189.588
R12752 a_4806_n1573.n3 a_4806_n1573.t0 89.1195
R12753 a_4806_n1573.n0 a_4806_n1573.t3 63.3338
R12754 a_4806_n1573.t1 a_4806_n1573.n3 41.0422
R12755 a_4806_n1573.n0 a_4806_n1573.t2 31.9797
R12756 a_4401_n10022.t1 a_4401_n10022.n3 370.026
R12757 a_4401_n10022.n0 a_4401_n10022.t2 351.356
R12758 a_4401_n10022.n1 a_4401_n10022.t5 334.717
R12759 a_4401_n10022.n3 a_4401_n10022.t0 325.971
R12760 a_4401_n10022.n1 a_4401_n10022.t3 309.935
R12761 a_4401_n10022.n0 a_4401_n10022.t4 305.683
R12762 a_4401_n10022.n2 a_4401_n10022.n0 16.879
R12763 a_4401_n10022.n3 a_4401_n10022.n2 10.8867
R12764 a_4401_n10022.n2 a_4401_n10022.n1 9.3005
R12765 a_n480_n9484.n3 a_n480_n9484.n2 636.953
R12766 a_n480_n9484.n1 a_n480_n9484.t5 366.856
R12767 a_n480_n9484.n2 a_n480_n9484.n0 300.2
R12768 a_n480_n9484.n2 a_n480_n9484.n1 225.036
R12769 a_n480_n9484.n1 a_n480_n9484.t4 174.056
R12770 a_n480_n9484.n0 a_n480_n9484.t2 70.0005
R12771 a_n480_n9484.n3 a_n480_n9484.t3 68.0124
R12772 a_n480_n9484.t0 a_n480_n9484.n3 63.3219
R12773 a_n480_n9484.n0 a_n480_n9484.t1 61.6672
R12774 a_n4647_n9662.t0 a_n4647_n9662.t1 60.0005
R12775 a_284_n4702.n3 a_284_n4702.n2 674.338
R12776 a_284_n4702.n1 a_284_n4702.t4 332.58
R12777 a_284_n4702.n2 a_284_n4702.n0 284.012
R12778 a_284_n4702.n2 a_284_n4702.n1 253.648
R12779 a_284_n4702.n1 a_284_n4702.t5 168.701
R12780 a_284_n4702.n3 a_284_n4702.t2 96.1553
R12781 a_284_n4702.t1 a_284_n4702.n3 65.6672
R12782 a_284_n4702.n0 a_284_n4702.t3 65.0005
R12783 a_284_n4702.n0 a_284_n4702.t0 45.0005
R12784 a_380_n4702.t1 a_380_n4702.t0 198.571
R12785 a_8739_n1599.n3 a_8739_n1599.n2 674.338
R12786 a_8739_n1599.n1 a_8739_n1599.t5 332.58
R12787 a_8739_n1599.n2 a_8739_n1599.n0 284.012
R12788 a_8739_n1599.n2 a_8739_n1599.n1 253.648
R12789 a_8739_n1599.n1 a_8739_n1599.t4 168.701
R12790 a_8739_n1599.t0 a_8739_n1599.n3 96.1553
R12791 a_8739_n1599.n3 a_8739_n1599.t3 65.6672
R12792 a_8739_n1599.n0 a_8739_n1599.t1 65.0005
R12793 a_8739_n1599.n0 a_8739_n1599.t2 45.0005
R12794 a_9302_n1573.n1 a_9302_n1573.n0 926.024
R12795 a_9302_n1573.t1 a_9302_n1573.n1 82.0838
R12796 a_9302_n1573.n0 a_9302_n1573.t0 63.3338
R12797 a_9302_n1573.n1 a_9302_n1573.t3 63.3219
R12798 a_9302_n1573.n0 a_9302_n1573.t2 29.7268
R12799 a_1627_n9724.n4 a_1627_n9724.n1 807.871
R12800 a_1627_n9724.n0 a_1627_n9724.t7 389.183
R12801 a_1627_n9724.n5 a_1627_n9724.n0 251.167
R12802 a_1627_n9724.t0 a_1627_n9724.n5 223.571
R12803 a_1627_n9724.n2 a_1627_n9724.t8 212.081
R12804 a_1627_n9724.n3 a_1627_n9724.t6 212.081
R12805 a_1627_n9724.n4 a_1627_n9724.n3 176.576
R12806 a_1627_n9724.n0 a_1627_n9724.t5 174.891
R12807 a_1627_n9724.n2 a_1627_n9724.t4 139.78
R12808 a_1627_n9724.n3 a_1627_n9724.t3 139.78
R12809 a_1627_n9724.n1 a_1627_n9724.t1 63.3219
R12810 a_1627_n9724.n1 a_1627_n9724.t2 63.3219
R12811 a_1627_n9724.n3 a_1627_n9724.n2 61.346
R12812 a_1627_n9724.n5 a_1627_n9724.n4 37.7195
R12813 SWN[5].n4 SWN[5].n3 585
R12814 SWN[5].n3 SWN[5].n2 585
R12815 SWN[5].n1 SWN[5].n0 185
R12816 SWN[5].n5 SWN[5].n1 53.3859
R12817 SWN[5].n3 SWN[5].t2 26.5955
R12818 SWN[5].n3 SWN[5].t3 26.5955
R12819 SWN[5].n0 SWN[5].t0 24.9236
R12820 SWN[5].n0 SWN[5].t1 24.9236
R12821 SWN[5] SWN[5].n5 14.676
R12822 SWN[5] SWN[5].n4 10.4965
R12823 SWN[5].n2 SWN[5] 10.4965
R12824 SWN[5].n4 SWN[5] 6.9125
R12825 SWN[5].n2 SWN[5] 6.9125
R12826 SWN[5].n5 SWN[5] 4.3525
R12827 SWN[5].n1 SWN[5] 1.7925
R12828 auto_sampling_0.x7.Q.n5 auto_sampling_0.x7.Q.n4 585
R12829 auto_sampling_0.x7.Q.n4 auto_sampling_0.x7.Q.n3 585
R12830 auto_sampling_0.x7.Q.n2 auto_sampling_0.x7.Q.t4 333.651
R12831 auto_sampling_0.x7.Q.n2 auto_sampling_0.x7.Q.t5 297.233
R12832 auto_sampling_0.x7.Q auto_sampling_0.x7.Q.n2 196.493
R12833 auto_sampling_0.x7.Q.n1 auto_sampling_0.x7.Q.n0 185
R12834 auto_sampling_0.x7.Q auto_sampling_0.x7.Q.n1 49.0339
R12835 auto_sampling_0.x7.Q.n3 auto_sampling_0.x7.Q 44.2533
R12836 auto_sampling_0.x7.Q.n4 auto_sampling_0.x7.Q.t2 26.5955
R12837 auto_sampling_0.x7.Q.n4 auto_sampling_0.x7.Q.t3 26.5955
R12838 auto_sampling_0.x7.Q.n0 auto_sampling_0.x7.Q.t0 24.9236
R12839 auto_sampling_0.x7.Q.n0 auto_sampling_0.x7.Q.t1 24.9236
R12840 auto_sampling_0.x7.Q.n5 auto_sampling_0.x7.Q 15.6165
R12841 auto_sampling_0.x7.Q.n1 auto_sampling_0.x7.Q 10.4965
R12842 auto_sampling_0.x7.Q.n3 auto_sampling_0.x7.Q 1.7925
R12843 auto_sampling_0.x7.Q auto_sampling_0.x7.Q.n5 1.7925
R12844 a_644_3557.n1 a_644_3557.n0 926.024
R12845 a_644_3557.t0 a_644_3557.n1 82.0838
R12846 a_644_3557.n0 a_644_3557.t1 63.3338
R12847 a_644_3557.n1 a_644_3557.t3 63.3219
R12848 a_644_3557.n0 a_644_3557.t2 29.7268
R12849 a_371_n10022.n1 a_371_n10022.t4 530.01
R12850 a_371_n10022.t1 a_371_n10022.n5 421.021
R12851 a_371_n10022.n0 a_371_n10022.t5 337.142
R12852 a_371_n10022.n3 a_371_n10022.t0 280.223
R12853 a_371_n10022.n4 a_371_n10022.t6 263.173
R12854 a_371_n10022.n4 a_371_n10022.t3 227.826
R12855 a_371_n10022.n0 a_371_n10022.t7 199.762
R12856 a_371_n10022.n2 a_371_n10022.n1 170.81
R12857 a_371_n10022.n2 a_371_n10022.n0 167.321
R12858 a_371_n10022.n5 a_371_n10022.n4 152
R12859 a_371_n10022.n1 a_371_n10022.t2 141.923
R12860 a_371_n10022.n3 a_371_n10022.n2 10.8376
R12861 a_371_n10022.n5 a_371_n10022.n3 2.50485
R12862 CKO.n2 CKO 586.253
R12863 CKO.n3 CKO.n2 585
R12864 CKO.n4 CKO.t3 339.418
R12865 CKO.n36 CKO.t17 294.557
R12866 CKO.n33 CKO.t16 294.557
R12867 CKO.n30 CKO.t8 294.557
R12868 CKO.n26 CKO.t9 294.557
R12869 CKO.n24 CKO.t23 294.557
R12870 CKO.n20 CKO.t6 294.557
R12871 CKO.n18 CKO.t14 294.557
R12872 CKO.n15 CKO.t7 294.557
R12873 CKO.n12 CKO.t20 294.557
R12874 CKO.n9 CKO.t12 294.557
R12875 CKO.n5 CKO.t2 274.06
R12876 CKO.n0 CKO.t1 274.06
R12877 CKO.n36 CKO.t13 211.01
R12878 CKO.n33 CKO.t10 211.01
R12879 CKO.n30 CKO.t4 211.01
R12880 CKO.n26 CKO.t5 211.01
R12881 CKO.n24 CKO.t21 211.01
R12882 CKO.n20 CKO.t11 211.01
R12883 CKO.n18 CKO.t19 211.01
R12884 CKO.n15 CKO.t15 211.01
R12885 CKO.n12 CKO.t22 211.01
R12886 CKO.n9 CKO.t18 211.01
R12887 CKO CKO.n36 156.207
R12888 CKO CKO.n33 156.207
R12889 CKO CKO.n30 156.207
R12890 CKO CKO.n26 156.207
R12891 CKO CKO.n24 156.207
R12892 CKO.n21 CKO.n20 152
R12893 CKO.n19 CKO.n18 152
R12894 CKO.n16 CKO.n15 152
R12895 CKO.n13 CKO.n12 152
R12896 CKO.n10 CKO.n9 152
R12897 CKO.n2 CKO.t0 46.2955
R12898 CKO.n22 CKO 18.9565
R12899 CKO.n28 CKO.n25 18.5908
R12900 CKO.n1 CKO 15.3605
R12901 CKO.n8 CKO 14.5568
R12902 CKO.n22 CKO 14.1662
R12903 CKO.n17 CKO 14.1662
R12904 CKO.n38 CKO.n37 13.8005
R12905 CKO.n35 CKO.n34 13.8005
R12906 CKO.n32 CKO.n31 13.8005
R12907 CKO.n28 CKO.n27 13.8005
R12908 CKO.n14 CKO 13.8005
R12909 CKO.n11 CKO 13.8005
R12910 CKO.n8 CKO.n7 13.8005
R12911 CKO CKO.n5 11.2645
R12912 CKO CKO.n21 10.4234
R12913 CKO CKO.n19 10.4234
R12914 CKO CKO.n16 10.4234
R12915 CKO CKO.n13 10.4234
R12916 CKO CKO.n10 10.4234
R12917 CKO.n3 CKO 8.2092
R12918 CKO.n6 CKO 6.6565
R12919 CKO.n31 CKO 6.58336
R12920 CKO.n27 CKO 6.58336
R12921 CKO.n25 CKO 6.58336
R12922 CKO.n37 CKO 6.21764
R12923 CKO.n37 CKO 6.21764
R12924 CKO.n34 CKO 6.21764
R12925 CKO.n34 CKO 6.21764
R12926 CKO.n5 CKO 6.1445
R12927 CKO.n31 CKO 5.85193
R12928 CKO.n27 CKO 5.85193
R12929 CKO.n25 CKO 5.85193
R12930 CKO.n14 CKO.n11 4.79078
R12931 CKO.n17 CKO.n14 4.79078
R12932 CKO.n35 CKO.n32 4.79078
R12933 CKO.n38 CKO.n35 4.79078
R12934 CKO.n6 CKO 3.61789
R12935 CKO.n7 CKO.n4 2.97835
R12936 CKO.n29 CKO.n28 2.88814
R12937 CKO.n5 CKO 2.86947
R12938 CKO.n0 CKO 2.86947
R12939 CKO.n23 CKO.n17 2.65814
R12940 CKO CKO.n0 2.5605
R12941 CKO.n23 CKO.n22 2.13314
R12942 CKO.n1 CKO 2.0485
R12943 CKO.n21 CKO 2.01193
R12944 CKO.n19 CKO 2.01193
R12945 CKO.n16 CKO 2.01193
R12946 CKO.n13 CKO 2.01193
R12947 CKO.n10 CKO 2.01193
R12948 CKO.n32 CKO.n29 1.90314
R12949 CKO.n4 CKO 1.74382
R12950 CKO CKO.n3 1.25267
R12951 CKO.n29 CKO.n23 1.1455
R12952 CKO.n7 CKO.n6 1.11354
R12953 CKO CKO.n1 1.11354
R12954 CKO CKO.n38 0.940597
R12955 CKO.n11 CKO.n8 0.383812
R12956 a_3632_n5074.n1 a_3632_n5074.t5 530.01
R12957 a_3632_n5074.t1 a_3632_n5074.n5 421.021
R12958 a_3632_n5074.n0 a_3632_n5074.t3 337.142
R12959 a_3632_n5074.n3 a_3632_n5074.t0 280.223
R12960 a_3632_n5074.n4 a_3632_n5074.t4 263.173
R12961 a_3632_n5074.n4 a_3632_n5074.t2 227.826
R12962 a_3632_n5074.n0 a_3632_n5074.t7 199.762
R12963 a_3632_n5074.n2 a_3632_n5074.n1 170.81
R12964 a_3632_n5074.n2 a_3632_n5074.n0 167.321
R12965 a_3632_n5074.n5 a_3632_n5074.n4 152
R12966 a_3632_n5074.n1 a_3632_n5074.t6 141.923
R12967 a_3632_n5074.n3 a_3632_n5074.n2 10.8376
R12968 a_3632_n5074.n5 a_3632_n5074.n3 2.50485
R12969 a_5491_n9510.n5 a_5491_n9510.n4 807.871
R12970 a_5491_n9510.n2 a_5491_n9510.t6 389.183
R12971 a_5491_n9510.n3 a_5491_n9510.n2 251.167
R12972 a_5491_n9510.n3 a_5491_n9510.t1 223.571
R12973 a_5491_n9510.n0 a_5491_n9510.t8 212.081
R12974 a_5491_n9510.n1 a_5491_n9510.t4 212.081
R12975 a_5491_n9510.n4 a_5491_n9510.n1 176.576
R12976 a_5491_n9510.n2 a_5491_n9510.t5 174.891
R12977 a_5491_n9510.n0 a_5491_n9510.t7 139.78
R12978 a_5491_n9510.n1 a_5491_n9510.t3 139.78
R12979 a_5491_n9510.t0 a_5491_n9510.n5 63.3219
R12980 a_5491_n9510.n5 a_5491_n9510.t2 63.3219
R12981 a_5491_n9510.n1 a_5491_n9510.n0 61.346
R12982 a_5491_n9510.n4 a_5491_n9510.n3 37.7195
R12983 SWP[7].n0 SWP[7].t4 333.651
R12984 SWP[7].n0 SWP[7].t5 297.233
R12985 SWP[7].n4 SWP[7].n3 289.096
R12986 SWP[7].n1 SWP[7].n0 196.493
R12987 SWP[7].n6 SWP[7].n5 185
R12988 SWP[7] SWP[7].n6 49.0339
R12989 SWP[7] SWP[7].n1 39.5081
R12990 SWP[7].n2 SWP[7] 37.6912
R12991 SWP[7].n3 SWP[7].t2 26.5955
R12992 SWP[7].n3 SWP[7].t3 26.5955
R12993 SWP[7].n5 SWP[7].t0 24.9236
R12994 SWP[7].n5 SWP[7].t1 24.9236
R12995 SWP[7] SWP[7].n7 14.6135
R12996 SWP[7].n2 SWP[7] 13.5849
R12997 SWP[7].n7 SWP[7] 13.0565
R12998 SWP[7].n6 SWP[7] 10.4965
R12999 SWP[7] SWP[7].n4 9.48653
R13000 SWP[7].n4 SWP[7] 7.7181
R13001 SWP[7] SWP[7].n2 5.10179
R13002 SWP[7].n7 SWP[7] 4.3525
R13003 SWP[7].n1 SWP[7] 0.24431
R13004 a_1304_3557.n3 a_1304_3557.n2 636.953
R13005 a_1304_3557.n1 a_1304_3557.t5 366.856
R13006 a_1304_3557.n2 a_1304_3557.n0 300.2
R13007 a_1304_3557.n2 a_1304_3557.n1 225.036
R13008 a_1304_3557.n1 a_1304_3557.t4 174.056
R13009 a_1304_3557.n0 a_1304_3557.t1 70.0005
R13010 a_1304_3557.n3 a_1304_3557.t2 68.0124
R13011 a_1304_3557.t0 a_1304_3557.n3 63.3219
R13012 a_1304_3557.n0 a_1304_3557.t3 61.6672
R13013 a_4087_3557.n1 a_4087_3557.t3 530.01
R13014 a_4087_3557.t1 a_4087_3557.n5 421.021
R13015 a_4087_3557.n0 a_4087_3557.t6 337.142
R13016 a_4087_3557.n3 a_4087_3557.t0 280.223
R13017 a_4087_3557.n4 a_4087_3557.t4 263.173
R13018 a_4087_3557.n4 a_4087_3557.t5 227.826
R13019 a_4087_3557.n0 a_4087_3557.t7 199.762
R13020 a_4087_3557.n2 a_4087_3557.n1 170.81
R13021 a_4087_3557.n2 a_4087_3557.n0 167.321
R13022 a_4087_3557.n5 a_4087_3557.n4 152
R13023 a_4087_3557.n1 a_4087_3557.t2 141.923
R13024 a_4087_3557.n3 a_4087_3557.n2 10.8376
R13025 a_4087_3557.n5 a_4087_3557.n3 2.50485
R13026 a_4508_3557.n1 a_4508_3557.n0 926.024
R13027 a_4508_3557.n0 a_4508_3557.t3 82.0838
R13028 a_4508_3557.n1 a_4508_3557.t0 63.3338
R13029 a_4508_3557.n0 a_4508_3557.t2 63.3219
R13030 a_4508_3557.n2 a_4508_3557.t1 26.3935
R13031 a_4508_3557.n3 a_4508_3557.n2 14.4005
R13032 a_4508_3557.n2 a_4508_3557.n1 3.33383
R13033 a_4603_3557.n3 a_4603_3557.n2 674.338
R13034 a_4603_3557.n1 a_4603_3557.t4 332.58
R13035 a_4603_3557.n2 a_4603_3557.n0 284.012
R13036 a_4603_3557.n2 a_4603_3557.n1 253.648
R13037 a_4603_3557.n1 a_4603_3557.t5 168.701
R13038 a_4603_3557.t0 a_4603_3557.n3 96.1553
R13039 a_4603_3557.n3 a_4603_3557.t2 65.6672
R13040 a_4603_3557.n0 a_4603_3557.t1 65.0005
R13041 a_4603_3557.n0 a_4603_3557.t3 45.0005
R13042 a_n9123_n10022.t0 a_n9123_n10022.n3 370.026
R13043 a_n9123_n10022.n0 a_n9123_n10022.t2 351.356
R13044 a_n9123_n10022.n1 a_n9123_n10022.t5 334.717
R13045 a_n9123_n10022.n3 a_n9123_n10022.t1 325.971
R13046 a_n9123_n10022.n1 a_n9123_n10022.t4 309.935
R13047 a_n9123_n10022.n0 a_n9123_n10022.t3 305.683
R13048 a_n9123_n10022.n2 a_n9123_n10022.n0 16.879
R13049 a_n9123_n10022.n3 a_n9123_n10022.n2 10.8867
R13050 a_n9123_n10022.n2 a_n9123_n10022.n1 9.3005
R13051 a_n8555_n10054.n3 a_n8555_n10054.n2 647.119
R13052 a_n8555_n10054.n1 a_n8555_n10054.t4 350.253
R13053 a_n8555_n10054.n2 a_n8555_n10054.n0 260.339
R13054 a_n8555_n10054.n2 a_n8555_n10054.n1 246.119
R13055 a_n8555_n10054.n1 a_n8555_n10054.t5 189.588
R13056 a_n8555_n10054.n3 a_n8555_n10054.t3 89.1195
R13057 a_n8555_n10054.n0 a_n8555_n10054.t1 63.3338
R13058 a_n8555_n10054.t2 a_n8555_n10054.n3 41.0422
R13059 a_n8555_n10054.n0 a_n8555_n10054.t0 31.9797
R13060 a_n8208_n9650.n3 a_n8208_n9650.n2 636.953
R13061 a_n8208_n9650.n1 a_n8208_n9650.t4 366.856
R13062 a_n8208_n9650.n2 a_n8208_n9650.n0 300.2
R13063 a_n8208_n9650.n2 a_n8208_n9650.n1 225.036
R13064 a_n8208_n9650.n1 a_n8208_n9650.t5 174.056
R13065 a_n8208_n9650.n0 a_n8208_n9650.t0 70.0005
R13066 a_n8208_n9650.n3 a_n8208_n9650.t2 68.0124
R13067 a_n8208_n9650.t1 a_n8208_n9650.n3 63.3219
R13068 a_n8208_n9650.n0 a_n8208_n9650.t3 61.6672
R13069 a_2787_n1331.n1 a_2787_n1331.t2 530.01
R13070 a_2787_n1331.t1 a_2787_n1331.n5 421.021
R13071 a_2787_n1331.n0 a_2787_n1331.t3 337.171
R13072 a_2787_n1331.n3 a_2787_n1331.t0 280.223
R13073 a_2787_n1331.n4 a_2787_n1331.t7 263.173
R13074 a_2787_n1331.n4 a_2787_n1331.t5 227.826
R13075 a_2787_n1331.n0 a_2787_n1331.t4 199.762
R13076 a_2787_n1331.n2 a_2787_n1331.n1 170.81
R13077 a_2787_n1331.n2 a_2787_n1331.n0 167.321
R13078 a_2787_n1331.n5 a_2787_n1331.n4 152
R13079 a_2787_n1331.n1 a_2787_n1331.t6 141.923
R13080 a_2787_n1331.n3 a_2787_n1331.n2 10.8376
R13081 a_2787_n1331.n5 a_2787_n1331.n3 2.50485
R13082 a_5330_3923.t0 a_5330_3923.t1 126.644
R13083 a_n7191_n10022.t1 a_n7191_n10022.n3 370.026
R13084 a_n7191_n10022.n0 a_n7191_n10022.t2 351.356
R13085 a_n7191_n10022.n1 a_n7191_n10022.t3 334.717
R13086 a_n7191_n10022.n3 a_n7191_n10022.t0 325.971
R13087 a_n7191_n10022.n1 a_n7191_n10022.t5 309.935
R13088 a_n7191_n10022.n0 a_n7191_n10022.t4 305.683
R13089 a_n7191_n10022.n2 a_n7191_n10022.n0 16.879
R13090 a_n7191_n10022.n3 a_n7191_n10022.n2 10.8867
R13091 a_n7191_n10022.n2 a_n7191_n10022.n1 9.3005
R13092 a_n4169_n9724.n4 a_n4169_n9724.n1 807.871
R13093 a_n4169_n9724.n0 a_n4169_n9724.t6 389.183
R13094 a_n4169_n9724.n5 a_n4169_n9724.n0 251.167
R13095 a_n4169_n9724.t0 a_n4169_n9724.n5 223.571
R13096 a_n4169_n9724.n2 a_n4169_n9724.t4 212.081
R13097 a_n4169_n9724.n3 a_n4169_n9724.t7 212.081
R13098 a_n4169_n9724.n4 a_n4169_n9724.n3 176.576
R13099 a_n4169_n9724.n0 a_n4169_n9724.t8 174.891
R13100 a_n4169_n9724.n2 a_n4169_n9724.t5 139.78
R13101 a_n4169_n9724.n3 a_n4169_n9724.t3 139.78
R13102 a_n4169_n9724.n1 a_n4169_n9724.t1 63.3219
R13103 a_n4169_n9724.n1 a_n4169_n9724.t2 63.3219
R13104 a_n4169_n9724.n3 a_n4169_n9724.n2 61.346
R13105 a_n4169_n9724.n5 a_n4169_n9724.n4 37.7195
R13106 a_4055_n1029.n1 a_4055_n1029.t7 530.01
R13107 a_4055_n1029.t1 a_4055_n1029.n5 421.021
R13108 a_4055_n1029.n0 a_4055_n1029.t3 337.142
R13109 a_4055_n1029.n3 a_4055_n1029.t0 280.223
R13110 a_4055_n1029.n4 a_4055_n1029.t6 263.173
R13111 a_4055_n1029.n4 a_4055_n1029.t5 227.826
R13112 a_4055_n1029.n0 a_4055_n1029.t2 199.762
R13113 a_4055_n1029.n2 a_4055_n1029.n1 170.81
R13114 a_4055_n1029.n2 a_4055_n1029.n0 167.321
R13115 a_4055_n1029.n5 a_4055_n1029.n4 152
R13116 a_4055_n1029.n1 a_4055_n1029.t4 141.923
R13117 a_4055_n1029.n3 a_4055_n1029.n2 10.8376
R13118 a_4055_n1029.n5 a_4055_n1029.n3 2.50485
R13119 a_n8033_n9510.n5 a_n8033_n9510.n4 807.871
R13120 a_n8033_n9510.n2 a_n8033_n9510.t4 389.183
R13121 a_n8033_n9510.n3 a_n8033_n9510.n2 251.167
R13122 a_n8033_n9510.n3 a_n8033_n9510.t1 223.571
R13123 a_n8033_n9510.n0 a_n8033_n9510.t8 212.081
R13124 a_n8033_n9510.n1 a_n8033_n9510.t6 212.081
R13125 a_n8033_n9510.n4 a_n8033_n9510.n1 176.576
R13126 a_n8033_n9510.n2 a_n8033_n9510.t3 174.891
R13127 a_n8033_n9510.n0 a_n8033_n9510.t7 139.78
R13128 a_n8033_n9510.n1 a_n8033_n9510.t5 139.78
R13129 a_n8033_n9510.t0 a_n8033_n9510.n5 63.3219
R13130 a_n8033_n9510.n5 a_n8033_n9510.t2 63.3219
R13131 a_n8033_n9510.n1 a_n8033_n9510.n0 61.346
R13132 a_n8033_n9510.n4 a_n8033_n9510.n3 37.7195
R13133 a_n8099_n9484.t1 a_n8099_n9484.t0 94.7268
R13134 a_n10393_n9484.n22 a_n10393_n9484.t2 286.348
R13135 a_n10393_n9484.n24 a_n10393_n9484.t3 271.051
R13136 a_n10393_n9484.n4 a_n10393_n9484.t18 221.72
R13137 a_n10393_n9484.n5 a_n10393_n9484.t15 221.72
R13138 a_n10393_n9484.n3 a_n10393_n9484.t21 221.72
R13139 a_n10393_n9484.n9 a_n10393_n9484.t19 221.72
R13140 a_n10393_n9484.n11 a_n10393_n9484.t9 221.72
R13141 a_n10393_n9484.n1 a_n10393_n9484.t7 221.72
R13142 a_n10393_n9484.n17 a_n10393_n9484.t13 221.72
R13143 a_n10393_n9484.n18 a_n10393_n9484.t11 221.72
R13144 a_n10393_n9484.n25 a_n10393_n9484.n24 206.055
R13145 a_n10393_n9484.n22 a_n10393_n9484.n21 198.177
R13146 a_n10393_n9484.n7 a_n10393_n9484.n6 177.601
R13147 a_n10393_n9484.n20 a_n10393_n9484.n19 152
R13148 a_n10393_n9484.n16 a_n10393_n9484.n0 152
R13149 a_n10393_n9484.n15 a_n10393_n9484.n14 152
R13150 a_n10393_n9484.n13 a_n10393_n9484.n12 152
R13151 a_n10393_n9484.n10 a_n10393_n9484.n2 152
R13152 a_n10393_n9484.n8 a_n10393_n9484.n7 152
R13153 a_n10393_n9484.n4 a_n10393_n9484.t16 149.421
R13154 a_n10393_n9484.n5 a_n10393_n9484.t14 149.421
R13155 a_n10393_n9484.n3 a_n10393_n9484.t20 149.421
R13156 a_n10393_n9484.n9 a_n10393_n9484.t17 149.421
R13157 a_n10393_n9484.n11 a_n10393_n9484.t8 149.421
R13158 a_n10393_n9484.n1 a_n10393_n9484.t6 149.421
R13159 a_n10393_n9484.n17 a_n10393_n9484.t12 149.421
R13160 a_n10393_n9484.n18 a_n10393_n9484.t10 149.421
R13161 a_n10393_n9484.n5 a_n10393_n9484.n4 74.9783
R13162 a_n10393_n9484.n6 a_n10393_n9484.n5 66.0523
R13163 a_n10393_n9484.n16 a_n10393_n9484.n15 60.6968
R13164 a_n10393_n9484.n19 a_n10393_n9484.n17 55.3412
R13165 a_n10393_n9484.n8 a_n10393_n9484.n3 51.7709
R13166 a_n10393_n9484.n12 a_n10393_n9484.n1 51.7709
R13167 a_n10393_n9484.n23 a_n10393_n9484.n22 48.9632
R13168 a_n10393_n9484.n24 a_n10393_n9484.n23 38.7339
R13169 a_n10393_n9484.n10 a_n10393_n9484.n9 37.4894
R13170 a_n10393_n9484.n11 a_n10393_n9484.n10 37.4894
R13171 a_n10393_n9484.t1 a_n10393_n9484.n25 26.5955
R13172 a_n10393_n9484.n25 a_n10393_n9484.t5 26.5955
R13173 a_n10393_n9484.n7 a_n10393_n9484.n2 25.6005
R13174 a_n10393_n9484.n13 a_n10393_n9484.n2 25.6005
R13175 a_n10393_n9484.n14 a_n10393_n9484.n13 25.6005
R13176 a_n10393_n9484.n14 a_n10393_n9484.n0 25.6005
R13177 a_n10393_n9484.n20 a_n10393_n9484.n0 25.6005
R13178 a_n10393_n9484.n21 a_n10393_n9484.t0 24.9236
R13179 a_n10393_n9484.n21 a_n10393_n9484.t4 24.9236
R13180 a_n10393_n9484.n9 a_n10393_n9484.n8 23.2079
R13181 a_n10393_n9484.n12 a_n10393_n9484.n11 23.2079
R13182 a_n10393_n9484.n19 a_n10393_n9484.n18 19.6375
R13183 a_n10393_n9484.n23 a_n10393_n9484.n20 18.4476
R13184 a_n10393_n9484.n6 a_n10393_n9484.n3 8.92643
R13185 a_n10393_n9484.n15 a_n10393_n9484.n1 8.92643
R13186 a_n10393_n9484.n17 a_n10393_n9484.n16 5.35606
R13187 cdac_ctrl_0.x1.X.n39 cdac_ctrl_0.x1.X.n37 374.966
R13188 cdac_ctrl_0.x1.X.n31 cdac_ctrl_0.x1.X.t22 333.651
R13189 cdac_ctrl_0.x1.X.n28 cdac_ctrl_0.x1.X.t29 333.651
R13190 cdac_ctrl_0.x1.X.n25 cdac_ctrl_0.x1.X.t33 333.651
R13191 cdac_ctrl_0.x1.X.n22 cdac_ctrl_0.x1.X.t16 333.651
R13192 cdac_ctrl_0.x1.X.n19 cdac_ctrl_0.x1.X.t21 333.651
R13193 cdac_ctrl_0.x1.X.n16 cdac_ctrl_0.x1.X.t31 333.651
R13194 cdac_ctrl_0.x1.X.n13 cdac_ctrl_0.x1.X.t24 333.651
R13195 cdac_ctrl_0.x1.X.n10 cdac_ctrl_0.x1.X.t27 333.651
R13196 cdac_ctrl_0.x1.X.n7 cdac_ctrl_0.x1.X.t18 333.651
R13197 cdac_ctrl_0.x1.X.n5 cdac_ctrl_0.x1.X.t30 333.651
R13198 cdac_ctrl_0.x1.X.n40 cdac_ctrl_0.x1.X.n36 311.717
R13199 cdac_ctrl_0.x1.X.n39 cdac_ctrl_0.x1.X.n38 311.717
R13200 cdac_ctrl_0.x1.X.n31 cdac_ctrl_0.x1.X.t28 297.233
R13201 cdac_ctrl_0.x1.X.n28 cdac_ctrl_0.x1.X.t32 297.233
R13202 cdac_ctrl_0.x1.X.n25 cdac_ctrl_0.x1.X.t35 297.233
R13203 cdac_ctrl_0.x1.X.n22 cdac_ctrl_0.x1.X.t17 297.233
R13204 cdac_ctrl_0.x1.X.n19 cdac_ctrl_0.x1.X.t25 297.233
R13205 cdac_ctrl_0.x1.X.n16 cdac_ctrl_0.x1.X.t20 297.233
R13206 cdac_ctrl_0.x1.X.n13 cdac_ctrl_0.x1.X.t19 297.233
R13207 cdac_ctrl_0.x1.X.n10 cdac_ctrl_0.x1.X.t34 297.233
R13208 cdac_ctrl_0.x1.X.n7 cdac_ctrl_0.x1.X.t23 297.233
R13209 cdac_ctrl_0.x1.X.n5 cdac_ctrl_0.x1.X.t26 297.233
R13210 cdac_ctrl_0.x1.X.n35 cdac_ctrl_0.x1.X.n34 284.19
R13211 cdac_ctrl_0.x1.X.n3 cdac_ctrl_0.x1.X.n2 261.425
R13212 cdac_ctrl_0.x1.X cdac_ctrl_0.x1.X.n43 199.683
R13213 cdac_ctrl_0.x1.X.n3 cdac_ctrl_0.x1.X.n1 198.177
R13214 cdac_ctrl_0.x1.X.n4 cdac_ctrl_0.x1.X.n0 198.177
R13215 cdac_ctrl_0.x1.X.n32 cdac_ctrl_0.x1.X.n31 196.493
R13216 cdac_ctrl_0.x1.X.n29 cdac_ctrl_0.x1.X.n28 196.493
R13217 cdac_ctrl_0.x1.X.n26 cdac_ctrl_0.x1.X.n25 196.493
R13218 cdac_ctrl_0.x1.X.n23 cdac_ctrl_0.x1.X.n22 196.493
R13219 cdac_ctrl_0.x1.X.n20 cdac_ctrl_0.x1.X.n19 196.493
R13220 cdac_ctrl_0.x1.X.n17 cdac_ctrl_0.x1.X.n16 196.493
R13221 cdac_ctrl_0.x1.X.n14 cdac_ctrl_0.x1.X.n13 196.493
R13222 cdac_ctrl_0.x1.X.n11 cdac_ctrl_0.x1.X.n10 196.493
R13223 cdac_ctrl_0.x1.X.n8 cdac_ctrl_0.x1.X.n7 196.493
R13224 cdac_ctrl_0.x1.X.n6 cdac_ctrl_0.x1.X.n5 196.493
R13225 cdac_ctrl_0.x1.X.n4 cdac_ctrl_0.x1.X.n3 63.2476
R13226 cdac_ctrl_0.x1.X.n40 cdac_ctrl_0.x1.X.n39 63.2476
R13227 cdac_ctrl_0.x1.X.n42 cdac_ctrl_0.x1.X.n4 50.4476
R13228 cdac_ctrl_0.x1.X.n41 cdac_ctrl_0.x1.X.n40 50.4476
R13229 cdac_ctrl_0.x1.X.n9 cdac_ctrl_0.x1.X.n6 38.2063
R13230 cdac_ctrl_0.x1.X.n41 cdac_ctrl_0.x1.X.n35 31.7955
R13231 cdac_ctrl_0.x1.X.n15 cdac_ctrl_0.x1.X.n14 31.3559
R13232 cdac_ctrl_0.x1.X.n12 cdac_ctrl_0.x1.X.n11 31.3559
R13233 cdac_ctrl_0.x1.X.n33 cdac_ctrl_0.x1.X.n32 31.159
R13234 cdac_ctrl_0.x1.X.n30 cdac_ctrl_0.x1.X.n29 31.159
R13235 cdac_ctrl_0.x1.X.n27 cdac_ctrl_0.x1.X.n26 31.159
R13236 cdac_ctrl_0.x1.X.n24 cdac_ctrl_0.x1.X.n23 31.159
R13237 cdac_ctrl_0.x1.X.n21 cdac_ctrl_0.x1.X.n20 31.159
R13238 cdac_ctrl_0.x1.X.n18 cdac_ctrl_0.x1.X.n17 31.159
R13239 cdac_ctrl_0.x1.X.n9 cdac_ctrl_0.x1.X.n8 31.159
R13240 cdac_ctrl_0.x1.X.n35 cdac_ctrl_0.x1.X.n33 28.2061
R13241 cdac_ctrl_0.x1.X.n34 cdac_ctrl_0.x1.X.t10 26.5955
R13242 cdac_ctrl_0.x1.X.n34 cdac_ctrl_0.x1.X.t11 26.5955
R13243 cdac_ctrl_0.x1.X.n36 cdac_ctrl_0.x1.X.t8 26.5955
R13244 cdac_ctrl_0.x1.X.n36 cdac_ctrl_0.x1.X.t9 26.5955
R13245 cdac_ctrl_0.x1.X.n37 cdac_ctrl_0.x1.X.t12 26.5955
R13246 cdac_ctrl_0.x1.X.n37 cdac_ctrl_0.x1.X.t13 26.5955
R13247 cdac_ctrl_0.x1.X.n38 cdac_ctrl_0.x1.X.t14 26.5955
R13248 cdac_ctrl_0.x1.X.n38 cdac_ctrl_0.x1.X.t15 26.5955
R13249 cdac_ctrl_0.x1.X.n2 cdac_ctrl_0.x1.X.t4 24.9236
R13250 cdac_ctrl_0.x1.X.n2 cdac_ctrl_0.x1.X.t5 24.9236
R13251 cdac_ctrl_0.x1.X.n1 cdac_ctrl_0.x1.X.t6 24.9236
R13252 cdac_ctrl_0.x1.X.n1 cdac_ctrl_0.x1.X.t7 24.9236
R13253 cdac_ctrl_0.x1.X.n0 cdac_ctrl_0.x1.X.t0 24.9236
R13254 cdac_ctrl_0.x1.X.n0 cdac_ctrl_0.x1.X.t1 24.9236
R13255 cdac_ctrl_0.x1.X.n43 cdac_ctrl_0.x1.X.t2 24.9236
R13256 cdac_ctrl_0.x1.X.n43 cdac_ctrl_0.x1.X.t3 24.9236
R13257 cdac_ctrl_0.x1.X.n42 cdac_ctrl_0.x1.X 14.3064
R13258 cdac_ctrl_0.x1.X.n12 cdac_ctrl_0.x1.X.n9 7.04781
R13259 cdac_ctrl_0.x1.X.n15 cdac_ctrl_0.x1.X.n12 7.04781
R13260 cdac_ctrl_0.x1.X.n18 cdac_ctrl_0.x1.X.n15 7.04781
R13261 cdac_ctrl_0.x1.X.n21 cdac_ctrl_0.x1.X.n18 7.04781
R13262 cdac_ctrl_0.x1.X.n24 cdac_ctrl_0.x1.X.n21 7.04781
R13263 cdac_ctrl_0.x1.X.n27 cdac_ctrl_0.x1.X.n24 7.04781
R13264 cdac_ctrl_0.x1.X.n30 cdac_ctrl_0.x1.X.n27 7.04781
R13265 cdac_ctrl_0.x1.X.n33 cdac_ctrl_0.x1.X.n30 7.04781
R13266 cdac_ctrl_0.x1.X cdac_ctrl_0.x1.X.n41 4.26717
R13267 cdac_ctrl_0.x1.X cdac_ctrl_0.x1.X.n42 2.76128
R13268 cdac_ctrl_0.x1.X.n32 cdac_ctrl_0.x1.X 0.24431
R13269 cdac_ctrl_0.x1.X.n29 cdac_ctrl_0.x1.X 0.24431
R13270 cdac_ctrl_0.x1.X.n26 cdac_ctrl_0.x1.X 0.24431
R13271 cdac_ctrl_0.x1.X.n23 cdac_ctrl_0.x1.X 0.24431
R13272 cdac_ctrl_0.x1.X.n20 cdac_ctrl_0.x1.X 0.24431
R13273 cdac_ctrl_0.x1.X.n17 cdac_ctrl_0.x1.X 0.24431
R13274 cdac_ctrl_0.x1.X.n14 cdac_ctrl_0.x1.X 0.24431
R13275 cdac_ctrl_0.x1.X.n11 cdac_ctrl_0.x1.X 0.24431
R13276 cdac_ctrl_0.x1.X.n8 cdac_ctrl_0.x1.X 0.24431
R13277 cdac_ctrl_0.x1.X.n6 cdac_ctrl_0.x1.X 0.24431
R13278 a_n2412_n9650.n3 a_n2412_n9650.n2 636.953
R13279 a_n2412_n9650.n1 a_n2412_n9650.t4 366.856
R13280 a_n2412_n9650.n2 a_n2412_n9650.n0 300.2
R13281 a_n2412_n9650.n2 a_n2412_n9650.n1 225.036
R13282 a_n2412_n9650.n1 a_n2412_n9650.t5 174.056
R13283 a_n2412_n9650.n0 a_n2412_n9650.t3 70.0005
R13284 a_n2412_n9650.n3 a_n2412_n9650.t2 68.0124
R13285 a_n2412_n9650.t1 a_n2412_n9650.n3 63.3219
R13286 a_n2412_n9650.n0 a_n2412_n9650.t0 61.6672
R13287 a_n2058_n9662.t0 a_n2058_n9662.t1 87.1434
R13288 a_n2237_n9724.n4 a_n2237_n9724.n1 807.871
R13289 a_n2237_n9724.n0 a_n2237_n9724.t7 389.183
R13290 a_n2237_n9724.n5 a_n2237_n9724.n0 251.167
R13291 a_n2237_n9724.t0 a_n2237_n9724.n5 223.571
R13292 a_n2237_n9724.n2 a_n2237_n9724.t6 212.081
R13293 a_n2237_n9724.n3 a_n2237_n9724.t8 212.081
R13294 a_n2237_n9724.n4 a_n2237_n9724.n3 176.576
R13295 a_n2237_n9724.n0 a_n2237_n9724.t3 174.891
R13296 a_n2237_n9724.n2 a_n2237_n9724.t5 139.78
R13297 a_n2237_n9724.n3 a_n2237_n9724.t4 139.78
R13298 a_n2237_n9724.n1 a_n2237_n9724.t1 63.3219
R13299 a_n2237_n9724.n1 a_n2237_n9724.t2 63.3219
R13300 a_n2237_n9724.n3 a_n2237_n9724.n2 61.346
R13301 a_n2237_n9724.n5 a_n2237_n9724.n4 37.7195
R13302 a_n3327_n10022.t1 a_n3327_n10022.n3 370.026
R13303 a_n3327_n10022.n0 a_n3327_n10022.t5 351.356
R13304 a_n3327_n10022.n1 a_n3327_n10022.t3 334.717
R13305 a_n3327_n10022.n3 a_n3327_n10022.t0 325.971
R13306 a_n3327_n10022.n1 a_n3327_n10022.t4 309.935
R13307 a_n3327_n10022.n0 a_n3327_n10022.t2 305.683
R13308 a_n3327_n10022.n2 a_n3327_n10022.n0 16.879
R13309 a_n3327_n10022.n3 a_n3327_n10022.n2 10.8867
R13310 a_n3327_n10022.n2 a_n3327_n10022.n1 9.3005
R13311 a_n2250_n10028.t0 a_n2250_n10028.t1 126.644
R13312 a_7556_n5650.n5 a_7556_n5650.n4 807.871
R13313 a_7556_n5650.n0 a_7556_n5650.t3 389.183
R13314 a_7556_n5650.n1 a_7556_n5650.n0 251.167
R13315 a_7556_n5650.n1 a_7556_n5650.t1 223.571
R13316 a_7556_n5650.n3 a_7556_n5650.t7 212.081
R13317 a_7556_n5650.n2 a_7556_n5650.t8 212.081
R13318 a_7556_n5650.n4 a_7556_n5650.n3 176.576
R13319 a_7556_n5650.n0 a_7556_n5650.t6 174.891
R13320 a_7556_n5650.n3 a_7556_n5650.t4 139.78
R13321 a_7556_n5650.n2 a_7556_n5650.t5 139.78
R13322 a_7556_n5650.t0 a_7556_n5650.n5 63.3219
R13323 a_7556_n5650.n5 a_7556_n5650.t2 63.3219
R13324 a_7556_n5650.n3 a_7556_n5650.n2 61.346
R13325 a_7556_n5650.n4 a_7556_n5650.n1 37.5061
R13326 a_2670_2717.n3 a_2670_2717.n2 674.338
R13327 a_2670_2717.n1 a_2670_2717.t5 332.58
R13328 a_2670_2717.n2 a_2670_2717.n0 284.012
R13329 a_2670_2717.n2 a_2670_2717.n1 253.648
R13330 a_2670_2717.n1 a_2670_2717.t4 168.701
R13331 a_2670_2717.n3 a_2670_2717.t3 96.1553
R13332 a_2670_2717.t0 a_2670_2717.n3 65.6672
R13333 a_2670_2717.n0 a_2670_2717.t2 65.0005
R13334 a_2670_2717.n0 a_2670_2717.t1 45.0005
R13335 a_3558_n1029.t0 a_3558_n1029.t1 87.1434
R13336 a_191_n1029.n1 a_191_n1029.t3 530.01
R13337 a_191_n1029.t1 a_191_n1029.n5 421.021
R13338 a_191_n1029.n0 a_191_n1029.t2 337.142
R13339 a_191_n1029.n3 a_191_n1029.t0 280.223
R13340 a_191_n1029.n4 a_191_n1029.t7 263.173
R13341 a_191_n1029.n4 a_191_n1029.t6 227.826
R13342 a_191_n1029.n0 a_191_n1029.t5 199.762
R13343 a_191_n1029.n2 a_191_n1029.n1 170.81
R13344 a_191_n1029.n2 a_191_n1029.n0 167.321
R13345 a_191_n1029.n5 a_191_n1029.n4 152
R13346 a_191_n1029.n1 a_191_n1029.t4 141.923
R13347 a_191_n1029.n3 a_191_n1029.n2 10.8376
R13348 a_191_n1029.n5 a_191_n1029.n3 2.50485
R13349 a_925_n787.n3 a_925_n787.n2 647.119
R13350 a_925_n787.n1 a_925_n787.t4 350.253
R13351 a_925_n787.n2 a_925_n787.n0 260.339
R13352 a_925_n787.n2 a_925_n787.n1 246.119
R13353 a_925_n787.n1 a_925_n787.t5 189.588
R13354 a_925_n787.n3 a_925_n787.t0 89.1195
R13355 a_925_n787.n0 a_925_n787.t3 63.3338
R13356 a_925_n787.t2 a_925_n787.n3 41.0422
R13357 a_925_n787.n0 a_925_n787.t1 31.9797
R13358 a_1272_n1029.n3 a_1272_n1029.n2 636.953
R13359 a_1272_n1029.n1 a_1272_n1029.t5 366.856
R13360 a_1272_n1029.n2 a_1272_n1029.n0 300.2
R13361 a_1272_n1029.n2 a_1272_n1029.n1 225.036
R13362 a_1272_n1029.n1 a_1272_n1029.t4 174.056
R13363 a_1272_n1029.n0 a_1272_n1029.t3 70.0005
R13364 a_1272_n1029.t0 a_1272_n1029.n3 68.0124
R13365 a_1272_n1029.n3 a_1272_n1029.t2 63.3219
R13366 a_1272_n1029.n0 a_1272_n1029.t1 61.6672
R13367 a_3410_2691.n5 a_3410_2691.n4 807.871
R13368 a_3410_2691.n2 a_3410_2691.t6 389.183
R13369 a_3410_2691.n3 a_3410_2691.n2 251.167
R13370 a_3410_2691.n3 a_3410_2691.t1 223.571
R13371 a_3410_2691.n0 a_3410_2691.t7 212.081
R13372 a_3410_2691.n1 a_3410_2691.t3 212.081
R13373 a_3410_2691.n4 a_3410_2691.n1 176.576
R13374 a_3410_2691.n2 a_3410_2691.t5 174.891
R13375 a_3410_2691.n0 a_3410_2691.t8 139.78
R13376 a_3410_2691.n1 a_3410_2691.t4 139.78
R13377 a_3410_2691.t0 a_3410_2691.n5 63.3219
R13378 a_3410_2691.n5 a_3410_2691.t2 63.3219
R13379 a_3410_2691.n1 a_3410_2691.n0 61.346
R13380 a_3410_2691.n4 a_3410_2691.n3 37.7195
R13381 auto_sampling_0.x15.D.n5 auto_sampling_0.x15.D.n4 585
R13382 auto_sampling_0.x15.D.n4 auto_sampling_0.x15.D.n3 585
R13383 auto_sampling_0.x15.D.n2 auto_sampling_0.x15.D.t5 333.651
R13384 auto_sampling_0.x15.D.n2 auto_sampling_0.x15.D.t4 297.233
R13385 auto_sampling_0.x15.D auto_sampling_0.x15.D.n2 196.493
R13386 auto_sampling_0.x15.D.n1 auto_sampling_0.x15.D.n0 185
R13387 auto_sampling_0.x15.D auto_sampling_0.x15.D.n1 49.0339
R13388 auto_sampling_0.x15.D.n3 auto_sampling_0.x15.D 44.2533
R13389 auto_sampling_0.x15.D.n4 auto_sampling_0.x15.D.t2 26.5955
R13390 auto_sampling_0.x15.D.n4 auto_sampling_0.x15.D.t3 26.5955
R13391 auto_sampling_0.x15.D.n0 auto_sampling_0.x15.D.t0 24.9236
R13392 auto_sampling_0.x15.D.n0 auto_sampling_0.x15.D.t1 24.9236
R13393 auto_sampling_0.x15.D.n5 auto_sampling_0.x15.D 15.6165
R13394 auto_sampling_0.x15.D.n1 auto_sampling_0.x15.D 10.4965
R13395 auto_sampling_0.x15.D.n3 auto_sampling_0.x15.D 1.7925
R13396 auto_sampling_0.x15.D auto_sampling_0.x15.D.n5 1.7925
R13397 a_8116_2717.t1 a_8116_2717.n3 370.026
R13398 a_8116_2717.n0 a_8116_2717.t2 351.356
R13399 a_8116_2717.n1 a_8116_2717.t4 334.717
R13400 a_8116_2717.n3 a_8116_2717.t0 325.971
R13401 a_8116_2717.n1 a_8116_2717.t3 309.935
R13402 a_8116_2717.n0 a_8116_2717.t5 305.683
R13403 a_8116_2717.n2 a_8116_2717.n0 16.879
R13404 a_8116_2717.n3 a_8116_2717.n2 10.8867
R13405 a_8116_2717.n2 a_8116_2717.n1 9.3005
R13406 a_8684_2959.n3 a_8684_2959.n2 647.119
R13407 a_8684_2959.n1 a_8684_2959.t4 350.253
R13408 a_8684_2959.n2 a_8684_2959.n0 260.339
R13409 a_8684_2959.n2 a_8684_2959.n1 246.119
R13410 a_8684_2959.n1 a_8684_2959.t5 189.588
R13411 a_8684_2959.n3 a_8684_2959.t0 89.1195
R13412 a_8684_2959.n0 a_8684_2959.t3 63.3338
R13413 a_8684_2959.t2 a_8684_2959.n3 41.0422
R13414 a_8684_2959.n0 a_8684_2959.t1 31.9797
R13415 a_9031_2717.n3 a_9031_2717.n2 636.953
R13416 a_9031_2717.n1 a_9031_2717.t4 366.856
R13417 a_9031_2717.n2 a_9031_2717.n0 300.2
R13418 a_9031_2717.n2 a_9031_2717.n1 225.036
R13419 a_9031_2717.n1 a_9031_2717.t5 174.056
R13420 a_9031_2717.n0 a_9031_2717.t3 70.0005
R13421 a_9031_2717.t1 a_9031_2717.n3 68.0124
R13422 a_9031_2717.n3 a_9031_2717.t2 63.3219
R13423 a_9031_2717.n0 a_9031_2717.t0 61.6672
R13424 a_9534_n9484.t0 a_9534_n9484.t1 87.1434
R13425 a_9355_n9510.n3 a_9355_n9510.n0 807.871
R13426 a_9355_n9510.n4 a_9355_n9510.t4 389.183
R13427 a_9355_n9510.n5 a_9355_n9510.n4 251.167
R13428 a_9355_n9510.t0 a_9355_n9510.n5 223.571
R13429 a_9355_n9510.n1 a_9355_n9510.t6 212.081
R13430 a_9355_n9510.n2 a_9355_n9510.t8 212.081
R13431 a_9355_n9510.n3 a_9355_n9510.n2 176.576
R13432 a_9355_n9510.n4 a_9355_n9510.t3 174.891
R13433 a_9355_n9510.n1 a_9355_n9510.t5 139.78
R13434 a_9355_n9510.n2 a_9355_n9510.t7 139.78
R13435 a_9355_n9510.n0 a_9355_n9510.t1 63.3219
R13436 a_9355_n9510.n0 a_9355_n9510.t2 63.3219
R13437 a_9355_n9510.n2 a_9355_n9510.n1 61.346
R13438 a_9355_n9510.n5 a_9355_n9510.n3 37.7195
R13439 a_6535_3557.n3 a_6535_3557.n2 674.338
R13440 a_6535_3557.n1 a_6535_3557.t4 332.58
R13441 a_6535_3557.n2 a_6535_3557.n0 284.012
R13442 a_6535_3557.n2 a_6535_3557.n1 253.648
R13443 a_6535_3557.n1 a_6535_3557.t5 168.701
R13444 a_6535_3557.n3 a_6535_3557.t3 96.1553
R13445 a_6535_3557.t1 a_6535_3557.n3 65.6672
R13446 a_6535_3557.n0 a_6535_3557.t2 65.0005
R13447 a_6535_3557.n0 a_6535_3557.t0 45.0005
R13448 a_7248_n9650.n3 a_7248_n9650.n2 636.953
R13449 a_7248_n9650.n1 a_7248_n9650.t5 366.856
R13450 a_7248_n9650.n2 a_7248_n9650.n0 300.2
R13451 a_7248_n9650.n2 a_7248_n9650.n1 225.036
R13452 a_7248_n9650.n1 a_7248_n9650.t4 174.056
R13453 a_7248_n9650.n0 a_7248_n9650.t3 70.0005
R13454 a_7248_n9650.t0 a_7248_n9650.n3 68.0124
R13455 a_7248_n9650.n3 a_7248_n9650.t2 63.3219
R13456 a_7248_n9650.n0 a_7248_n9650.t1 61.6672
R13457 a_7357_n9650.n0 a_7357_n9650.t1 68.3338
R13458 a_7357_n9650.n0 a_7357_n9650.t0 26.3935
R13459 a_7357_n9650.n1 a_7357_n9650.n0 14.4005
R13460 a_9355_n9724.n5 a_9355_n9724.n4 807.871
R13461 a_9355_n9724.n2 a_9355_n9724.t8 389.183
R13462 a_9355_n9724.n3 a_9355_n9724.n2 251.167
R13463 a_9355_n9724.n3 a_9355_n9724.t1 223.571
R13464 a_9355_n9724.n0 a_9355_n9724.t5 212.081
R13465 a_9355_n9724.n1 a_9355_n9724.t3 212.081
R13466 a_9355_n9724.n4 a_9355_n9724.n1 176.576
R13467 a_9355_n9724.n2 a_9355_n9724.t7 174.891
R13468 a_9355_n9724.n0 a_9355_n9724.t4 139.78
R13469 a_9355_n9724.n1 a_9355_n9724.t6 139.78
R13470 a_9355_n9724.t0 a_9355_n9724.n5 63.3219
R13471 a_9355_n9724.n5 a_9355_n9724.t2 63.3219
R13472 a_9355_n9724.n1 a_9355_n9724.n0 61.346
R13473 a_9355_n9724.n4 a_9355_n9724.n3 37.7195
R13474 SWN[9].n4 SWN[9].n3 585
R13475 SWN[9].n3 SWN[9].n2 585
R13476 SWN[9].n1 SWN[9].n0 185
R13477 SWN[9].n5 SWN[9].n1 53.3859
R13478 SWN[9].n3 SWN[9].t2 26.5955
R13479 SWN[9].n3 SWN[9].t3 26.5955
R13480 SWN[9].n0 SWN[9].t1 24.9236
R13481 SWN[9].n0 SWN[9].t0 24.9236
R13482 SWN[9] SWN[9].n5 14.6674
R13483 SWN[9] SWN[9].n4 10.4965
R13484 SWN[9].n2 SWN[9] 10.4965
R13485 SWN[9].n4 SWN[9] 6.9125
R13486 SWN[9].n2 SWN[9] 6.9125
R13487 SWN[9].n5 SWN[9] 4.3525
R13488 SWN[9].n1 SWN[9] 1.7925
R13489 a_1658_3557.t0 a_1658_3557.t1 87.1434
R13490 a_8833_n10054.n3 a_8833_n10054.n2 647.119
R13491 a_8833_n10054.n1 a_8833_n10054.t5 350.253
R13492 a_8833_n10054.n2 a_8833_n10054.n0 260.339
R13493 a_8833_n10054.n2 a_8833_n10054.n1 246.119
R13494 a_8833_n10054.n1 a_8833_n10054.t4 189.588
R13495 a_8833_n10054.n3 a_8833_n10054.t0 89.1195
R13496 a_8833_n10054.n0 a_8833_n10054.t1 63.3338
R13497 a_8833_n10054.t3 a_8833_n10054.n3 41.0422
R13498 a_8833_n10054.n0 a_8833_n10054.t2 31.9797
R13499 a_3088_n1573.n0 a_3088_n1573.t2 1327.82
R13500 a_3088_n1573.t0 a_3088_n1573.n0 194.655
R13501 a_3088_n1573.n0 a_3088_n1573.t1 63.3219
R13502 a_2943_n1599.n3 a_2943_n1599.n2 674.338
R13503 a_2943_n1599.n1 a_2943_n1599.t5 332.58
R13504 a_2943_n1599.n2 a_2943_n1599.n0 284.012
R13505 a_2943_n1599.n2 a_2943_n1599.n1 253.648
R13506 a_2943_n1599.n1 a_2943_n1599.t4 168.701
R13507 a_2943_n1599.t1 a_2943_n1599.n3 96.1553
R13508 a_2943_n1599.n3 a_2943_n1599.t3 65.6672
R13509 a_2943_n1599.n0 a_2943_n1599.t0 65.0005
R13510 a_2943_n1599.n0 a_2943_n1599.t2 45.0005
R13511 a_n6841_n9650.n3 a_n6841_n9650.n2 674.338
R13512 a_n6841_n9650.n1 a_n6841_n9650.t5 332.58
R13513 a_n6841_n9650.n2 a_n6841_n9650.n0 284.012
R13514 a_n6841_n9650.n2 a_n6841_n9650.n1 253.648
R13515 a_n6841_n9650.n1 a_n6841_n9650.t4 168.701
R13516 a_n6841_n9650.n3 a_n6841_n9650.t3 96.1553
R13517 a_n6841_n9650.t0 a_n6841_n9650.n3 65.6672
R13518 a_n6841_n9650.n0 a_n6841_n9650.t2 65.0005
R13519 a_n6841_n9650.n0 a_n6841_n9650.t1 45.0005
R13520 a_n6623_n10054.n3 a_n6623_n10054.n2 647.119
R13521 a_n6623_n10054.n1 a_n6623_n10054.t4 350.253
R13522 a_n6623_n10054.n2 a_n6623_n10054.n0 260.339
R13523 a_n6623_n10054.n2 a_n6623_n10054.n1 246.119
R13524 a_n6623_n10054.n1 a_n6623_n10054.t5 189.588
R13525 a_n6623_n10054.n3 a_n6623_n10054.t3 89.1195
R13526 a_n6623_n10054.n0 a_n6623_n10054.t2 63.3338
R13527 a_n6623_n10054.t1 a_n6623_n10054.n3 41.0422
R13528 a_n6623_n10054.n0 a_n6623_n10054.t0 31.9797
R13529 a_9207_3531.n5 a_9207_3531.n4 807.871
R13530 a_9207_3531.n2 a_9207_3531.t3 389.183
R13531 a_9207_3531.n3 a_9207_3531.n2 251.167
R13532 a_9207_3531.n3 a_9207_3531.t2 223.571
R13533 a_9207_3531.n0 a_9207_3531.t4 212.081
R13534 a_9207_3531.n1 a_9207_3531.t8 212.081
R13535 a_9207_3531.n4 a_9207_3531.n1 176.576
R13536 a_9207_3531.n2 a_9207_3531.t5 174.891
R13537 a_9207_3531.n0 a_9207_3531.t7 139.78
R13538 a_9207_3531.n1 a_9207_3531.t6 139.78
R13539 a_9207_3531.n5 a_9207_3531.t1 63.3219
R13540 a_9207_3531.t0 a_9207_3531.n5 63.3219
R13541 a_9207_3531.n1 a_9207_3531.n0 61.346
R13542 a_9207_3531.n4 a_9207_3531.n3 37.7195
R13543 a_4115_n1599.n5 a_4115_n1599.n4 807.871
R13544 a_4115_n1599.n0 a_4115_n1599.t6 389.183
R13545 a_4115_n1599.n1 a_4115_n1599.n0 251.167
R13546 a_4115_n1599.n1 a_4115_n1599.t2 223.571
R13547 a_4115_n1599.n3 a_4115_n1599.t4 212.081
R13548 a_4115_n1599.n2 a_4115_n1599.t5 212.081
R13549 a_4115_n1599.n4 a_4115_n1599.n3 176.576
R13550 a_4115_n1599.n0 a_4115_n1599.t3 174.891
R13551 a_4115_n1599.n3 a_4115_n1599.t7 139.78
R13552 a_4115_n1599.n2 a_4115_n1599.t8 139.78
R13553 a_4115_n1599.t0 a_4115_n1599.n5 63.3219
R13554 a_4115_n1599.n5 a_4115_n1599.t1 63.3219
R13555 a_4115_n1599.n3 a_4115_n1599.n2 61.346
R13556 a_4115_n1599.n4 a_4115_n1599.n1 37.5061
R13557 a_4677_n1207.t1 a_4677_n1207.t0 94.7268
R13558 a_251_n1599.n4 a_251_n1599.n1 807.871
R13559 a_251_n1599.n0 a_251_n1599.t3 389.183
R13560 a_251_n1599.n5 a_251_n1599.n0 251.167
R13561 a_251_n1599.t0 a_251_n1599.n5 223.571
R13562 a_251_n1599.n3 a_251_n1599.t8 212.081
R13563 a_251_n1599.n2 a_251_n1599.t7 212.081
R13564 a_251_n1599.n4 a_251_n1599.n3 176.576
R13565 a_251_n1599.n0 a_251_n1599.t5 174.891
R13566 a_251_n1599.n3 a_251_n1599.t6 139.78
R13567 a_251_n1599.n2 a_251_n1599.t4 139.78
R13568 a_251_n1599.n1 a_251_n1599.t2 63.3219
R13569 a_251_n1599.n1 a_251_n1599.t1 63.3219
R13570 a_251_n1599.n3 a_251_n1599.n2 61.346
R13571 a_251_n1599.n5 a_251_n1599.n4 37.5061
R13572 a_772_n1573.t0 a_772_n1573.t1 126.644
R13573 a_537_n9484.t1 a_537_n9484.n3 370.026
R13574 a_537_n9484.n0 a_537_n9484.t5 351.356
R13575 a_537_n9484.n1 a_537_n9484.t3 334.717
R13576 a_537_n9484.n3 a_537_n9484.t0 325.971
R13577 a_537_n9484.n1 a_537_n9484.t4 309.935
R13578 a_537_n9484.n0 a_537_n9484.t2 305.683
R13579 a_537_n9484.n2 a_537_n9484.n0 16.879
R13580 a_537_n9484.n3 a_537_n9484.n2 10.8867
R13581 a_537_n9484.n2 a_537_n9484.n1 9.3005
R13582 a_1452_n9484.n3 a_1452_n9484.n2 636.953
R13583 a_1452_n9484.n1 a_1452_n9484.t4 366.856
R13584 a_1452_n9484.n2 a_1452_n9484.n0 300.2
R13585 a_1452_n9484.n2 a_1452_n9484.n1 225.036
R13586 a_1452_n9484.n1 a_1452_n9484.t5 174.056
R13587 a_1452_n9484.n0 a_1452_n9484.t3 70.0005
R13588 a_1452_n9484.t1 a_1452_n9484.n3 68.0124
R13589 a_1452_n9484.n3 a_1452_n9484.t2 63.3219
R13590 a_1452_n9484.n0 a_1452_n9484.t0 61.6672
R13591 a_1614_n9118.t0 a_1614_n9118.t1 126.644
R13592 a_4719_n1331.n1 a_4719_n1331.t3 530.01
R13593 a_4719_n1331.t1 a_4719_n1331.n5 421.021
R13594 a_4719_n1331.n0 a_4719_n1331.t7 337.171
R13595 a_4719_n1331.n3 a_4719_n1331.t0 280.223
R13596 a_4719_n1331.n4 a_4719_n1331.t5 263.173
R13597 a_4719_n1331.n4 a_4719_n1331.t4 227.826
R13598 a_4719_n1331.n0 a_4719_n1331.t2 199.762
R13599 a_4719_n1331.n2 a_4719_n1331.n1 170.81
R13600 a_4719_n1331.n2 a_4719_n1331.n0 167.321
R13601 a_4719_n1331.n5 a_4719_n1331.n4 152
R13602 a_4719_n1331.n1 a_4719_n1331.t6 141.923
R13603 a_4719_n1331.n3 a_4719_n1331.n2 10.8376
R13604 a_4719_n1331.n5 a_4719_n1331.n3 2.50485
R13605 a_n467_3083.t0 a_n467_3083.t1 126.644
R13606 a_3559_n9510.n5 a_3559_n9510.n4 807.871
R13607 a_3559_n9510.n2 a_3559_n9510.t3 389.183
R13608 a_3559_n9510.n3 a_3559_n9510.n2 251.167
R13609 a_3559_n9510.n3 a_3559_n9510.t1 223.571
R13610 a_3559_n9510.n0 a_3559_n9510.t7 212.081
R13611 a_3559_n9510.n1 a_3559_n9510.t5 212.081
R13612 a_3559_n9510.n4 a_3559_n9510.n1 176.576
R13613 a_3559_n9510.n2 a_3559_n9510.t8 174.891
R13614 a_3559_n9510.n0 a_3559_n9510.t6 139.78
R13615 a_3559_n9510.n1 a_3559_n9510.t4 139.78
R13616 a_3559_n9510.t0 a_3559_n9510.n5 63.3219
R13617 a_3559_n9510.n5 a_3559_n9510.t2 63.3219
R13618 a_3559_n9510.n1 a_3559_n9510.n0 61.346
R13619 a_3559_n9510.n4 a_3559_n9510.n3 37.7195
R13620 a_3546_n9118.t0 a_3546_n9118.t1 126.644
R13621 a_n9289_n9484.n1 a_n9289_n9484.t6 530.01
R13622 a_n9289_n9484.t1 a_n9289_n9484.n5 421.021
R13623 a_n9289_n9484.n0 a_n9289_n9484.t7 337.142
R13624 a_n9289_n9484.n3 a_n9289_n9484.t0 280.223
R13625 a_n9289_n9484.n4 a_n9289_n9484.t3 263.173
R13626 a_n9289_n9484.n4 a_n9289_n9484.t5 227.826
R13627 a_n9289_n9484.n0 a_n9289_n9484.t4 199.762
R13628 a_n9289_n9484.n2 a_n9289_n9484.n1 170.81
R13629 a_n9289_n9484.n2 a_n9289_n9484.n0 167.321
R13630 a_n9289_n9484.n5 a_n9289_n9484.n4 152
R13631 a_n9289_n9484.n1 a_n9289_n9484.t2 141.923
R13632 a_n9289_n9484.n3 a_n9289_n9484.n2 10.8376
R13633 a_n9289_n9484.n5 a_n9289_n9484.n3 2.50485
R13634 a_n8868_n9484.n1 a_n8868_n9484.n0 926.024
R13635 a_n8868_n9484.t1 a_n8868_n9484.n1 82.0838
R13636 a_n8868_n9484.n0 a_n8868_n9484.t0 63.3338
R13637 a_n8868_n9484.n1 a_n8868_n9484.t3 63.3219
R13638 a_n8868_n9484.n0 a_n8868_n9484.t2 29.7268
R13639 a_1011_n1599.n3 a_1011_n1599.n2 674.338
R13640 a_1011_n1599.n1 a_1011_n1599.t5 332.58
R13641 a_1011_n1599.n2 a_1011_n1599.n0 284.012
R13642 a_1011_n1599.n2 a_1011_n1599.n1 253.648
R13643 a_1011_n1599.n1 a_1011_n1599.t4 168.701
R13644 a_1011_n1599.n3 a_1011_n1599.t2 96.1553
R13645 a_1011_n1599.t0 a_1011_n1599.n3 65.6672
R13646 a_1011_n1599.n0 a_1011_n1599.t3 65.0005
R13647 a_1011_n1599.n0 a_1011_n1599.t1 45.0005
R13648 a_1574_n1573.n1 a_1574_n1573.n0 926.024
R13649 a_1574_n1573.t0 a_1574_n1573.n1 82.0838
R13650 a_1574_n1573.n0 a_1574_n1573.t3 63.3338
R13651 a_1574_n1573.n1 a_1574_n1573.t1 63.3219
R13652 a_1574_n1573.n0 a_1574_n1573.t2 29.7268
R13653 a_8739_n5080.t0 a_8739_n5080.t1 126.644
R13654 a_n9289_n10022.n1 a_n9289_n10022.t3 530.01
R13655 a_n9289_n10022.t0 a_n9289_n10022.n5 421.021
R13656 a_n9289_n10022.n0 a_n9289_n10022.t4 337.142
R13657 a_n9289_n10022.n3 a_n9289_n10022.t1 280.223
R13658 a_n9289_n10022.n4 a_n9289_n10022.t5 263.173
R13659 a_n9289_n10022.n4 a_n9289_n10022.t7 227.826
R13660 a_n9289_n10022.n0 a_n9289_n10022.t2 199.762
R13661 a_n9289_n10022.n2 a_n9289_n10022.n1 170.81
R13662 a_n9289_n10022.n2 a_n9289_n10022.n0 167.321
R13663 a_n9289_n10022.n5 a_n9289_n10022.n4 152
R13664 a_n9289_n10022.n1 a_n9289_n10022.t6 141.923
R13665 a_n9289_n10022.n3 a_n9289_n10022.n2 10.8376
R13666 a_n9289_n10022.n5 a_n9289_n10022.n3 2.50485
R13667 a_n8099_n9650.n0 a_n8099_n9650.t0 68.3338
R13668 a_n8099_n9650.n0 a_n8099_n9650.t1 26.3935
R13669 a_n8099_n9650.n1 a_n8099_n9650.n0 14.4005
R13670 a_6503_n1029.n3 a_6503_n1029.n2 674.338
R13671 a_6503_n1029.n1 a_6503_n1029.t5 332.58
R13672 a_6503_n1029.n2 a_6503_n1029.n0 284.012
R13673 a_6503_n1029.n2 a_6503_n1029.n1 253.648
R13674 a_6503_n1029.n1 a_6503_n1029.t4 168.701
R13675 a_6503_n1029.n3 a_6503_n1029.t3 96.1553
R13676 a_6503_n1029.t1 a_6503_n1029.n3 65.6672
R13677 a_6503_n1029.n0 a_6503_n1029.t2 65.0005
R13678 a_6503_n1029.n0 a_6503_n1029.t0 45.0005
R13679 a_1105_n9242.n3 a_1105_n9242.n2 647.119
R13680 a_1105_n9242.n1 a_1105_n9242.t5 350.253
R13681 a_1105_n9242.n2 a_1105_n9242.n0 260.339
R13682 a_1105_n9242.n2 a_1105_n9242.n1 246.119
R13683 a_1105_n9242.n1 a_1105_n9242.t4 189.588
R13684 a_1105_n9242.n3 a_1105_n9242.t0 89.1195
R13685 a_1105_n9242.n0 a_1105_n9242.t3 63.3338
R13686 a_1105_n9242.t2 a_1105_n9242.n3 41.0422
R13687 a_1105_n9242.n0 a_1105_n9242.t1 31.9797
R13688 a_546_n4714.t0 a_546_n4714.t1 60.0005
R13689 a_9162_n663.t0 a_9162_n663.t1 126.644
R13690 a_942_n1573.n3 a_942_n1573.n2 647.119
R13691 a_942_n1573.n1 a_942_n1573.t4 350.253
R13692 a_942_n1573.n2 a_942_n1573.n0 260.339
R13693 a_942_n1573.n2 a_942_n1573.n1 246.119
R13694 a_942_n1573.n1 a_942_n1573.t5 189.588
R13695 a_942_n1573.n3 a_942_n1573.t1 89.1195
R13696 a_942_n1573.n0 a_942_n1573.t0 63.3338
R13697 a_942_n1573.t3 a_942_n1573.n3 41.0422
R13698 a_942_n1573.n0 a_942_n1573.t2 31.9797
R13699 a_1249_n1207.t0 a_1249_n1207.t1 60.0005
R13700 a_1321_n1207.t1 a_1321_n1207.t0 198.571
R13701 a_6188_n5080.t0 a_6188_n5080.n0 1327.82
R13702 a_6188_n5080.n0 a_6188_n5080.t1 194.655
R13703 a_6188_n5080.n0 a_6188_n5080.t2 63.3219
R13704 DOUT[9].n3 DOUT[9].n2 585
R13705 DOUT[9].n4 DOUT[9].n3 585
R13706 DOUT[9].n1 DOUT[9].n0 185
R13707 DOUT[9] DOUT[9].n1 57.7379
R13708 DOUT[9].n3 DOUT[9].t3 26.5955
R13709 DOUT[9].n3 DOUT[9].t2 26.5955
R13710 DOUT[9].n0 DOUT[9].t1 24.9236
R13711 DOUT[9].n0 DOUT[9].t0 24.9236
R13712 DOUT[9] DOUT[9].n5 17.8815
R13713 DOUT[9].n2 DOUT[9] 10.4965
R13714 DOUT[9].n4 DOUT[9] 10.4965
R13715 DOUT[9].n2 DOUT[9] 6.9125
R13716 DOUT[9].n5 DOUT[9] 4.3525
R13717 DOUT[9].n5 DOUT[9].n4 2.5605
R13718 DOUT[9].n1 DOUT[9] 1.7925
R13719 a_7370_n1573.n1 a_7370_n1573.n0 926.024
R13720 a_7370_n1573.n0 a_7370_n1573.t3 82.0838
R13721 a_7370_n1573.n1 a_7370_n1573.t0 63.3338
R13722 a_7370_n1573.n0 a_7370_n1573.t2 63.3219
R13723 a_7370_n1573.n2 a_7370_n1573.t1 26.3935
R13724 a_7370_n1573.n3 a_7370_n1573.n2 14.4005
R13725 a_7370_n1573.n2 a_7370_n1573.n1 3.33383
R13726 a_n2977_n9484.n3 a_n2977_n9484.n2 674.338
R13727 a_n2977_n9484.n1 a_n2977_n9484.t5 332.58
R13728 a_n2977_n9484.n2 a_n2977_n9484.n0 284.012
R13729 a_n2977_n9484.n2 a_n2977_n9484.n1 253.648
R13730 a_n2977_n9484.n1 a_n2977_n9484.t4 168.701
R13731 a_n2977_n9484.n3 a_n2977_n9484.t3 96.1553
R13732 a_n2977_n9484.t2 a_n2977_n9484.n3 65.6672
R13733 a_n2977_n9484.n0 a_n2977_n9484.t0 65.0005
R13734 a_n2977_n9484.n0 a_n2977_n9484.t1 45.0005
R13735 a_n2759_n9242.n3 a_n2759_n9242.n2 647.119
R13736 a_n2759_n9242.n1 a_n2759_n9242.t5 350.253
R13737 a_n2759_n9242.n2 a_n2759_n9242.n0 260.339
R13738 a_n2759_n9242.n2 a_n2759_n9242.n1 246.119
R13739 a_n2759_n9242.n1 a_n2759_n9242.t4 189.588
R13740 a_n2759_n9242.n3 a_n2759_n9242.t1 89.1195
R13741 a_n2759_n9242.n0 a_n2759_n9242.t0 63.3338
R13742 a_n2759_n9242.t3 a_n2759_n9242.n3 41.0422
R13743 a_n2759_n9242.n0 a_n2759_n9242.t2 31.9797
R13744 a_n6101_n9510.n5 a_n6101_n9510.n4 807.871
R13745 a_n6101_n9510.n2 a_n6101_n9510.t8 389.183
R13746 a_n6101_n9510.n3 a_n6101_n9510.n2 251.167
R13747 a_n6101_n9510.n3 a_n6101_n9510.t1 223.571
R13748 a_n6101_n9510.n0 a_n6101_n9510.t6 212.081
R13749 a_n6101_n9510.n1 a_n6101_n9510.t4 212.081
R13750 a_n6101_n9510.n4 a_n6101_n9510.n1 176.576
R13751 a_n6101_n9510.n2 a_n6101_n9510.t7 174.891
R13752 a_n6101_n9510.n0 a_n6101_n9510.t5 139.78
R13753 a_n6101_n9510.n1 a_n6101_n9510.t3 139.78
R13754 a_n6101_n9510.n5 a_n6101_n9510.t2 63.3219
R13755 a_n6101_n9510.t0 a_n6101_n9510.n5 63.3219
R13756 a_n6101_n9510.n1 a_n6101_n9510.n0 61.346
R13757 a_n6101_n9510.n4 a_n6101_n9510.n3 37.7195
R13758 SWP[1].n0 SWP[1].t4 333.651
R13759 SWP[1].n0 SWP[1].t5 297.233
R13760 SWP[1].n5 SWP[1].n4 289.096
R13761 SWP[1].n1 SWP[1].n0 196.493
R13762 SWP[1].n7 SWP[1].n6 185
R13763 SWP[1].n3 SWP[1] 52.0428
R13764 SWP[1] SWP[1].n7 49.0339
R13765 SWP[1].n2 SWP[1].n1 39.5123
R13766 SWP[1].n4 SWP[1].t2 26.5955
R13767 SWP[1].n4 SWP[1].t3 26.5955
R13768 SWP[1].n6 SWP[1].t0 24.9236
R13769 SWP[1].n6 SWP[1].t1 24.9236
R13770 SWP[1] SWP[1].n3 19.0876
R13771 SWP[1] SWP[1].n8 14.6049
R13772 SWP[1].n8 SWP[1] 13.0565
R13773 SWP[1].n3 SWP[1].n2 11.4605
R13774 SWP[1].n7 SWP[1] 10.4965
R13775 SWP[1] SWP[1].n5 9.48653
R13776 SWP[1].n5 SWP[1] 7.7181
R13777 SWP[1].n8 SWP[1] 4.3525
R13778 SWP[1].n1 SWP[1] 0.24431
R13779 SWP[1].n2 SWP[1] 0.0022625
R13780 a_n6623_n9242.n3 a_n6623_n9242.n2 647.119
R13781 a_n6623_n9242.n1 a_n6623_n9242.t5 350.253
R13782 a_n6623_n9242.n2 a_n6623_n9242.n0 260.339
R13783 a_n6623_n9242.n2 a_n6623_n9242.n1 246.119
R13784 a_n6623_n9242.n1 a_n6623_n9242.t4 189.588
R13785 a_n6623_n9242.n3 a_n6623_n9242.t0 89.1195
R13786 a_n6623_n9242.n0 a_n6623_n9242.t3 63.3338
R13787 a_n6623_n9242.t2 a_n6623_n9242.n3 41.0422
R13788 a_n6623_n9242.n0 a_n6623_n9242.t1 31.9797
R13789 a_5670_n9662.t0 a_5670_n9662.t1 87.1434
R13790 a_1203_n4714.t0 a_1203_n4714.t1 87.1434
R13791 a_8723_n10028.n0 a_8723_n10028.t2 1327.82
R13792 a_8723_n10028.t0 a_8723_n10028.n0 194.655
R13793 a_8723_n10028.n0 a_8723_n10028.t1 63.3219
R13794 auto_sampling_0.x11.D.n5 auto_sampling_0.x11.D.n4 585
R13795 auto_sampling_0.x11.D.n4 auto_sampling_0.x11.D.n3 585
R13796 auto_sampling_0.x11.D.n2 auto_sampling_0.x11.D.t4 333.651
R13797 auto_sampling_0.x11.D.n2 auto_sampling_0.x11.D.t5 297.233
R13798 auto_sampling_0.x11.D auto_sampling_0.x11.D.n2 196.493
R13799 auto_sampling_0.x11.D.n1 auto_sampling_0.x11.D.n0 185
R13800 auto_sampling_0.x11.D auto_sampling_0.x11.D.n1 49.0339
R13801 auto_sampling_0.x11.D.n3 auto_sampling_0.x11.D 44.2533
R13802 auto_sampling_0.x11.D.n4 auto_sampling_0.x11.D.t2 26.5955
R13803 auto_sampling_0.x11.D.n4 auto_sampling_0.x11.D.t3 26.5955
R13804 auto_sampling_0.x11.D.n0 auto_sampling_0.x11.D.t1 24.9236
R13805 auto_sampling_0.x11.D.n0 auto_sampling_0.x11.D.t0 24.9236
R13806 auto_sampling_0.x11.D.n5 auto_sampling_0.x11.D 15.6165
R13807 auto_sampling_0.x11.D.n1 auto_sampling_0.x11.D 10.4965
R13808 auto_sampling_0.x11.D.n3 auto_sampling_0.x11.D 1.7925
R13809 auto_sampling_0.x11.D auto_sampling_0.x11.D.n5 1.7925
R13810 a_n4169_n9510.n3 a_n4169_n9510.n0 807.871
R13811 a_n4169_n9510.n4 a_n4169_n9510.t3 389.183
R13812 a_n4169_n9510.n5 a_n4169_n9510.n4 251.167
R13813 a_n4169_n9510.t0 a_n4169_n9510.n5 223.571
R13814 a_n4169_n9510.n1 a_n4169_n9510.t7 212.081
R13815 a_n4169_n9510.n2 a_n4169_n9510.t5 212.081
R13816 a_n4169_n9510.n3 a_n4169_n9510.n2 176.576
R13817 a_n4169_n9510.n4 a_n4169_n9510.t8 174.891
R13818 a_n4169_n9510.n1 a_n4169_n9510.t6 139.78
R13819 a_n4169_n9510.n2 a_n4169_n9510.t4 139.78
R13820 a_n4169_n9510.n0 a_n4169_n9510.t1 63.3219
R13821 a_n4169_n9510.n0 a_n4169_n9510.t2 63.3219
R13822 a_n4169_n9510.n2 a_n4169_n9510.n1 61.346
R13823 a_n4169_n9510.n5 a_n4169_n9510.n3 37.7195
R13824 CF[7].n11 CF[7].n10 585
R13825 CF[7].n12 CF[7].n11 585
R13826 CF[7].n6 CF[7].t9 333.651
R13827 CF[7].n6 CF[7].t5 297.233
R13828 CF[7].n3 CF[7].t7 294.557
R13829 CF[7].n0 CF[7].t8 294.557
R13830 CF[7].n3 CF[7].t6 211.01
R13831 CF[7].n0 CF[7].t4 211.01
R13832 CF[7].n7 CF[7].n6 196.493
R13833 CF[7].n9 CF[7].n8 185
R13834 CF[7].n4 CF[7].n3 153.097
R13835 CF[7].n1 CF[7].n0 152
R13836 CF[7] CF[7].n9 49.0339
R13837 CF[7] CF[7].n14 45.4935
R13838 CF[7].n13 CF[7].n7 35.37
R13839 CF[7].n11 CF[7].t3 26.5955
R13840 CF[7].n11 CF[7].t2 26.5955
R13841 CF[7].n14 CF[7] 25.3611
R13842 CF[7].n8 CF[7].t1 24.9236
R13843 CF[7].n8 CF[7].t0 24.9236
R13844 CF[7].n13 CF[7].n12 17.2879
R13845 CF[7].n10 CF[7] 15.6165
R13846 CF[7].n5 CF[7].n2 14.9321
R13847 CF[7].n5 CF[7].n4 13.9063
R13848 CF[7].n9 CF[7] 10.4965
R13849 CF[7].n2 CF[7] 9.32621
R13850 CF[7].n14 CF[7] 5.77425
R13851 CF[7].n4 CF[7] 3.10907
R13852 CF[7].n1 CF[7] 2.01193
R13853 CF[7].n12 CF[7] 1.7925
R13854 CF[7].n10 CF[7] 1.7925
R13855 CF[7].n2 CF[7].n1 1.09764
R13856 CF[7] CF[7].n5 0.851793
R13857 CF[7] CF[7].n13 0.740885
R13858 CF[7].n7 CF[7] 0.24431
R13859 DOUT[8].n3 DOUT[8].n2 585
R13860 DOUT[8].n4 DOUT[8].n3 585
R13861 DOUT[8].n1 DOUT[8].n0 185
R13862 DOUT[8] DOUT[8].n1 49.0339
R13863 DOUT[8].n3 DOUT[8].t3 26.5955
R13864 DOUT[8].n3 DOUT[8].t2 26.5955
R13865 DOUT[8].n0 DOUT[8].t1 24.9236
R13866 DOUT[8].n0 DOUT[8].t0 24.9236
R13867 DOUT[8] DOUT[8].n4 20.4383
R13868 DOUT[8].n2 DOUT[8] 15.6165
R13869 DOUT[8].n1 DOUT[8] 10.4965
R13870 DOUT[8].n4 DOUT[8] 1.7925
R13871 DOUT[8].n2 DOUT[8] 1.7925
R13872 a_2469_n10022.t1 a_2469_n10022.n3 370.026
R13873 a_2469_n10022.n0 a_2469_n10022.t3 351.356
R13874 a_2469_n10022.n1 a_2469_n10022.t5 334.717
R13875 a_2469_n10022.n3 a_2469_n10022.t0 325.971
R13876 a_2469_n10022.n1 a_2469_n10022.t4 309.935
R13877 a_2469_n10022.n0 a_2469_n10022.t2 305.683
R13878 a_2469_n10022.n2 a_2469_n10022.n0 16.879
R13879 a_2469_n10022.n3 a_2469_n10022.n2 10.8867
R13880 a_2469_n10022.n2 a_2469_n10022.n1 9.3005
R13881 a_3384_n9650.n3 a_3384_n9650.n2 636.953
R13882 a_3384_n9650.n1 a_3384_n9650.t4 366.856
R13883 a_3384_n9650.n2 a_3384_n9650.n0 300.2
R13884 a_3384_n9650.n2 a_3384_n9650.n1 225.036
R13885 a_3384_n9650.n1 a_3384_n9650.t5 174.056
R13886 a_3384_n9650.n0 a_3384_n9650.t2 70.0005
R13887 a_3384_n9650.t0 a_3384_n9650.n3 68.0124
R13888 a_3384_n9650.n3 a_3384_n9650.t3 63.3219
R13889 a_3384_n9650.n0 a_3384_n9650.t1 61.6672
R13890 a_3546_n10028.t0 a_3546_n10028.t1 126.644
R13891 a_n453_3531.n5 a_n453_3531.n4 807.871
R13892 a_n453_3531.n2 a_n453_3531.t5 389.183
R13893 a_n453_3531.n3 a_n453_3531.n2 251.167
R13894 a_n453_3531.n3 a_n453_3531.t1 223.571
R13895 a_n453_3531.n0 a_n453_3531.t6 212.081
R13896 a_n453_3531.n1 a_n453_3531.t8 212.081
R13897 a_n453_3531.n4 a_n453_3531.n1 176.576
R13898 a_n453_3531.n2 a_n453_3531.t7 174.891
R13899 a_n453_3531.n0 a_n453_3531.t3 139.78
R13900 a_n453_3531.n1 a_n453_3531.t4 139.78
R13901 a_n453_3531.n5 a_n453_3531.t2 63.3219
R13902 a_n453_3531.t0 a_n453_3531.n5 63.3219
R13903 a_n453_3531.n1 a_n453_3531.n0 61.346
R13904 a_n453_3531.n4 a_n453_3531.n3 37.7195
R13905 a_n6114_n10028.t0 a_n6114_n10028.t1 126.644
R13906 a_n3493_n10022.n1 a_n3493_n10022.t7 530.01
R13907 a_n3493_n10022.t1 a_n3493_n10022.n5 421.021
R13908 a_n3493_n10022.n0 a_n3493_n10022.t2 337.142
R13909 a_n3493_n10022.n3 a_n3493_n10022.t0 280.223
R13910 a_n3493_n10022.n4 a_n3493_n10022.t3 263.173
R13911 a_n3493_n10022.n4 a_n3493_n10022.t5 227.826
R13912 a_n3493_n10022.n0 a_n3493_n10022.t6 199.762
R13913 a_n3493_n10022.n2 a_n3493_n10022.n1 170.81
R13914 a_n3493_n10022.n2 a_n3493_n10022.n0 167.321
R13915 a_n3493_n10022.n5 a_n3493_n10022.n4 152
R13916 a_n3493_n10022.n1 a_n3493_n10022.t4 141.923
R13917 a_n3493_n10022.n3 a_n3493_n10022.n2 10.8376
R13918 a_n3493_n10022.n5 a_n3493_n10022.n3 2.50485
R13919 a_n126_n9484.t0 a_n126_n9484.t1 87.1434
R13920 a_6167_n9484.n1 a_6167_n9484.t3 530.01
R13921 a_6167_n9484.t1 a_6167_n9484.n5 421.021
R13922 a_6167_n9484.n0 a_6167_n9484.t7 337.142
R13923 a_6167_n9484.n3 a_6167_n9484.t0 280.223
R13924 a_6167_n9484.n4 a_6167_n9484.t6 263.173
R13925 a_6167_n9484.n4 a_6167_n9484.t2 227.826
R13926 a_6167_n9484.n0 a_6167_n9484.t4 199.762
R13927 a_6167_n9484.n2 a_6167_n9484.n1 170.81
R13928 a_6167_n9484.n2 a_6167_n9484.n0 167.321
R13929 a_6167_n9484.n5 a_6167_n9484.n4 152
R13930 a_6167_n9484.n1 a_6167_n9484.t5 141.923
R13931 a_6167_n9484.n3 a_6167_n9484.n2 10.8376
R13932 a_6167_n9484.n5 a_6167_n9484.n3 2.50485
R13933 a_958_n4702.n0 a_958_n4702.t1 68.3338
R13934 a_958_n4702.n0 a_958_n4702.t0 26.3935
R13935 a_958_n4702.n1 a_958_n4702.n0 14.4005
R13936 a_7422_n1029.t0 a_7422_n1029.t1 87.1434
R13937 a_1806_n9484.t0 a_1806_n9484.t1 87.1434
R13938 a_1627_n9510.n5 a_1627_n9510.n4 807.871
R13939 a_1627_n9510.n2 a_1627_n9510.t6 389.183
R13940 a_1627_n9510.n3 a_1627_n9510.n2 251.167
R13941 a_1627_n9510.n3 a_1627_n9510.t2 223.571
R13942 a_1627_n9510.n0 a_1627_n9510.t8 212.081
R13943 a_1627_n9510.n1 a_1627_n9510.t4 212.081
R13944 a_1627_n9510.n4 a_1627_n9510.n1 176.576
R13945 a_1627_n9510.n2 a_1627_n9510.t5 174.891
R13946 a_1627_n9510.n0 a_1627_n9510.t7 139.78
R13947 a_1627_n9510.n1 a_1627_n9510.t3 139.78
R13948 a_1627_n9510.n5 a_1627_n9510.t1 63.3219
R13949 a_1627_n9510.t0 a_1627_n9510.n5 63.3219
R13950 a_1627_n9510.n1 a_1627_n9510.n0 61.346
R13951 a_1627_n9510.n4 a_1627_n9510.n3 37.7195
R13952 a_6333_n10022.t1 a_6333_n10022.n3 370.026
R13953 a_6333_n10022.n0 a_6333_n10022.t2 351.356
R13954 a_6333_n10022.n1 a_6333_n10022.t4 334.717
R13955 a_6333_n10022.n3 a_6333_n10022.t0 325.971
R13956 a_6333_n10022.n1 a_6333_n10022.t3 309.935
R13957 a_6333_n10022.n0 a_6333_n10022.t5 305.683
R13958 a_6333_n10022.n2 a_6333_n10022.n0 16.879
R13959 a_6333_n10022.n3 a_6333_n10022.n2 10.8867
R13960 a_6333_n10022.n2 a_6333_n10022.n1 9.3005
R13961 a_6153_n1029.t1 a_6153_n1029.n3 370.026
R13962 a_6153_n1029.n0 a_6153_n1029.t3 351.356
R13963 a_6153_n1029.n1 a_6153_n1029.t4 334.717
R13964 a_6153_n1029.n3 a_6153_n1029.t0 325.971
R13965 a_6153_n1029.n1 a_6153_n1029.t5 309.935
R13966 a_6153_n1029.n0 a_6153_n1029.t2 305.683
R13967 a_6153_n1029.n2 a_6153_n1029.n0 16.879
R13968 a_6153_n1029.n3 a_6153_n1029.n2 10.8867
R13969 a_6153_n1029.n2 a_6153_n1029.n1 9.3005
R13970 a_7230_n663.t0 a_7230_n663.t1 126.644
R13971 a_792_n9662.n1 a_792_n9662.n0 926.024
R13972 a_792_n9662.t0 a_792_n9662.n1 82.0838
R13973 a_792_n9662.n0 a_792_n9662.t1 63.3338
R13974 a_792_n9662.n1 a_792_n9662.t3 63.3219
R13975 a_792_n9662.n0 a_792_n9662.t2 29.7268
R13976 a_n3072_n9484.n1 a_n3072_n9484.n0 926.024
R13977 a_n3072_n9484.n0 a_n3072_n9484.t3 82.0838
R13978 a_n3072_n9484.n1 a_n3072_n9484.t0 63.3338
R13979 a_n3072_n9484.n0 a_n3072_n9484.t2 63.3219
R13980 a_n3072_n9484.n2 a_n3072_n9484.t1 26.3935
R13981 a_n3072_n9484.n3 a_n3072_n9484.n2 14.4005
R13982 a_n3072_n9484.n2 a_n3072_n9484.n1 3.33383
R13983 a_1760_n5650.n5 a_1760_n5650.n4 807.871
R13984 a_1760_n5650.n0 a_1760_n5650.t4 389.183
R13985 a_1760_n5650.n1 a_1760_n5650.n0 251.167
R13986 a_1760_n5650.n1 a_1760_n5650.t2 223.571
R13987 a_1760_n5650.n3 a_1760_n5650.t3 212.081
R13988 a_1760_n5650.n2 a_1760_n5650.t8 212.081
R13989 a_1760_n5650.n4 a_1760_n5650.n3 176.576
R13990 a_1760_n5650.n0 a_1760_n5650.t6 174.891
R13991 a_1760_n5650.n3 a_1760_n5650.t7 139.78
R13992 a_1760_n5650.n2 a_1760_n5650.t5 139.78
R13993 a_1760_n5650.t0 a_1760_n5650.n5 63.3219
R13994 a_1760_n5650.n5 a_1760_n5650.t1 63.3219
R13995 a_1760_n5650.n3 a_1760_n5650.n2 61.346
R13996 a_1760_n5650.n4 a_1760_n5650.n1 37.5061
R13997 DOUT[2].n3 DOUT[2].n2 585
R13998 DOUT[2].n4 DOUT[2].n3 585
R13999 DOUT[2].n1 DOUT[2].n0 185
R14000 DOUT[2] DOUT[2].n1 49.0339
R14001 DOUT[2].n3 DOUT[2].t3 26.5955
R14002 DOUT[2].n3 DOUT[2].t2 26.5955
R14003 DOUT[2].n0 DOUT[2].t0 24.9236
R14004 DOUT[2].n0 DOUT[2].t1 24.9236
R14005 DOUT[2] DOUT[2].n4 20.4366
R14006 DOUT[2].n2 DOUT[2] 15.6165
R14007 DOUT[2].n1 DOUT[2] 10.4965
R14008 DOUT[2].n4 DOUT[2] 1.7925
R14009 DOUT[2].n2 DOUT[2] 1.7925
R14010 a_7951_3557.n1 a_7951_3557.t3 530.01
R14011 a_7951_3557.t1 a_7951_3557.n5 421.021
R14012 a_7951_3557.n0 a_7951_3557.t6 337.142
R14013 a_7951_3557.n3 a_7951_3557.t0 280.223
R14014 a_7951_3557.n4 a_7951_3557.t4 263.173
R14015 a_7951_3557.n4 a_7951_3557.t5 227.826
R14016 a_7951_3557.n0 a_7951_3557.t7 199.762
R14017 a_7951_3557.n2 a_7951_3557.n1 170.81
R14018 a_7951_3557.n2 a_7951_3557.n0 167.321
R14019 a_7951_3557.n5 a_7951_3557.n4 152
R14020 a_7951_3557.n1 a_7951_3557.t2 141.923
R14021 a_7951_3557.n3 a_7951_3557.n2 10.8376
R14022 a_7951_3557.n5 a_7951_3557.n3 2.50485
R14023 a_8372_3557.n1 a_8372_3557.n0 926.024
R14024 a_8372_3557.n0 a_8372_3557.t3 82.0838
R14025 a_8372_3557.n1 a_8372_3557.t0 63.3338
R14026 a_8372_3557.n0 a_8372_3557.t2 63.3219
R14027 a_8372_3557.n2 a_8372_3557.t1 26.3935
R14028 a_8372_3557.n3 a_8372_3557.n2 14.4005
R14029 a_8372_3557.n2 a_8372_3557.n1 3.33383
R14030 a_8467_3557.n3 a_8467_3557.n2 674.338
R14031 a_8467_3557.n1 a_8467_3557.t4 332.58
R14032 a_8467_3557.n2 a_8467_3557.n0 284.012
R14033 a_8467_3557.n2 a_8467_3557.n1 253.648
R14034 a_8467_3557.n1 a_8467_3557.t5 168.701
R14035 a_8467_3557.t1 a_8467_3557.n3 96.1553
R14036 a_8467_3557.n3 a_8467_3557.t2 65.6672
R14037 a_8467_3557.n0 a_8467_3557.t0 65.0005
R14038 a_8467_3557.n0 a_8467_3557.t3 45.0005
R14039 a_9194_3923.t0 a_9194_3923.t1 126.644
R14040 a_3181_n1207.t0 a_3181_n1207.t1 60.0005
R14041 a_3559_n9724.n4 a_3559_n9724.n1 807.871
R14042 a_3559_n9724.n0 a_3559_n9724.t6 389.183
R14043 a_3559_n9724.n5 a_3559_n9724.n0 251.167
R14044 a_3559_n9724.t0 a_3559_n9724.n5 223.571
R14045 a_3559_n9724.n2 a_3559_n9724.t8 212.081
R14046 a_3559_n9724.n3 a_3559_n9724.t4 212.081
R14047 a_3559_n9724.n4 a_3559_n9724.n3 176.576
R14048 a_3559_n9724.n0 a_3559_n9724.t5 174.891
R14049 a_3559_n9724.n2 a_3559_n9724.t7 139.78
R14050 a_3559_n9724.n3 a_3559_n9724.t3 139.78
R14051 a_3559_n9724.n1 a_3559_n9724.t1 63.3219
R14052 a_3559_n9724.n1 a_3559_n9724.t2 63.3219
R14053 a_3559_n9724.n3 a_3559_n9724.n2 61.346
R14054 a_3559_n9724.n5 a_3559_n9724.n4 37.7195
R14055 SWN[6].n4 SWN[6].n3 585
R14056 SWN[6].n3 SWN[6].n2 585
R14057 SWN[6].n1 SWN[6].n0 185
R14058 SWN[6].n5 SWN[6].n1 53.3859
R14059 SWN[6].n3 SWN[6].t2 26.5955
R14060 SWN[6].n3 SWN[6].t3 26.5955
R14061 SWN[6].n0 SWN[6].t0 24.9236
R14062 SWN[6].n0 SWN[6].t1 24.9236
R14063 SWN[6] SWN[6].n5 14.676
R14064 SWN[6] SWN[6].n4 10.4965
R14065 SWN[6].n2 SWN[6] 10.4965
R14066 SWN[6].n4 SWN[6] 6.9125
R14067 SWN[6].n2 SWN[6] 6.9125
R14068 SWN[6].n5 SWN[6] 4.3525
R14069 SWN[6].n1 SWN[6] 1.7925
R14070 a_2325_n5356.t1 a_2325_n5356.n3 370.026
R14071 a_2325_n5356.n0 a_2325_n5356.t2 351.356
R14072 a_2325_n5356.n1 a_2325_n5356.t4 334.717
R14073 a_2325_n5356.n3 a_2325_n5356.t0 325.971
R14074 a_2325_n5356.n1 a_2325_n5356.t3 309.935
R14075 a_2325_n5356.n0 a_2325_n5356.t5 305.683
R14076 a_2325_n5356.n2 a_2325_n5356.n0 16.879
R14077 a_2325_n5356.n3 a_2325_n5356.n2 10.8867
R14078 a_2325_n5356.n2 a_2325_n5356.n1 9.3005
R14079 a_2047_n5372.n3 a_2047_n5372.n2 636.953
R14080 a_2047_n5372.n1 a_2047_n5372.t5 366.856
R14081 a_2047_n5372.n2 a_2047_n5372.n0 300.2
R14082 a_2047_n5372.n2 a_2047_n5372.n1 225.036
R14083 a_2047_n5372.n1 a_2047_n5372.t4 174.056
R14084 a_2047_n5372.n0 a_2047_n5372.t0 70.0005
R14085 a_2047_n5372.n3 a_2047_n5372.t2 68.0124
R14086 a_2047_n5372.t1 a_2047_n5372.n3 63.3219
R14087 a_2047_n5372.n0 a_2047_n5372.t3 61.6672
R14088 a_2183_n1599.n4 a_2183_n1599.n1 807.871
R14089 a_2183_n1599.n0 a_2183_n1599.t7 389.183
R14090 a_2183_n1599.n5 a_2183_n1599.n0 251.167
R14091 a_2183_n1599.t0 a_2183_n1599.n5 223.571
R14092 a_2183_n1599.n3 a_2183_n1599.t6 212.081
R14093 a_2183_n1599.n2 a_2183_n1599.t4 212.081
R14094 a_2183_n1599.n4 a_2183_n1599.n3 176.576
R14095 a_2183_n1599.n0 a_2183_n1599.t5 174.891
R14096 a_2183_n1599.n3 a_2183_n1599.t3 139.78
R14097 a_2183_n1599.n2 a_2183_n1599.t8 139.78
R14098 a_2183_n1599.n1 a_2183_n1599.t2 63.3219
R14099 a_2183_n1599.n1 a_2183_n1599.t1 63.3219
R14100 a_2183_n1599.n3 a_2183_n1599.n2 61.346
R14101 a_2183_n1599.n5 a_2183_n1599.n4 37.5061
R14102 CF[1].n9 CF[1].n8 585
R14103 CF[1].n10 CF[1].n9 585
R14104 CF[1].n12 CF[1].t7 332.312
R14105 CF[1].n12 CF[1].t4 295.627
R14106 CF[1].n3 CF[1].t8 294.557
R14107 CF[1].n0 CF[1].t6 294.557
R14108 CF[1].n3 CF[1].t5 211.01
R14109 CF[1].n0 CF[1].t9 211.01
R14110 CF[1] CF[1].n12 196.004
R14111 CF[1].n7 CF[1].n6 185
R14112 CF[1].n4 CF[1].n3 153.097
R14113 CF[1].n1 CF[1].n0 152
R14114 CF[1] CF[1].n14 67.7696
R14115 CF[1] CF[1].n7 57.7379
R14116 CF[1].n13 CF[1] 37.1376
R14117 CF[1].n14 CF[1] 33.3154
R14118 CF[1].n9 CF[1].t2 26.5955
R14119 CF[1].n9 CF[1].t3 26.5955
R14120 CF[1].n6 CF[1].t1 24.9236
R14121 CF[1].n6 CF[1].t0 24.9236
R14122 CF[1].n5 CF[1].n2 14.9321
R14123 CF[1].n13 CF[1].n11 14.7279
R14124 CF[1].n5 CF[1].n4 13.9063
R14125 CF[1].n8 CF[1] 10.4965
R14126 CF[1].n10 CF[1] 10.4965
R14127 CF[1].n2 CF[1] 9.32621
R14128 CF[1].n14 CF[1] 8.568
R14129 CF[1].n8 CF[1] 6.9125
R14130 CF[1].n11 CF[1] 4.3525
R14131 CF[1].n4 CF[1] 3.10907
R14132 CF[1].n11 CF[1].n10 2.5605
R14133 CF[1].n1 CF[1] 2.01193
R14134 CF[1].n7 CF[1] 1.7925
R14135 CF[1].n2 CF[1].n1 1.09764
R14136 CF[1] CF[1].n13 0.885115
R14137 CF[1] CF[1].n5 0.830241
R14138 a_519_n5258.n3 a_519_n5258.n2 647.119
R14139 a_519_n5258.n1 a_519_n5258.t5 350.253
R14140 a_519_n5258.n2 a_519_n5258.n0 260.339
R14141 a_519_n5258.n2 a_519_n5258.n1 246.119
R14142 a_519_n5258.n1 a_519_n5258.t4 189.588
R14143 a_519_n5258.n3 a_519_n5258.t2 89.1195
R14144 a_519_n5258.n0 a_519_n5258.t1 63.3338
R14145 a_519_n5258.t3 a_519_n5258.n3 41.0422
R14146 a_519_n5258.n0 a_519_n5258.t0 31.9797
R14147 a_733_n5258.t0 a_733_n5258.n0 1327.82
R14148 a_733_n5258.n0 a_733_n5258.t1 194.655
R14149 a_733_n5258.n0 a_733_n5258.t2 63.3219
R14150 a_5985_n4714.n1 a_5985_n4714.n0 926.024
R14151 a_5985_n4714.t1 a_5985_n4714.n1 82.0838
R14152 a_5985_n4714.n0 a_5985_n4714.t0 63.3338
R14153 a_5985_n4714.n1 a_5985_n4714.t3 63.3219
R14154 a_5985_n4714.n0 a_5985_n4714.t2 29.7268
R14155 a_6080_n4702.n3 a_6080_n4702.n2 674.338
R14156 a_6080_n4702.n1 a_6080_n4702.t5 332.58
R14157 a_6080_n4702.n2 a_6080_n4702.n0 284.012
R14158 a_6080_n4702.n2 a_6080_n4702.n1 253.648
R14159 a_6080_n4702.n1 a_6080_n4702.t4 168.701
R14160 a_6080_n4702.t1 a_6080_n4702.n3 96.1553
R14161 a_6080_n4702.n3 a_6080_n4702.t2 65.6672
R14162 a_6080_n4702.n0 a_6080_n4702.t0 65.0005
R14163 a_6080_n4702.n0 a_6080_n4702.t3 45.0005
R14164 a_8265_n10022.t1 a_8265_n10022.n3 370.026
R14165 a_8265_n10022.n0 a_8265_n10022.t4 351.356
R14166 a_8265_n10022.n1 a_8265_n10022.t2 334.717
R14167 a_8265_n10022.n3 a_8265_n10022.t0 325.971
R14168 a_8265_n10022.n1 a_8265_n10022.t5 309.935
R14169 a_8265_n10022.n0 a_8265_n10022.t3 305.683
R14170 a_8265_n10022.n2 a_8265_n10022.n0 16.879
R14171 a_8265_n10022.n3 a_8265_n10022.n2 10.8867
R14172 a_8265_n10022.n2 a_8265_n10022.n1 9.3005
R14173 a_8711_n9650.t0 a_8711_n9650.t1 198.571
R14174 a_n5004_n9662.n1 a_n5004_n9662.n0 926.024
R14175 a_n5004_n9662.t1 a_n5004_n9662.n1 82.0838
R14176 a_n5004_n9662.n0 a_n5004_n9662.t0 63.3338
R14177 a_n5004_n9662.n1 a_n5004_n9662.t3 63.3219
R14178 a_n5004_n9662.n0 a_n5004_n9662.t2 29.7268
R14179 a_1105_n10054.n3 a_1105_n10054.n2 647.119
R14180 a_1105_n10054.n1 a_1105_n10054.t5 350.253
R14181 a_1105_n10054.n2 a_1105_n10054.n0 260.339
R14182 a_1105_n10054.n2 a_1105_n10054.n1 246.119
R14183 a_1105_n10054.n1 a_1105_n10054.t4 189.588
R14184 a_1105_n10054.n3 a_1105_n10054.t3 89.1195
R14185 a_1105_n10054.n0 a_1105_n10054.t2 63.3338
R14186 a_1105_n10054.t0 a_1105_n10054.n3 41.0422
R14187 a_1105_n10054.n0 a_1105_n10054.t1 31.9797
R14188 a_995_n10028.n0 a_995_n10028.t2 1327.82
R14189 a_995_n10028.n0 a_995_n10028.t1 194.655
R14190 a_995_n10028.t0 a_995_n10028.n0 63.3219
R14191 a_2303_n9484.n1 a_2303_n9484.t6 530.01
R14192 a_2303_n9484.t0 a_2303_n9484.n5 421.021
R14193 a_2303_n9484.n0 a_2303_n9484.t4 337.142
R14194 a_2303_n9484.n3 a_2303_n9484.t1 280.223
R14195 a_2303_n9484.n4 a_2303_n9484.t3 263.173
R14196 a_2303_n9484.n4 a_2303_n9484.t5 227.826
R14197 a_2303_n9484.n0 a_2303_n9484.t7 199.762
R14198 a_2303_n9484.n2 a_2303_n9484.n1 170.81
R14199 a_2303_n9484.n2 a_2303_n9484.n0 167.321
R14200 a_2303_n9484.n5 a_2303_n9484.n4 152
R14201 a_2303_n9484.n1 a_2303_n9484.t2 141.923
R14202 a_2303_n9484.n3 a_2303_n9484.n2 10.8376
R14203 a_2303_n9484.n5 a_2303_n9484.n3 2.50485
R14204 a_2724_n9484.n1 a_2724_n9484.n0 926.024
R14205 a_2724_n9484.n0 a_2724_n9484.t2 82.0838
R14206 a_2724_n9484.n1 a_2724_n9484.t3 63.3338
R14207 a_2724_n9484.n0 a_2724_n9484.t1 63.3219
R14208 a_2724_n9484.n2 a_2724_n9484.t0 26.3935
R14209 a_2724_n9484.n3 a_2724_n9484.n2 14.4005
R14210 a_2724_n9484.n2 a_2724_n9484.n1 3.33383
R14211 a_2819_n9484.n3 a_2819_n9484.n2 674.338
R14212 a_2819_n9484.n1 a_2819_n9484.t4 332.58
R14213 a_2819_n9484.n2 a_2819_n9484.n0 284.012
R14214 a_2819_n9484.n2 a_2819_n9484.n1 253.648
R14215 a_2819_n9484.n1 a_2819_n9484.t5 168.701
R14216 a_2819_n9484.n3 a_2819_n9484.t3 96.1553
R14217 a_2819_n9484.t1 a_2819_n9484.n3 65.6672
R14218 a_2819_n9484.n0 a_2819_n9484.t2 65.0005
R14219 a_2819_n9484.n0 a_2819_n9484.t0 45.0005
R14220 a_n4344_n9650.n3 a_n4344_n9650.n2 636.953
R14221 a_n4344_n9650.n1 a_n4344_n9650.t4 366.856
R14222 a_n4344_n9650.n2 a_n4344_n9650.n0 300.2
R14223 a_n4344_n9650.n2 a_n4344_n9650.n1 225.036
R14224 a_n4344_n9650.n1 a_n4344_n9650.t5 174.056
R14225 a_n4344_n9650.n0 a_n4344_n9650.t3 70.0005
R14226 a_n4344_n9650.t1 a_n4344_n9650.n3 68.0124
R14227 a_n4344_n9650.n3 a_n4344_n9650.t2 63.3219
R14228 a_n4344_n9650.n0 a_n4344_n9650.t0 61.6672
R14229 a_n3990_n9662.t0 a_n3990_n9662.t1 87.1434
R14230 a_390_n5624.n0 a_390_n5624.t1 68.3338
R14231 a_390_n5624.n0 a_390_n5624.t0 26.3935
R14232 a_390_n5624.n1 a_390_n5624.n0 14.4005
R14233 a_n5922_n9484.t0 a_n5922_n9484.t1 87.1434
R14234 a_6018_2717.n1 a_6018_2717.t5 530.01
R14235 a_6018_2717.t1 a_6018_2717.n5 421.021
R14236 a_6018_2717.n0 a_6018_2717.t3 337.142
R14237 a_6018_2717.n3 a_6018_2717.t0 280.223
R14238 a_6018_2717.n4 a_6018_2717.t7 263.173
R14239 a_6018_2717.n4 a_6018_2717.t6 227.826
R14240 a_6018_2717.n0 a_6018_2717.t2 199.762
R14241 a_6018_2717.n2 a_6018_2717.n1 170.81
R14242 a_6018_2717.n2 a_6018_2717.n0 167.321
R14243 a_6018_2717.n5 a_6018_2717.n4 152
R14244 a_6018_2717.n1 a_6018_2717.t4 141.923
R14245 a_6018_2717.n3 a_6018_2717.n2 10.8376
R14246 a_6018_2717.n5 a_6018_2717.n3 2.50485
R14247 a_7099_2717.n3 a_7099_2717.n2 636.953
R14248 a_7099_2717.n1 a_7099_2717.t4 366.856
R14249 a_7099_2717.n2 a_7099_2717.n0 300.2
R14250 a_7099_2717.n2 a_7099_2717.n1 225.036
R14251 a_7099_2717.n1 a_7099_2717.t5 174.056
R14252 a_7099_2717.n0 a_7099_2717.t1 70.0005
R14253 a_7099_2717.n3 a_7099_2717.t2 68.0124
R14254 a_7099_2717.t0 a_7099_2717.n3 63.3219
R14255 a_7099_2717.n0 a_7099_2717.t3 61.6672
R14256 a_7208_2717.t1 a_7208_2717.t0 94.7268
R14257 a_887_n9650.n3 a_887_n9650.n2 674.338
R14258 a_887_n9650.n1 a_887_n9650.t4 332.58
R14259 a_887_n9650.n2 a_887_n9650.n0 284.012
R14260 a_887_n9650.n2 a_887_n9650.n1 253.648
R14261 a_887_n9650.n1 a_887_n9650.t5 168.701
R14262 a_887_n9650.n3 a_887_n9650.t2 96.1553
R14263 a_887_n9650.t0 a_887_n9650.n3 65.6672
R14264 a_887_n9650.n0 a_887_n9650.t3 65.0005
R14265 a_887_n9650.n0 a_887_n9650.t1 45.0005
R14266 a_393_n5356.t0 a_393_n5356.n3 370.026
R14267 a_393_n5356.n0 a_393_n5356.t4 351.356
R14268 a_393_n5356.n1 a_393_n5356.t5 334.717
R14269 a_393_n5356.n3 a_393_n5356.t1 325.971
R14270 a_393_n5356.n1 a_393_n5356.t3 309.935
R14271 a_393_n5356.n0 a_393_n5356.t2 305.683
R14272 a_393_n5356.n2 a_393_n5356.n0 16.879
R14273 a_393_n5356.n3 a_393_n5356.n2 10.8867
R14274 a_393_n5356.n2 a_393_n5356.n1 9.3005
R14275 a_349_n5258.t0 a_349_n5258.t1 126.644
R14276 a_115_n5372.n3 a_115_n5372.n2 636.953
R14277 a_115_n5372.n1 a_115_n5372.t4 366.856
R14278 a_115_n5372.n2 a_115_n5372.n0 300.2
R14279 a_115_n5372.n2 a_115_n5372.n1 225.036
R14280 a_115_n5372.n1 a_115_n5372.t5 174.056
R14281 a_115_n5372.n0 a_115_n5372.t1 70.0005
R14282 a_115_n5372.n3 a_115_n5372.t2 68.0124
R14283 a_115_n5372.t0 a_115_n5372.n3 63.3219
R14284 a_115_n5372.n0 a_115_n5372.t3 61.6672
R14285 a_1149_n9662.t0 a_1149_n9662.t1 60.0005
R14286 a_6185_3557.t1 a_6185_3557.n3 370.026
R14287 a_6185_3557.n0 a_6185_3557.t5 351.356
R14288 a_6185_3557.n1 a_6185_3557.t3 334.717
R14289 a_6185_3557.n3 a_6185_3557.t0 325.971
R14290 a_6185_3557.n1 a_6185_3557.t4 309.935
R14291 a_6185_3557.n0 a_6185_3557.t2 305.683
R14292 a_6185_3557.n2 a_6185_3557.n0 16.879
R14293 a_6185_3557.n3 a_6185_3557.n2 10.8867
R14294 a_6185_3557.n2 a_6185_3557.n1 9.3005
R14295 a_7262_3923.t0 a_7262_3923.t1 126.644
R14296 a_150_n5624.t0 a_150_n5624.t1 87.1434
R14297 a_4865_3557.t0 a_4865_3557.t1 60.0005
R14298 a_3083_n5258.n1 a_3083_n5258.n0 926.024
R14299 a_3083_n5258.t0 a_3083_n5258.n1 82.0838
R14300 a_3083_n5258.n0 a_3083_n5258.t1 63.3338
R14301 a_3083_n5258.n1 a_3083_n5258.t3 63.3219
R14302 a_3083_n5258.n0 a_3083_n5258.t2 29.7268
R14303 a_6611_n663.n0 a_6611_n663.t2 1327.82
R14304 a_6611_n663.n0 a_6611_n663.t1 194.655
R14305 a_6611_n663.t0 a_6611_n663.n0 63.3219
R14306 DOUT[1].n3 DOUT[1].n2 585
R14307 DOUT[1].n4 DOUT[1].n3 585
R14308 DOUT[1].n1 DOUT[1].n0 185
R14309 DOUT[1] DOUT[1].n1 57.7379
R14310 DOUT[1].n3 DOUT[1].t2 26.5955
R14311 DOUT[1].n3 DOUT[1].t3 26.5955
R14312 DOUT[1].n0 DOUT[1].t1 24.9236
R14313 DOUT[1].n0 DOUT[1].t0 24.9236
R14314 DOUT[1] DOUT[1].n5 17.8877
R14315 DOUT[1].n2 DOUT[1] 10.4965
R14316 DOUT[1].n4 DOUT[1] 10.4965
R14317 DOUT[1].n2 DOUT[1] 6.9125
R14318 DOUT[1].n5 DOUT[1] 4.3525
R14319 DOUT[1].n5 DOUT[1].n4 2.5605
R14320 DOUT[1].n1 DOUT[1] 1.7925
R14321 a_n2303_n9650.n0 a_n2303_n9650.t1 68.3338
R14322 a_n2303_n9650.n0 a_n2303_n9650.t0 26.3935
R14323 a_n2303_n9650.n1 a_n2303_n9650.n0 14.4005
R14324 a_2123_n1029.n1 a_2123_n1029.t3 530.01
R14325 a_2123_n1029.t1 a_2123_n1029.n5 421.021
R14326 a_2123_n1029.n0 a_2123_n1029.t6 337.142
R14327 a_2123_n1029.n3 a_2123_n1029.t0 280.223
R14328 a_2123_n1029.n4 a_2123_n1029.t7 263.173
R14329 a_2123_n1029.n4 a_2123_n1029.t4 227.826
R14330 a_2123_n1029.n0 a_2123_n1029.t5 199.762
R14331 a_2123_n1029.n2 a_2123_n1029.n1 170.81
R14332 a_2123_n1029.n2 a_2123_n1029.n0 167.321
R14333 a_2123_n1029.n5 a_2123_n1029.n4 152
R14334 a_2123_n1029.n1 a_2123_n1029.t2 141.923
R14335 a_2123_n1029.n3 a_2123_n1029.n2 10.8376
R14336 a_2123_n1029.n5 a_2123_n1029.n3 2.50485
R14337 a_n2977_n9650.n3 a_n2977_n9650.n2 674.338
R14338 a_n2977_n9650.n1 a_n2977_n9650.t5 332.58
R14339 a_n2977_n9650.n2 a_n2977_n9650.n0 284.012
R14340 a_n2977_n9650.n2 a_n2977_n9650.n1 253.648
R14341 a_n2977_n9650.n1 a_n2977_n9650.t4 168.701
R14342 a_n2977_n9650.n3 a_n2977_n9650.t2 96.1553
R14343 a_n2977_n9650.t1 a_n2977_n9650.n3 65.6672
R14344 a_n2977_n9650.n0 a_n2977_n9650.t3 65.0005
R14345 a_n2977_n9650.n0 a_n2977_n9650.t0 45.0005
R14346 a_n8033_n9724.n5 a_n8033_n9724.n4 807.871
R14347 a_n8033_n9724.n2 a_n8033_n9724.t5 389.183
R14348 a_n8033_n9724.n3 a_n8033_n9724.n2 251.167
R14349 a_n8033_n9724.n3 a_n8033_n9724.t1 223.571
R14350 a_n8033_n9724.n0 a_n8033_n9724.t7 212.081
R14351 a_n8033_n9724.n1 a_n8033_n9724.t3 212.081
R14352 a_n8033_n9724.n4 a_n8033_n9724.n1 176.576
R14353 a_n8033_n9724.n2 a_n8033_n9724.t4 174.891
R14354 a_n8033_n9724.n0 a_n8033_n9724.t8 139.78
R14355 a_n8033_n9724.n1 a_n8033_n9724.t6 139.78
R14356 a_n8033_n9724.t0 a_n8033_n9724.n5 63.3219
R14357 a_n8033_n9724.n5 a_n8033_n9724.t2 63.3219
R14358 a_n8033_n9724.n1 a_n8033_n9724.n0 61.346
R14359 a_n8033_n9724.n4 a_n8033_n9724.n3 37.7195
R14360 SWN[0].n4 SWN[0].n3 585
R14361 SWN[0].n3 SWN[0].n2 585
R14362 SWN[0].n1 SWN[0].n0 185
R14363 SWN[0].n5 SWN[0].n1 53.3859
R14364 SWN[0].n3 SWN[0].t2 26.5955
R14365 SWN[0].n3 SWN[0].t3 26.5955
R14366 SWN[0].n0 SWN[0].t0 24.9236
R14367 SWN[0].n0 SWN[0].t1 24.9236
R14368 SWN[0] SWN[0].n5 14.6437
R14369 SWN[0] SWN[0].n4 10.4965
R14370 SWN[0].n2 SWN[0] 10.4965
R14371 SWN[0].n4 SWN[0] 6.9125
R14372 SWN[0].n2 SWN[0] 6.9125
R14373 SWN[0].n5 SWN[0] 4.3525
R14374 SWN[0].n1 SWN[0] 1.7925
R14375 a_5020_n1573.n0 a_5020_n1573.t1 1327.82
R14376 a_5020_n1573.t0 a_5020_n1573.n0 194.655
R14377 a_5020_n1573.n0 a_5020_n1573.t2 63.3219
R14378 a_4875_n1599.n3 a_4875_n1599.n2 674.338
R14379 a_4875_n1599.n1 a_4875_n1599.t4 332.58
R14380 a_4875_n1599.n2 a_4875_n1599.n0 284.012
R14381 a_4875_n1599.n2 a_4875_n1599.n1 253.648
R14382 a_4875_n1599.n1 a_4875_n1599.t5 168.701
R14383 a_4875_n1599.t0 a_4875_n1599.n3 96.1553
R14384 a_4875_n1599.n3 a_4875_n1599.t3 65.6672
R14385 a_4875_n1599.n0 a_4875_n1599.t1 65.0005
R14386 a_4875_n1599.n0 a_4875_n1599.t2 45.0005
R14387 CF[6].n11 CF[6].n10 585
R14388 CF[6].n12 CF[6].n11 585
R14389 CF[6].n6 CF[6].t8 333.651
R14390 CF[6].n6 CF[6].t6 297.233
R14391 CF[6].n3 CF[6].t9 294.557
R14392 CF[6].n0 CF[6].t4 294.557
R14393 CF[6].n3 CF[6].t7 211.01
R14394 CF[6].n0 CF[6].t5 211.01
R14395 CF[6].n7 CF[6].n6 196.493
R14396 CF[6].n9 CF[6].n8 185
R14397 CF[6].n4 CF[6].n3 153.097
R14398 CF[6].n1 CF[6].n0 152
R14399 CF[6] CF[6].n14 49.5617
R14400 CF[6] CF[6].n9 49.0339
R14401 CF[6].n13 CF[6].n7 35.37
R14402 CF[6].n11 CF[6].t2 26.5955
R14403 CF[6].n11 CF[6].t3 26.5955
R14404 CF[6].n8 CF[6].t0 24.9236
R14405 CF[6].n8 CF[6].t1 24.9236
R14406 CF[6].n14 CF[6] 19.7736
R14407 CF[6].n13 CF[6].n12 17.2879
R14408 CF[6].n10 CF[6] 15.6165
R14409 CF[6].n5 CF[6].n2 14.9321
R14410 CF[6].n5 CF[6].n4 13.9063
R14411 CF[6].n9 CF[6] 10.4965
R14412 CF[6].n2 CF[6] 9.32621
R14413 CF[6].n14 CF[6] 5.928
R14414 CF[6].n4 CF[6] 3.10907
R14415 CF[6].n1 CF[6] 2.01193
R14416 CF[6].n12 CF[6] 1.7925
R14417 CF[6].n10 CF[6] 1.7925
R14418 CF[6].n2 CF[6].n1 1.09764
R14419 CF[6] CF[6].n5 0.834552
R14420 CF[6] CF[6].n13 0.712038
R14421 CF[6].n7 CF[6] 0.24431
R14422 a_6184_2717.t1 a_6184_2717.n3 370.026
R14423 a_6184_2717.n0 a_6184_2717.t4 351.356
R14424 a_6184_2717.n1 a_6184_2717.t2 334.717
R14425 a_6184_2717.n3 a_6184_2717.t0 325.971
R14426 a_6184_2717.n1 a_6184_2717.t5 309.935
R14427 a_6184_2717.n0 a_6184_2717.t3 305.683
R14428 a_6184_2717.n2 a_6184_2717.n0 16.879
R14429 a_6184_2717.n3 a_6184_2717.n2 10.8867
R14430 a_6184_2717.n2 a_6184_2717.n1 9.3005
R14431 a_6534_2717.n3 a_6534_2717.n2 674.338
R14432 a_6534_2717.n1 a_6534_2717.t4 332.58
R14433 a_6534_2717.n2 a_6534_2717.n0 284.012
R14434 a_6534_2717.n2 a_6534_2717.n1 253.648
R14435 a_6534_2717.n1 a_6534_2717.t5 168.701
R14436 a_6534_2717.t1 a_6534_2717.n3 96.1553
R14437 a_6534_2717.n3 a_6534_2717.t3 65.6672
R14438 a_6534_2717.n0 a_6534_2717.t0 65.0005
R14439 a_6534_2717.n0 a_6534_2717.t2 45.0005
R14440 a_6630_2717.t0 a_6630_2717.t1 198.571
R14441 a_n1561_n9484.n1 a_n1561_n9484.t6 530.01
R14442 a_n1561_n9484.t1 a_n1561_n9484.n5 421.021
R14443 a_n1561_n9484.n0 a_n1561_n9484.t7 337.142
R14444 a_n1561_n9484.n3 a_n1561_n9484.t0 280.223
R14445 a_n1561_n9484.n4 a_n1561_n9484.t3 263.173
R14446 a_n1561_n9484.n4 a_n1561_n9484.t4 227.826
R14447 a_n1561_n9484.n0 a_n1561_n9484.t2 199.762
R14448 a_n1561_n9484.n2 a_n1561_n9484.n1 170.81
R14449 a_n1561_n9484.n2 a_n1561_n9484.n0 167.321
R14450 a_n1561_n9484.n5 a_n1561_n9484.n4 152
R14451 a_n1561_n9484.n1 a_n1561_n9484.t5 141.923
R14452 a_n1561_n9484.n3 a_n1561_n9484.n2 10.8376
R14453 a_n1561_n9484.n5 a_n1561_n9484.n3 2.50485
R14454 a_7453_2717.t0 a_7453_2717.t1 87.1434
R14455 a_2874_n1573.n3 a_2874_n1573.n2 647.119
R14456 a_2874_n1573.n1 a_2874_n1573.t5 350.253
R14457 a_2874_n1573.n2 a_2874_n1573.n0 260.339
R14458 a_2874_n1573.n2 a_2874_n1573.n1 246.119
R14459 a_2874_n1573.n1 a_2874_n1573.t4 189.588
R14460 a_2874_n1573.n3 a_2874_n1573.t2 89.1195
R14461 a_2874_n1573.n0 a_2874_n1573.t3 63.3338
R14462 a_2874_n1573.t1 a_2874_n1573.n3 41.0422
R14463 a_2874_n1573.n0 a_2874_n1573.t0 31.9797
R14464 a_2469_n9484.t1 a_2469_n9484.n3 370.026
R14465 a_2469_n9484.n0 a_2469_n9484.t5 351.356
R14466 a_2469_n9484.n1 a_2469_n9484.t3 334.717
R14467 a_2469_n9484.n3 a_2469_n9484.t0 325.971
R14468 a_2469_n9484.n1 a_2469_n9484.t4 309.935
R14469 a_2469_n9484.n0 a_2469_n9484.t2 305.683
R14470 a_2469_n9484.n2 a_2469_n9484.n0 16.879
R14471 a_2469_n9484.n3 a_2469_n9484.n2 10.8867
R14472 a_2469_n9484.n2 a_2469_n9484.n1 9.3005
R14473 a_3384_n9484.n3 a_3384_n9484.n2 636.953
R14474 a_3384_n9484.n1 a_3384_n9484.t5 366.856
R14475 a_3384_n9484.n2 a_3384_n9484.n0 300.2
R14476 a_3384_n9484.n2 a_3384_n9484.n1 225.036
R14477 a_3384_n9484.n1 a_3384_n9484.t4 174.056
R14478 a_3384_n9484.n0 a_3384_n9484.t1 70.0005
R14479 a_3384_n9484.n3 a_3384_n9484.t3 68.0124
R14480 a_3384_n9484.t0 a_3384_n9484.n3 63.3219
R14481 a_3384_n9484.n0 a_3384_n9484.t2 61.6672
R14482 a_3738_n9662.t0 a_3738_n9662.t1 87.1434
R14483 COMP_N.n6 COMP_N.t4 235.763
R14484 COMP_N.n1 COMP_N.t5 221.72
R14485 COMP_N.n0 COMP_N.t0 221.72
R14486 COMP_N.n6 COMP_N.t2 163.464
R14487 COMP_N.n3 COMP_N.n2 152
R14488 COMP_N.n5 COMP_N.n4 152
R14489 COMP_N.n7 COMP_N.n6 152
R14490 COMP_N.n1 COMP_N.t1 149.421
R14491 COMP_N.n0 COMP_N.t3 149.421
R14492 COMP_N.n2 COMP_N.n1 58.019
R14493 COMP_N.n5 COMP_N.n0 43.7375
R14494 COMP_N.n4 COMP_N.n3 21.7605
R14495 COMP_N.n7 COMP_N 19.5205
R14496 COMP_N.n6 COMP_N.n5 17.8524
R14497 COMP_N.n2 COMP_N.n0 16.9598
R14498 COMP_N COMP_N.n8 10.7837
R14499 COMP_N.n3 COMP_N 5.4405
R14500 COMP_N.n8 COMP_N 5.4405
R14501 COMP_N.n8 COMP_N.n7 4.4805
R14502 COMP_N.n4 COMP_N 2.2405
R14503 a_9289_n9484.t1 a_9289_n9484.t0 94.7268
R14504 a_3037_n10054.n3 a_3037_n10054.n2 647.119
R14505 a_3037_n10054.n1 a_3037_n10054.t4 350.253
R14506 a_3037_n10054.n2 a_3037_n10054.n0 260.339
R14507 a_3037_n10054.n2 a_3037_n10054.n1 246.119
R14508 a_3037_n10054.n1 a_3037_n10054.t5 189.588
R14509 a_3037_n10054.n3 a_3037_n10054.t2 89.1195
R14510 a_3037_n10054.n0 a_3037_n10054.t3 63.3338
R14511 a_3037_n10054.t0 a_3037_n10054.n3 41.0422
R14512 a_3037_n10054.n0 a_3037_n10054.t1 31.9797
R14513 a_2915_n9650.t0 a_2915_n9650.t1 198.571
R14514 a_3081_n9662.t0 a_3081_n9662.t1 60.0005
R14515 a_357_n1029.t1 a_357_n1029.n3 370.026
R14516 a_357_n1029.n0 a_357_n1029.t5 351.356
R14517 a_357_n1029.n1 a_357_n1029.t4 334.717
R14518 a_357_n1029.n3 a_357_n1029.t0 325.971
R14519 a_357_n1029.n1 a_357_n1029.t3 309.935
R14520 a_357_n1029.n0 a_357_n1029.t2 305.683
R14521 a_357_n1029.n2 a_357_n1029.n0 16.879
R14522 a_357_n1029.n3 a_357_n1029.n2 10.8867
R14523 a_357_n1029.n2 a_357_n1029.n1 9.3005
R14524 a_1434_n663.t0 a_1434_n663.t1 126.644
R14525 a_2322_n5624.n0 a_2322_n5624.t1 68.3338
R14526 a_2322_n5624.n0 a_2322_n5624.t0 26.3935
R14527 a_2322_n5624.n1 a_2322_n5624.n0 14.4005
R14528 a_6643_3923.t0 a_6643_3923.n0 1327.82
R14529 a_6643_3923.n0 a_6643_3923.t2 194.655
R14530 a_6643_3923.n0 a_6643_3923.t1 63.3219
R14531 a_n976_2959.n3 a_n976_2959.n2 647.119
R14532 a_n976_2959.n1 a_n976_2959.t4 350.253
R14533 a_n976_2959.n2 a_n976_2959.n0 260.339
R14534 a_n976_2959.n2 a_n976_2959.n1 246.119
R14535 a_n976_2959.n1 a_n976_2959.t5 189.588
R14536 a_n976_2959.n3 a_n976_2959.t3 89.1195
R14537 a_n976_2959.n0 a_n976_2959.t0 63.3338
R14538 a_n976_2959.t2 a_n976_2959.n3 41.0422
R14539 a_n976_2959.n0 a_n976_2959.t1 31.9797
R14540 a_n1098_2717.t1 a_n1098_2717.t0 198.571
R14541 a_n932_2717.t0 a_n932_2717.t1 60.0005
R14542 a_3253_n1207.t0 a_3253_n1207.t1 198.571
R14543 a_n520_2717.t0 a_n520_2717.t1 94.7268
R14544 CF[2].n9 CF[2].n8 585
R14545 CF[2].n10 CF[2].n9 585
R14546 CF[2].n12 CF[2].t6 332.312
R14547 CF[2].n12 CF[2].t8 295.627
R14548 CF[2].n3 CF[2].t5 294.557
R14549 CF[2].n0 CF[2].t7 294.557
R14550 CF[2].n3 CF[2].t4 211.01
R14551 CF[2].n0 CF[2].t9 211.01
R14552 CF[2] CF[2].n12 196.004
R14553 CF[2].n7 CF[2].n6 185
R14554 CF[2].n4 CF[2].n3 153.097
R14555 CF[2].n1 CF[2].n0 152
R14556 CF[2] CF[2].n14 63.7558
R14557 CF[2] CF[2].n7 57.7379
R14558 CF[2].n13 CF[2] 37.1376
R14559 CF[2].n14 CF[2] 28.8178
R14560 CF[2].n9 CF[2].t3 26.5955
R14561 CF[2].n9 CF[2].t2 26.5955
R14562 CF[2].n6 CF[2].t1 24.9236
R14563 CF[2].n6 CF[2].t0 24.9236
R14564 CF[2].n5 CF[2].n2 14.9321
R14565 CF[2].n13 CF[2].n11 14.7279
R14566 CF[2].n5 CF[2].n4 13.9063
R14567 CF[2].n8 CF[2] 10.4965
R14568 CF[2].n10 CF[2] 10.4965
R14569 CF[2].n2 CF[2] 9.32621
R14570 CF[2].n14 CF[2] 8.41175
R14571 CF[2].n8 CF[2] 6.9125
R14572 CF[2].n11 CF[2] 4.3525
R14573 CF[2].n4 CF[2] 3.10907
R14574 CF[2].n11 CF[2].n10 2.5605
R14575 CF[2].n1 CF[2] 2.01193
R14576 CF[2].n7 CF[2] 1.7925
R14577 CF[2].n2 CF[2].n1 1.09764
R14578 CF[2] CF[2].n13 0.909154
R14579 CF[2] CF[2].n5 0.834552
R14580 a_3135_n4714.t0 a_3135_n4714.t1 87.1434
R14581 a_4086_2717.n1 a_4086_2717.t4 530.01
R14582 a_4086_2717.t1 a_4086_2717.n5 421.021
R14583 a_4086_2717.n0 a_4086_2717.t6 337.142
R14584 a_4086_2717.n3 a_4086_2717.t0 280.223
R14585 a_4086_2717.n4 a_4086_2717.t3 263.173
R14586 a_4086_2717.n4 a_4086_2717.t2 227.826
R14587 a_4086_2717.n0 a_4086_2717.t5 199.762
R14588 a_4086_2717.n2 a_4086_2717.n1 170.81
R14589 a_4086_2717.n2 a_4086_2717.n0 167.321
R14590 a_4086_2717.n5 a_4086_2717.n4 152
R14591 a_4086_2717.n1 a_4086_2717.t7 141.923
R14592 a_4086_2717.n3 a_4086_2717.n2 10.8376
R14593 a_4086_2717.n5 a_4086_2717.n3 2.50485
R14594 a_4252_2717.t1 a_4252_2717.n3 370.026
R14595 a_4252_2717.n0 a_4252_2717.t5 351.356
R14596 a_4252_2717.n1 a_4252_2717.t3 334.717
R14597 a_4252_2717.n3 a_4252_2717.t0 325.971
R14598 a_4252_2717.n1 a_4252_2717.t2 309.935
R14599 a_4252_2717.n0 a_4252_2717.t4 305.683
R14600 a_4252_2717.n2 a_4252_2717.n0 16.879
R14601 a_4252_2717.n3 a_4252_2717.n2 10.8867
R14602 a_4252_2717.n2 a_4252_2717.n1 9.3005
R14603 a_4476_n1029.n1 a_4476_n1029.n0 926.024
R14604 a_4476_n1029.t0 a_4476_n1029.n1 82.0838
R14605 a_4476_n1029.n0 a_4476_n1029.t3 63.3338
R14606 a_4476_n1029.n1 a_4476_n1029.t2 63.3219
R14607 a_4476_n1029.n0 a_4476_n1029.t1 29.7268
R14608 a_n7854_n9662.t0 a_n7854_n9662.t1 87.1434
R14609 a_8247_n5258.n3 a_8247_n5258.n2 647.119
R14610 a_8247_n5258.n1 a_8247_n5258.t4 350.253
R14611 a_8247_n5258.n2 a_8247_n5258.n0 260.339
R14612 a_8247_n5258.n2 a_8247_n5258.n1 246.119
R14613 a_8247_n5258.n1 a_8247_n5258.t5 189.588
R14614 a_8247_n5258.n3 a_8247_n5258.t3 89.1195
R14615 a_8247_n5258.n0 a_8247_n5258.t2 63.3338
R14616 a_8247_n5258.t0 a_8247_n5258.n3 41.0422
R14617 a_8247_n5258.n0 a_8247_n5258.t1 31.9797
R14618 a_8554_n5624.t0 a_8554_n5624.t1 60.0005
R14619 a_8626_n5624.t0 a_8626_n5624.t1 198.571
R14620 a_9000_n1029.n3 a_9000_n1029.n2 636.953
R14621 a_9000_n1029.n1 a_9000_n1029.t4 366.856
R14622 a_9000_n1029.n2 a_9000_n1029.n0 300.2
R14623 a_9000_n1029.n2 a_9000_n1029.n1 225.036
R14624 a_9000_n1029.n1 a_9000_n1029.t5 174.056
R14625 a_9000_n1029.n0 a_9000_n1029.t2 70.0005
R14626 a_9000_n1029.t0 a_9000_n1029.n3 68.0124
R14627 a_9000_n1029.n3 a_9000_n1029.t1 63.3219
R14628 a_9000_n1029.n0 a_9000_n1029.t3 61.6672
R14629 a_9354_n1029.t0 a_9354_n1029.t1 87.1434
R14630 a_389_3557.t0 a_389_3557.n3 370.026
R14631 a_389_3557.n0 a_389_3557.t4 351.356
R14632 a_389_3557.n1 a_389_3557.t3 334.717
R14633 a_389_3557.n3 a_389_3557.t1 325.971
R14634 a_389_3557.n1 a_389_3557.t5 309.935
R14635 a_389_3557.n0 a_389_3557.t2 305.683
R14636 a_389_3557.n2 a_389_3557.n0 16.879
R14637 a_389_3557.n3 a_389_3557.n2 10.8867
R14638 a_389_3557.n2 a_389_3557.n1 9.3005
R14639 a_1466_3923.t0 a_1466_3923.t1 126.644
R14640 a_n3493_n9484.n1 a_n3493_n9484.t3 530.01
R14641 a_n3493_n9484.t1 a_n3493_n9484.n5 421.021
R14642 a_n3493_n9484.n0 a_n3493_n9484.t4 337.142
R14643 a_n3493_n9484.n3 a_n3493_n9484.t0 280.223
R14644 a_n3493_n9484.n4 a_n3493_n9484.t7 263.173
R14645 a_n3493_n9484.n4 a_n3493_n9484.t2 227.826
R14646 a_n3493_n9484.n0 a_n3493_n9484.t6 199.762
R14647 a_n3493_n9484.n2 a_n3493_n9484.n1 170.81
R14648 a_n3493_n9484.n2 a_n3493_n9484.n0 167.321
R14649 a_n3493_n9484.n5 a_n3493_n9484.n4 152
R14650 a_n3493_n9484.n1 a_n3493_n9484.t5 141.923
R14651 a_n3493_n9484.n3 a_n3493_n9484.n2 10.8376
R14652 a_n3493_n9484.n5 a_n3493_n9484.n3 2.50485
R14653 auto_sampling_0.x23.A.n3 auto_sampling_0.x23.A.t7 212.081
R14654 auto_sampling_0.x23.A.n5 auto_sampling_0.x23.A.t9 212.081
R14655 auto_sampling_0.x23.A.n2 auto_sampling_0.x23.A.t4 212.081
R14656 auto_sampling_0.x23.A.n10 auto_sampling_0.x23.A.t11 212.081
R14657 auto_sampling_0.x23.A.n15 auto_sampling_0.x23.A.n14 208.965
R14658 auto_sampling_0.x23.A.n11 auto_sampling_0.x23.A.n10 188.516
R14659 auto_sampling_0.x23.A.n4 auto_sampling_0.x23.A 154.304
R14660 auto_sampling_0.x23.A.n9 auto_sampling_0.x23.A.n8 152
R14661 auto_sampling_0.x23.A.n7 auto_sampling_0.x23.A.n6 152
R14662 auto_sampling_0.x23.A.n3 auto_sampling_0.x23.A.t10 139.78
R14663 auto_sampling_0.x23.A.n5 auto_sampling_0.x23.A.t5 139.78
R14664 auto_sampling_0.x23.A.n2 auto_sampling_0.x23.A.t8 139.78
R14665 auto_sampling_0.x23.A.n10 auto_sampling_0.x23.A.t6 139.78
R14666 auto_sampling_0.x23.A auto_sampling_0.x23.A.n0 96.8352
R14667 auto_sampling_0.x23.A.n4 auto_sampling_0.x23.A.n3 30.6732
R14668 auto_sampling_0.x23.A.n5 auto_sampling_0.x23.A.n4 30.6732
R14669 auto_sampling_0.x23.A.n6 auto_sampling_0.x23.A.n5 30.6732
R14670 auto_sampling_0.x23.A.n6 auto_sampling_0.x23.A.n2 30.6732
R14671 auto_sampling_0.x23.A.n9 auto_sampling_0.x23.A.n2 30.6732
R14672 auto_sampling_0.x23.A.n10 auto_sampling_0.x23.A.n9 30.6732
R14673 auto_sampling_0.x23.A.n14 auto_sampling_0.x23.A.t3 26.5955
R14674 auto_sampling_0.x23.A.n14 auto_sampling_0.x23.A.t2 26.5955
R14675 auto_sampling_0.x23.A.n0 auto_sampling_0.x23.A.t0 24.9236
R14676 auto_sampling_0.x23.A.n0 auto_sampling_0.x23.A.t1 24.9236
R14677 auto_sampling_0.x23.A.n7 auto_sampling_0.x23.A 19.2005
R14678 auto_sampling_0.x23.A.n13 auto_sampling_0.x23.A.n12 19.1625
R14679 auto_sampling_0.x23.A.n8 auto_sampling_0.x23.A 17.1525
R14680 auto_sampling_0.x23.A.n11 auto_sampling_0.x23.A 17.1525
R14681 auto_sampling_0.x23.A auto_sampling_0.x23.A.n13 13.0565
R14682 auto_sampling_0.x23.A auto_sampling_0.x23.A.n1 11.2645
R14683 auto_sampling_0.x23.A.n8 auto_sampling_0.x23.A 6.4005
R14684 auto_sampling_0.x23.A.n1 auto_sampling_0.x23.A 6.1445
R14685 auto_sampling_0.x23.A.n1 auto_sampling_0.x23.A 4.65505
R14686 auto_sampling_0.x23.A auto_sampling_0.x23.A.n7 4.3525
R14687 auto_sampling_0.x23.A.n12 auto_sampling_0.x23.A 4.3525
R14688 auto_sampling_0.x23.A.n13 auto_sampling_0.x23.A 4.3525
R14689 auto_sampling_0.x23.A.n12 auto_sampling_0.x23.A.n11 2.0485
R14690 auto_sampling_0.x23.A.n15 auto_sampling_0.x23.A 2.0485
R14691 auto_sampling_0.x23.A auto_sampling_0.x23.A.n15 1.55202
R14692 SWP[5].n0 SWP[5].t4 333.651
R14693 SWP[5].n0 SWP[5].t5 297.233
R14694 SWP[5].n4 SWP[5].n3 289.096
R14695 SWP[5].n1 SWP[5].n0 196.493
R14696 SWP[5].n6 SWP[5].n5 185
R14697 SWP[5] SWP[5].n6 49.0339
R14698 SWP[5].n2 SWP[5] 42.7158
R14699 SWP[5] SWP[5].n1 39.5065
R14700 SWP[5].n3 SWP[5].t2 26.5955
R14701 SWP[5].n3 SWP[5].t3 26.5955
R14702 SWP[5].n5 SWP[5].t0 24.9236
R14703 SWP[5].n5 SWP[5].t1 24.9236
R14704 SWP[5] SWP[5].n7 14.6178
R14705 SWP[5].n7 SWP[5] 13.0565
R14706 SWP[5].n2 SWP[5] 12.6429
R14707 SWP[5].n6 SWP[5] 10.4965
R14708 SWP[5] SWP[5].n2 9.5329
R14709 SWP[5] SWP[5].n4 9.48653
R14710 SWP[5].n4 SWP[5] 7.7181
R14711 SWP[5].n7 SWP[5] 4.3525
R14712 SWP[5].n1 SWP[5] 0.24431
R14713 a_8117_3557.t1 a_8117_3557.n3 370.026
R14714 a_8117_3557.n0 a_8117_3557.t2 351.356
R14715 a_8117_3557.n1 a_8117_3557.t5 334.717
R14716 a_8117_3557.n3 a_8117_3557.t0 325.971
R14717 a_8117_3557.n1 a_8117_3557.t3 309.935
R14718 a_8117_3557.n0 a_8117_3557.t4 305.683
R14719 a_8117_3557.n2 a_8117_3557.n0 16.879
R14720 a_8117_3557.n3 a_8117_3557.n2 10.8867
R14721 a_8117_3557.n2 a_8117_3557.n1 9.3005
R14722 a_8685_3799.n3 a_8685_3799.n2 647.119
R14723 a_8685_3799.n1 a_8685_3799.t4 350.253
R14724 a_8685_3799.n2 a_8685_3799.n0 260.339
R14725 a_8685_3799.n2 a_8685_3799.n1 246.119
R14726 a_8685_3799.n1 a_8685_3799.t5 189.588
R14727 a_8685_3799.n3 a_8685_3799.t0 89.1195
R14728 a_8685_3799.n0 a_8685_3799.t1 63.3338
R14729 a_8685_3799.t3 a_8685_3799.n3 41.0422
R14730 a_8685_3799.n0 a_8685_3799.t2 31.9797
R14731 a_9032_3557.n3 a_9032_3557.n2 636.953
R14732 a_9032_3557.n1 a_9032_3557.t5 366.856
R14733 a_9032_3557.n2 a_9032_3557.n0 300.2
R14734 a_9032_3557.n2 a_9032_3557.n1 225.036
R14735 a_9032_3557.n1 a_9032_3557.t4 174.056
R14736 a_9032_3557.n0 a_9032_3557.t2 70.0005
R14737 a_9032_3557.t0 a_9032_3557.n3 68.0124
R14738 a_9032_3557.n3 a_9032_3557.t3 63.3219
R14739 a_9032_3557.n0 a_9032_3557.t1 61.6672
R14740 a_8500_n1573.t0 a_8500_n1573.t1 126.644
R14741 a_8266_n1441.n3 a_8266_n1441.n2 636.953
R14742 a_8266_n1441.n1 a_8266_n1441.t4 366.856
R14743 a_8266_n1441.n2 a_8266_n1441.n0 300.2
R14744 a_8266_n1441.n2 a_8266_n1441.n1 225.036
R14745 a_8266_n1441.n1 a_8266_n1441.t5 174.056
R14746 a_8266_n1441.n0 a_8266_n1441.t2 70.0005
R14747 a_8266_n1441.t0 a_8266_n1441.n3 68.0124
R14748 a_8266_n1441.n3 a_8266_n1441.t3 63.3219
R14749 a_8266_n1441.n0 a_8266_n1441.t1 61.6672
R14750 a_6791_n9118.n0 a_6791_n9118.t2 1327.82
R14751 a_6791_n9118.n0 a_6791_n9118.t1 194.655
R14752 a_6791_n9118.t0 a_6791_n9118.n0 63.3219
R14753 a_8723_n9118.n0 a_8723_n9118.t2 1327.82
R14754 a_8723_n9118.t0 a_8723_n9118.n0 194.655
R14755 a_8723_n9118.n0 a_8723_n9118.t1 63.3219
R14756 a_4257_n5356.t0 a_4257_n5356.n3 370.026
R14757 a_4257_n5356.n0 a_4257_n5356.t2 351.356
R14758 a_4257_n5356.n1 a_4257_n5356.t3 334.717
R14759 a_4257_n5356.n3 a_4257_n5356.t1 325.971
R14760 a_4257_n5356.n1 a_4257_n5356.t5 309.935
R14761 a_4257_n5356.n0 a_4257_n5356.t4 305.683
R14762 a_4257_n5356.n2 a_4257_n5356.n0 16.879
R14763 a_4257_n5356.n3 a_4257_n5356.n2 10.8867
R14764 a_4257_n5356.n2 a_4257_n5356.n1 9.3005
R14765 a_3979_n5372.n3 a_3979_n5372.n2 636.953
R14766 a_3979_n5372.n1 a_3979_n5372.t4 366.856
R14767 a_3979_n5372.n2 a_3979_n5372.n0 300.2
R14768 a_3979_n5372.n2 a_3979_n5372.n1 225.036
R14769 a_3979_n5372.n1 a_3979_n5372.t5 174.056
R14770 a_3979_n5372.n0 a_3979_n5372.t2 70.0005
R14771 a_3979_n5372.n3 a_3979_n5372.t3 68.0124
R14772 a_3979_n5372.t1 a_3979_n5372.n3 63.3219
R14773 a_3979_n5372.n0 a_3979_n5372.t0 61.6672
R14774 a_388_2717.t1 a_388_2717.n3 370.026
R14775 a_388_2717.n0 a_388_2717.t5 351.356
R14776 a_388_2717.n1 a_388_2717.t4 334.717
R14777 a_388_2717.n3 a_388_2717.t0 325.971
R14778 a_388_2717.n1 a_388_2717.t2 309.935
R14779 a_388_2717.n0 a_388_2717.t3 305.683
R14780 a_388_2717.n2 a_388_2717.n0 16.879
R14781 a_388_2717.n3 a_388_2717.n2 10.8867
R14782 a_388_2717.n2 a_388_2717.n1 9.3005
R14783 a_643_2717.n1 a_643_2717.n0 926.024
R14784 a_643_2717.n0 a_643_2717.t3 82.0838
R14785 a_643_2717.n1 a_643_2717.t2 63.3338
R14786 a_643_2717.n0 a_643_2717.t1 63.3219
R14787 a_643_2717.n2 a_643_2717.t0 26.3935
R14788 a_643_2717.n3 a_643_2717.n2 14.4005
R14789 a_643_2717.n2 a_643_2717.n1 3.33383
R14790 a_738_2717.n3 a_738_2717.n2 674.338
R14791 a_738_2717.n1 a_738_2717.t4 332.58
R14792 a_738_2717.n2 a_738_2717.n0 284.012
R14793 a_738_2717.n2 a_738_2717.n1 253.648
R14794 a_738_2717.n1 a_738_2717.t5 168.701
R14795 a_738_2717.t0 a_738_2717.n3 96.1553
R14796 a_738_2717.n3 a_738_2717.t3 65.6672
R14797 a_738_2717.n0 a_738_2717.t1 65.0005
R14798 a_738_2717.n0 a_738_2717.t2 45.0005
R14799 a_n8511_n9484.t0 a_n8511_n9484.t1 60.0005
R14800 a_1866_n5074.t1 a_1866_n5074.n3 370.026
R14801 a_1866_n5074.n0 a_1866_n5074.t3 351.356
R14802 a_1866_n5074.n1 a_1866_n5074.t4 334.717
R14803 a_1866_n5074.n3 a_1866_n5074.t0 325.971
R14804 a_1866_n5074.n1 a_1866_n5074.t2 309.935
R14805 a_1866_n5074.n0 a_1866_n5074.t5 305.683
R14806 a_1866_n5074.n2 a_1866_n5074.n0 16.879
R14807 a_1866_n5074.n3 a_1866_n5074.n2 10.8867
R14808 a_1866_n5074.n2 a_1866_n5074.n1 9.3005
R14809 a_2121_n4714.n1 a_2121_n4714.n0 926.024
R14810 a_2121_n4714.n0 a_2121_n4714.t3 82.0838
R14811 a_2121_n4714.n1 a_2121_n4714.t2 63.3338
R14812 a_2121_n4714.n0 a_2121_n4714.t1 63.3219
R14813 a_2121_n4714.t0 a_2121_n4714.n1 29.7268
R14814 a_2216_n4702.n3 a_2216_n4702.n2 674.338
R14815 a_2216_n4702.n1 a_2216_n4702.t4 332.58
R14816 a_2216_n4702.n2 a_2216_n4702.n0 284.012
R14817 a_2216_n4702.n2 a_2216_n4702.n1 253.648
R14818 a_2216_n4702.n1 a_2216_n4702.t5 168.701
R14819 a_2216_n4702.t0 a_2216_n4702.n3 96.1553
R14820 a_2216_n4702.n3 a_2216_n4702.t3 65.6672
R14821 a_2216_n4702.n0 a_2216_n4702.t1 65.0005
R14822 a_2216_n4702.n0 a_2216_n4702.t2 45.0005
R14823 a_4253_3557.t1 a_4253_3557.n3 370.026
R14824 a_4253_3557.n0 a_4253_3557.t5 351.356
R14825 a_4253_3557.n1 a_4253_3557.t4 334.717
R14826 a_4253_3557.n3 a_4253_3557.t0 325.971
R14827 a_4253_3557.n1 a_4253_3557.t2 309.935
R14828 a_4253_3557.n0 a_4253_3557.t3 305.683
R14829 a_4253_3557.n2 a_4253_3557.n0 16.879
R14830 a_4253_3557.n3 a_4253_3557.n2 10.8867
R14831 a_4253_3557.n2 a_4253_3557.n1 9.3005
R14832 a_1657_2717.t0 a_1657_2717.t1 87.1434
R14833 a_4296_n5482.n1 a_4296_n5482.t4 530.01
R14834 a_4296_n5482.t1 a_4296_n5482.n5 421.021
R14835 a_4296_n5482.n0 a_4296_n5482.t5 337.171
R14836 a_4296_n5482.n3 a_4296_n5482.t0 280.223
R14837 a_4296_n5482.n4 a_4296_n5482.t7 263.173
R14838 a_4296_n5482.n4 a_4296_n5482.t2 227.826
R14839 a_4296_n5482.n0 a_4296_n5482.t6 199.762
R14840 a_4296_n5482.n2 a_4296_n5482.n1 170.81
R14841 a_4296_n5482.n2 a_4296_n5482.n0 167.321
R14842 a_4296_n5482.n5 a_4296_n5482.n4 152
R14843 a_4296_n5482.n1 a_4296_n5482.t3 141.923
R14844 a_4296_n5482.n3 a_4296_n5482.n2 10.8376
R14845 a_4296_n5482.n5 a_4296_n5482.n3 2.50485
R14846 a_2470_n1441.n3 a_2470_n1441.n2 636.953
R14847 a_2470_n1441.n1 a_2470_n1441.t4 366.856
R14848 a_2470_n1441.n2 a_2470_n1441.n0 300.2
R14849 a_2470_n1441.n2 a_2470_n1441.n1 225.036
R14850 a_2470_n1441.n1 a_2470_n1441.t5 174.056
R14851 a_2470_n1441.n0 a_2470_n1441.t2 70.0005
R14852 a_2470_n1441.t0 a_2470_n1441.n3 68.0124
R14853 a_2470_n1441.n3 a_2470_n1441.t3 63.3219
R14854 a_2470_n1441.n0 a_2470_n1441.t1 61.6672
R14855 a_2819_n9650.n3 a_2819_n9650.n2 674.338
R14856 a_2819_n9650.n1 a_2819_n9650.t4 332.58
R14857 a_2819_n9650.n2 a_2819_n9650.n0 284.012
R14858 a_2819_n9650.n2 a_2819_n9650.n1 253.648
R14859 a_2819_n9650.n1 a_2819_n9650.t5 168.701
R14860 a_2819_n9650.t1 a_2819_n9650.n3 96.1553
R14861 a_2819_n9650.n3 a_2819_n9650.t3 65.6672
R14862 a_2819_n9650.n0 a_2819_n9650.t0 65.0005
R14863 a_2819_n9650.n0 a_2819_n9650.t2 45.0005
R14864 a_8686_n4702.n0 a_8686_n4702.t1 68.3338
R14865 a_8686_n4702.n0 a_8686_n4702.t0 26.3935
R14866 a_8686_n4702.n1 a_8686_n4702.n0 14.4005
R14867 a_7177_n1029.t1 a_7177_n1029.t0 94.7268
R14868 a_4256_n5080.t0 a_4256_n5080.n0 1327.82
R14869 a_4256_n5080.n0 a_4256_n5080.t1 194.655
R14870 a_4256_n5080.n0 a_4256_n5080.t2 63.3219
R14871 a_222_2717.n1 a_222_2717.t2 530.01
R14872 a_222_2717.t1 a_222_2717.n5 421.021
R14873 a_222_2717.n0 a_222_2717.t5 337.142
R14874 a_222_2717.n3 a_222_2717.t0 280.223
R14875 a_222_2717.n4 a_222_2717.t4 263.173
R14876 a_222_2717.n4 a_222_2717.t3 227.826
R14877 a_222_2717.n0 a_222_2717.t6 199.762
R14878 a_222_2717.n2 a_222_2717.n1 170.81
R14879 a_222_2717.n2 a_222_2717.n0 167.321
R14880 a_222_2717.n5 a_222_2717.n4 152
R14881 a_222_2717.n1 a_222_2717.t7 141.923
R14882 a_222_2717.n3 a_222_2717.n2 10.8376
R14883 a_222_2717.n5 a_222_2717.n3 2.50485
R14884 a_846_3083.t0 a_846_3083.n0 1327.82
R14885 a_846_3083.n0 a_846_3083.t2 194.655
R14886 a_846_3083.n0 a_846_3083.t1 63.3219
R14887 a_n783_n9662.t0 a_n783_n9662.t1 60.0005
R14888 a_3590_3557.t0 a_3590_3557.t1 87.1434
R14889 a_n8208_n9484.n3 a_n8208_n9484.n2 636.953
R14890 a_n8208_n9484.n1 a_n8208_n9484.t5 366.856
R14891 a_n8208_n9484.n2 a_n8208_n9484.n0 300.2
R14892 a_n8208_n9484.n2 a_n8208_n9484.n1 225.036
R14893 a_n8208_n9484.n1 a_n8208_n9484.t4 174.056
R14894 a_n8208_n9484.n0 a_n8208_n9484.t3 70.0005
R14895 a_n8208_n9484.t0 a_n8208_n9484.n3 68.0124
R14896 a_n8208_n9484.n3 a_n8208_n9484.t2 63.3219
R14897 a_n8208_n9484.n0 a_n8208_n9484.t1 61.6672
R14898 a_2154_2717.n1 a_2154_2717.t4 530.01
R14899 a_2154_2717.t1 a_2154_2717.n5 421.021
R14900 a_2154_2717.n0 a_2154_2717.t2 337.142
R14901 a_2154_2717.n3 a_2154_2717.t0 280.223
R14902 a_2154_2717.n4 a_2154_2717.t6 263.173
R14903 a_2154_2717.n4 a_2154_2717.t5 227.826
R14904 a_2154_2717.n0 a_2154_2717.t7 199.762
R14905 a_2154_2717.n2 a_2154_2717.n1 170.81
R14906 a_2154_2717.n2 a_2154_2717.n0 167.321
R14907 a_2154_2717.n5 a_2154_2717.n4 152
R14908 a_2154_2717.n1 a_2154_2717.t3 141.923
R14909 a_2154_2717.n3 a_2154_2717.n2 10.8376
R14910 a_2154_2717.n5 a_2154_2717.n3 2.50485
R14911 a_4711_3923.t0 a_4711_3923.n0 1327.82
R14912 a_4711_3923.n0 a_4711_3923.t1 194.655
R14913 a_4711_3923.n0 a_4711_3923.t2 63.3219
R14914 a_8653_n787.n3 a_8653_n787.n2 647.119
R14915 a_8653_n787.n1 a_8653_n787.t4 350.253
R14916 a_8653_n787.n2 a_8653_n787.n0 260.339
R14917 a_8653_n787.n2 a_8653_n787.n1 246.119
R14918 a_8653_n787.n1 a_8653_n787.t5 189.588
R14919 a_8653_n787.n3 a_8653_n787.t2 89.1195
R14920 a_8653_n787.n0 a_8653_n787.t3 63.3338
R14921 a_8653_n787.t1 a_8653_n787.n3 41.0422
R14922 a_8653_n787.n0 a_8653_n787.t0 31.9797
R14923 a_8531_n1029.t0 a_8531_n1029.t1 198.571
R14924 a_8697_n1029.t0 a_8697_n1029.t1 60.0005
R14925 a_7662_n5074.t1 a_7662_n5074.n3 370.026
R14926 a_7662_n5074.n0 a_7662_n5074.t5 351.356
R14927 a_7662_n5074.n1 a_7662_n5074.t2 334.717
R14928 a_7662_n5074.n3 a_7662_n5074.t0 325.971
R14929 a_7662_n5074.n1 a_7662_n5074.t4 309.935
R14930 a_7662_n5074.n0 a_7662_n5074.t3 305.683
R14931 a_7662_n5074.n2 a_7662_n5074.n0 16.879
R14932 a_7662_n5074.n3 a_7662_n5074.n2 10.8867
R14933 a_7662_n5074.n2 a_7662_n5074.n1 9.3005
R14934 a_8108_n4702.t0 a_8108_n4702.t1 198.571
R14935 a_8562_2717.t1 a_8562_2717.t0 198.571
R14936 a_8728_2717.t0 a_8728_2717.t1 60.0005
R14937 a_n1710_2717.n1 a_n1710_2717.t3 530.01
R14938 a_n1710_2717.t1 a_n1710_2717.n5 421.021
R14939 a_n1710_2717.n0 a_n1710_2717.t5 337.142
R14940 a_n1710_2717.n3 a_n1710_2717.t0 280.223
R14941 a_n1710_2717.n4 a_n1710_2717.t7 263.173
R14942 a_n1710_2717.n4 a_n1710_2717.t6 227.826
R14943 a_n1710_2717.n0 a_n1710_2717.t4 199.762
R14944 a_n1710_2717.n2 a_n1710_2717.n1 170.81
R14945 a_n1710_2717.n2 a_n1710_2717.n0 167.321
R14946 a_n1710_2717.n5 a_n1710_2717.n4 152
R14947 a_n1710_2717.n1 a_n1710_2717.t2 141.923
R14948 a_n1710_2717.n3 a_n1710_2717.n2 10.8376
R14949 a_n1710_2717.n5 a_n1710_2717.n3 2.50485
R14950 a_n1289_2717.n1 a_n1289_2717.n0 926.024
R14951 a_n1289_2717.t0 a_n1289_2717.n1 82.0838
R14952 a_n1289_2717.n0 a_n1289_2717.t3 63.3338
R14953 a_n1289_2717.n1 a_n1289_2717.t1 63.3219
R14954 a_n1289_2717.n0 a_n1289_2717.t2 29.7268
R14955 a_n1194_2717.n3 a_n1194_2717.n2 674.338
R14956 a_n1194_2717.n1 a_n1194_2717.t5 332.58
R14957 a_n1194_2717.n2 a_n1194_2717.n0 284.012
R14958 a_n1194_2717.n2 a_n1194_2717.n1 253.648
R14959 a_n1194_2717.n1 a_n1194_2717.t4 168.701
R14960 a_n1194_2717.n3 a_n1194_2717.t2 96.1553
R14961 a_n1194_2717.t0 a_n1194_2717.n3 65.6672
R14962 a_n1194_2717.n0 a_n1194_2717.t3 65.0005
R14963 a_n1194_2717.n0 a_n1194_2717.t1 45.0005
R14964 a_6999_n4714.t0 a_6999_n4714.t1 87.1434
R14965 a_6820_n4776.n5 a_6820_n4776.n4 807.871
R14966 a_6820_n4776.n2 a_6820_n4776.t3 389.183
R14967 a_6820_n4776.n3 a_6820_n4776.n2 251.167
R14968 a_6820_n4776.n3 a_6820_n4776.t1 223.571
R14969 a_6820_n4776.n0 a_6820_n4776.t7 212.081
R14970 a_6820_n4776.n1 a_6820_n4776.t8 212.081
R14971 a_6820_n4776.n4 a_6820_n4776.n1 176.576
R14972 a_6820_n4776.n2 a_6820_n4776.t6 174.891
R14973 a_6820_n4776.n0 a_6820_n4776.t4 139.78
R14974 a_6820_n4776.n1 a_6820_n4776.t5 139.78
R14975 a_6820_n4776.n5 a_6820_n4776.t2 63.3219
R14976 a_6820_n4776.t0 a_6820_n4776.n5 63.3219
R14977 a_6820_n4776.n1 a_6820_n4776.n0 61.346
R14978 a_6820_n4776.n4 a_6820_n4776.n3 37.7195
R14979 a_2781_n4702.n3 a_2781_n4702.n2 636.953
R14980 a_2781_n4702.n1 a_2781_n4702.t5 366.856
R14981 a_2781_n4702.n2 a_2781_n4702.n0 300.2
R14982 a_2781_n4702.n2 a_2781_n4702.n1 225.036
R14983 a_2781_n4702.n1 a_2781_n4702.t4 174.056
R14984 a_2781_n4702.n0 a_2781_n4702.t2 70.0005
R14985 a_2781_n4702.t0 a_2781_n4702.n3 68.0124
R14986 a_2781_n4702.n3 a_2781_n4702.t3 63.3219
R14987 a_2781_n4702.n0 a_2781_n4702.t1 61.6672
R14988 a_2956_n4776.n5 a_2956_n4776.n4 807.871
R14989 a_2956_n4776.n2 a_2956_n4776.t5 389.183
R14990 a_2956_n4776.n3 a_2956_n4776.n2 251.167
R14991 a_2956_n4776.n3 a_2956_n4776.t2 223.571
R14992 a_2956_n4776.n0 a_2956_n4776.t3 212.081
R14993 a_2956_n4776.n1 a_2956_n4776.t4 212.081
R14994 a_2956_n4776.n4 a_2956_n4776.n1 176.576
R14995 a_2956_n4776.n2 a_2956_n4776.t7 174.891
R14996 a_2956_n4776.n0 a_2956_n4776.t6 139.78
R14997 a_2956_n4776.n1 a_2956_n4776.t8 139.78
R14998 a_2956_n4776.n5 a_2956_n4776.t1 63.3219
R14999 a_2956_n4776.t0 a_2956_n4776.n5 63.3219
R15000 a_2956_n4776.n1 a_2956_n4776.n0 61.346
R15001 a_2956_n4776.n4 a_2956_n4776.n3 37.7195
R15002 a_n5425_n10022.n1 a_n5425_n10022.t7 530.01
R15003 a_n5425_n10022.t1 a_n5425_n10022.n5 421.021
R15004 a_n5425_n10022.n0 a_n5425_n10022.t5 337.142
R15005 a_n5425_n10022.n3 a_n5425_n10022.t0 280.223
R15006 a_n5425_n10022.n4 a_n5425_n10022.t6 263.173
R15007 a_n5425_n10022.n4 a_n5425_n10022.t3 227.826
R15008 a_n5425_n10022.n0 a_n5425_n10022.t4 199.762
R15009 a_n5425_n10022.n2 a_n5425_n10022.n1 170.81
R15010 a_n5425_n10022.n2 a_n5425_n10022.n0 167.321
R15011 a_n5425_n10022.n5 a_n5425_n10022.n4 152
R15012 a_n5425_n10022.n1 a_n5425_n10022.t2 141.923
R15013 a_n5425_n10022.n3 a_n5425_n10022.n2 10.8376
R15014 a_n5425_n10022.n5 a_n5425_n10022.n3 2.50485
R15015 a_9180_n9650.n3 a_9180_n9650.n2 636.953
R15016 a_9180_n9650.n1 a_9180_n9650.t5 366.856
R15017 a_9180_n9650.n2 a_9180_n9650.n0 300.2
R15018 a_9180_n9650.n2 a_9180_n9650.n1 225.036
R15019 a_9180_n9650.n1 a_9180_n9650.t4 174.056
R15020 a_9180_n9650.n0 a_9180_n9650.t2 70.0005
R15021 a_9180_n9650.t0 a_9180_n9650.n3 68.0124
R15022 a_9180_n9650.n3 a_9180_n9650.t3 63.3219
R15023 a_9180_n9650.n0 a_9180_n9650.t1 61.6672
R15024 a_956_2959.n3 a_956_2959.n2 647.119
R15025 a_956_2959.n1 a_956_2959.t4 350.253
R15026 a_956_2959.n2 a_956_2959.n0 260.339
R15027 a_956_2959.n2 a_956_2959.n1 246.119
R15028 a_956_2959.n1 a_956_2959.t5 189.588
R15029 a_956_2959.n3 a_956_2959.t3 89.1195
R15030 a_956_2959.n0 a_956_2959.t2 63.3338
R15031 a_956_2959.t1 a_956_2959.n3 41.0422
R15032 a_956_2959.n0 a_956_2959.t0 31.9797
R15033 a_834_2717.t0 a_834_2717.t1 198.571
R15034 a_1000_2717.t0 a_1000_2717.t1 60.0005
R15035 a_537_n10022.t1 a_537_n10022.n3 370.026
R15036 a_537_n10022.n0 a_537_n10022.t5 351.356
R15037 a_537_n10022.n1 a_537_n10022.t3 334.717
R15038 a_537_n10022.n3 a_537_n10022.t0 325.971
R15039 a_537_n10022.n1 a_537_n10022.t2 309.935
R15040 a_537_n10022.n0 a_537_n10022.t4 305.683
R15041 a_537_n10022.n2 a_537_n10022.n0 16.879
R15042 a_537_n10022.n3 a_537_n10022.n2 10.8867
R15043 a_537_n10022.n2 a_537_n10022.n1 9.3005
R15044 a_432_n5482.n1 a_432_n5482.t2 530.01
R15045 a_432_n5482.t1 a_432_n5482.n5 421.021
R15046 a_432_n5482.n0 a_432_n5482.t4 337.171
R15047 a_432_n5482.n3 a_432_n5482.t0 280.223
R15048 a_432_n5482.n4 a_432_n5482.t3 263.173
R15049 a_432_n5482.n4 a_432_n5482.t5 227.826
R15050 a_432_n5482.n0 a_432_n5482.t6 199.762
R15051 a_432_n5482.n2 a_432_n5482.n1 170.81
R15052 a_432_n5482.n2 a_432_n5482.n0 167.321
R15053 a_432_n5482.n5 a_432_n5482.n4 152
R15054 a_432_n5482.n1 a_432_n5482.t7 141.923
R15055 a_432_n5482.n3 a_432_n5482.n2 10.8376
R15056 a_432_n5482.n5 a_432_n5482.n3 2.50485
R15057 a_588_n5387.n3 a_588_n5387.n2 674.338
R15058 a_588_n5387.n1 a_588_n5387.t4 332.58
R15059 a_588_n5387.n2 a_588_n5387.n0 284.012
R15060 a_588_n5387.n2 a_588_n5387.n1 253.648
R15061 a_588_n5387.n1 a_588_n5387.t5 168.701
R15062 a_588_n5387.t1 a_588_n5387.n3 96.1553
R15063 a_588_n5387.n3 a_588_n5387.t3 65.6672
R15064 a_588_n5387.n0 a_588_n5387.t0 65.0005
R15065 a_588_n5387.n0 a_588_n5387.t2 45.0005
R15066 a_6612_n1457.t1 a_6612_n1457.n3 370.026
R15067 a_6612_n1457.n0 a_6612_n1457.t4 351.356
R15068 a_6612_n1457.n1 a_6612_n1457.t2 334.717
R15069 a_6612_n1457.n3 a_6612_n1457.t0 325.971
R15070 a_6612_n1457.n1 a_6612_n1457.t5 309.935
R15071 a_6612_n1457.n0 a_6612_n1457.t3 305.683
R15072 a_6612_n1457.n2 a_6612_n1457.n0 16.879
R15073 a_6612_n1457.n3 a_6612_n1457.n2 10.8867
R15074 a_6612_n1457.n2 a_6612_n1457.n1 9.3005
R15075 auto_sampling_0.x2.D.n5 auto_sampling_0.x2.D.n4 585
R15076 auto_sampling_0.x2.D.n4 auto_sampling_0.x2.D.n3 585
R15077 auto_sampling_0.x2.D.n2 auto_sampling_0.x2.D.t4 333.651
R15078 auto_sampling_0.x2.D.n2 auto_sampling_0.x2.D.t5 297.233
R15079 auto_sampling_0.x2.D auto_sampling_0.x2.D.n2 196.493
R15080 auto_sampling_0.x2.D.n1 auto_sampling_0.x2.D.n0 185
R15081 auto_sampling_0.x2.D auto_sampling_0.x2.D.n1 49.0339
R15082 auto_sampling_0.x2.D.n3 auto_sampling_0.x2.D 44.2533
R15083 auto_sampling_0.x2.D.n4 auto_sampling_0.x2.D.t3 26.5955
R15084 auto_sampling_0.x2.D.n4 auto_sampling_0.x2.D.t2 26.5955
R15085 auto_sampling_0.x2.D.n0 auto_sampling_0.x2.D.t1 24.9236
R15086 auto_sampling_0.x2.D.n0 auto_sampling_0.x2.D.t0 24.9236
R15087 auto_sampling_0.x2.D.n5 auto_sampling_0.x2.D 15.6165
R15088 auto_sampling_0.x2.D.n1 auto_sampling_0.x2.D 10.4965
R15089 auto_sampling_0.x2.D.n3 auto_sampling_0.x2.D 1.7925
R15090 auto_sampling_0.x2.D auto_sampling_0.x2.D.n5 1.7925
R15091 a_2639_n1029.n3 a_2639_n1029.n2 674.338
R15092 a_2639_n1029.n1 a_2639_n1029.t5 332.58
R15093 a_2639_n1029.n2 a_2639_n1029.n0 284.012
R15094 a_2639_n1029.n2 a_2639_n1029.n1 253.648
R15095 a_2639_n1029.n1 a_2639_n1029.t4 168.701
R15096 a_2639_n1029.t2 a_2639_n1029.n3 96.1553
R15097 a_2639_n1029.n3 a_2639_n1029.t3 65.6672
R15098 a_2639_n1029.n0 a_2639_n1029.t1 65.0005
R15099 a_2639_n1029.n0 a_2639_n1029.t0 45.0005
R15100 a_2857_n787.n3 a_2857_n787.n2 647.119
R15101 a_2857_n787.n1 a_2857_n787.t4 350.253
R15102 a_2857_n787.n2 a_2857_n787.n0 260.339
R15103 a_2857_n787.n2 a_2857_n787.n1 246.119
R15104 a_2857_n787.n1 a_2857_n787.t5 189.588
R15105 a_2857_n787.n3 a_2857_n787.t3 89.1195
R15106 a_2857_n787.n0 a_2857_n787.t0 63.3338
R15107 a_2857_n787.t2 a_2857_n787.n3 41.0422
R15108 a_2857_n787.n0 a_2857_n787.t1 31.9797
R15109 a_6145_n5258.t0 a_6145_n5258.t1 126.644
R15110 a_2321_3557.t1 a_2321_3557.n3 370.026
R15111 a_2321_3557.n0 a_2321_3557.t2 351.356
R15112 a_2321_3557.n1 a_2321_3557.t5 334.717
R15113 a_2321_3557.n3 a_2321_3557.t0 325.971
R15114 a_2321_3557.n1 a_2321_3557.t3 309.935
R15115 a_2321_3557.n0 a_2321_3557.t4 305.683
R15116 a_2321_3557.n2 a_2321_3557.n0 16.879
R15117 a_2321_3557.n3 a_2321_3557.n2 10.8867
R15118 a_2321_3557.n2 a_2321_3557.n1 9.3005
R15119 a_6588_n9662.n1 a_6588_n9662.n0 926.024
R15120 a_6588_n9662.t1 a_6588_n9662.n1 82.0838
R15121 a_6588_n9662.n0 a_6588_n9662.t0 63.3338
R15122 a_6588_n9662.n1 a_6588_n9662.t3 63.3219
R15123 a_6588_n9662.n0 a_6588_n9662.t2 29.7268
R15124 a_6683_n9650.n3 a_6683_n9650.n2 674.338
R15125 a_6683_n9650.n1 a_6683_n9650.t5 332.58
R15126 a_6683_n9650.n2 a_6683_n9650.n0 284.012
R15127 a_6683_n9650.n2 a_6683_n9650.n1 253.648
R15128 a_6683_n9650.n1 a_6683_n9650.t4 168.701
R15129 a_6683_n9650.t1 a_6683_n9650.n3 96.1553
R15130 a_6683_n9650.n3 a_6683_n9650.t2 65.6672
R15131 a_6683_n9650.n0 a_6683_n9650.t0 65.0005
R15132 a_6683_n9650.n0 a_6683_n9650.t3 45.0005
R15133 a_n4909_n9484.n3 a_n4909_n9484.n2 674.338
R15134 a_n4909_n9484.n1 a_n4909_n9484.t4 332.58
R15135 a_n4909_n9484.n2 a_n4909_n9484.n0 284.012
R15136 a_n4909_n9484.n2 a_n4909_n9484.n1 253.648
R15137 a_n4909_n9484.n1 a_n4909_n9484.t5 168.701
R15138 a_n4909_n9484.n3 a_n4909_n9484.t3 96.1553
R15139 a_n4909_n9484.t0 a_n4909_n9484.n3 65.6672
R15140 a_n4909_n9484.n0 a_n4909_n9484.t2 65.0005
R15141 a_n4909_n9484.n0 a_n4909_n9484.t1 45.0005
R15142 a_n4813_n9484.t1 a_n4813_n9484.t0 198.571
R15143 a_n3072_n9662.n1 a_n3072_n9662.n0 926.024
R15144 a_n3072_n9662.t0 a_n3072_n9662.n1 82.0838
R15145 a_n3072_n9662.n0 a_n3072_n9662.t1 63.3338
R15146 a_n3072_n9662.n1 a_n3072_n9662.t3 63.3219
R15147 a_n3072_n9662.n0 a_n3072_n9662.t2 29.7268
R15148 a_8085_n1029.t1 a_8085_n1029.n3 370.026
R15149 a_8085_n1029.n0 a_8085_n1029.t5 351.356
R15150 a_8085_n1029.n1 a_8085_n1029.t3 334.717
R15151 a_8085_n1029.n3 a_8085_n1029.t0 325.971
R15152 a_8085_n1029.n1 a_8085_n1029.t2 309.935
R15153 a_8085_n1029.n0 a_8085_n1029.t4 305.683
R15154 a_8085_n1029.n2 a_8085_n1029.n0 16.879
R15155 a_8085_n1029.n3 a_8085_n1029.n2 10.8867
R15156 a_8085_n1029.n2 a_8085_n1029.n1 9.3005
R15157 a_8340_n1029.n1 a_8340_n1029.n0 926.024
R15158 a_8340_n1029.t0 a_8340_n1029.n1 82.0838
R15159 a_8340_n1029.n0 a_8340_n1029.t3 63.3338
R15160 a_8340_n1029.n1 a_8340_n1029.t2 63.3219
R15161 a_8340_n1029.n0 a_8340_n1029.t1 29.7268
R15162 a_8435_n1029.n3 a_8435_n1029.n2 674.338
R15163 a_8435_n1029.n1 a_8435_n1029.t5 332.58
R15164 a_8435_n1029.n2 a_8435_n1029.n0 284.012
R15165 a_8435_n1029.n2 a_8435_n1029.n1 253.648
R15166 a_8435_n1029.n1 a_8435_n1029.t4 168.701
R15167 a_8435_n1029.n3 a_8435_n1029.t2 96.1553
R15168 a_8435_n1029.t1 a_8435_n1029.n3 65.6672
R15169 a_8435_n1029.n0 a_8435_n1029.t3 65.0005
R15170 a_8435_n1029.n0 a_8435_n1029.t0 45.0005
R15171 a_6588_n9484.n1 a_6588_n9484.n0 926.024
R15172 a_6588_n9484.n0 a_6588_n9484.t3 82.0838
R15173 a_6588_n9484.n1 a_6588_n9484.t2 63.3338
R15174 a_6588_n9484.n0 a_6588_n9484.t1 63.3219
R15175 a_6588_n9484.n2 a_6588_n9484.t0 26.3935
R15176 a_6588_n9484.n3 a_6588_n9484.n2 14.4005
R15177 a_6588_n9484.n2 a_6588_n9484.n1 3.33383
R15178 a_2544_n1029.n1 a_2544_n1029.n0 926.024
R15179 a_2544_n1029.n0 a_2544_n1029.t3 82.0838
R15180 a_2544_n1029.n1 a_2544_n1029.t2 63.3338
R15181 a_2544_n1029.n0 a_2544_n1029.t1 63.3219
R15182 a_2544_n1029.n2 a_2544_n1029.t0 26.3935
R15183 a_2544_n1029.n3 a_2544_n1029.n2 14.4005
R15184 a_2544_n1029.n2 a_2544_n1029.n1 3.33383
R15185 a_612_n1029.n1 a_612_n1029.n0 926.024
R15186 a_612_n1029.n0 a_612_n1029.t3 82.0838
R15187 a_612_n1029.n1 a_612_n1029.t2 63.3338
R15188 a_612_n1029.n0 a_612_n1029.t1 63.3219
R15189 a_612_n1029.n2 a_612_n1029.t0 26.3935
R15190 a_612_n1029.n3 a_612_n1029.n2 14.4005
R15191 a_612_n1029.n2 a_612_n1029.n1 3.33383
R15192 a_707_n1029.n3 a_707_n1029.n2 674.338
R15193 a_707_n1029.n1 a_707_n1029.t5 332.58
R15194 a_707_n1029.n2 a_707_n1029.n0 284.012
R15195 a_707_n1029.n2 a_707_n1029.n1 253.648
R15196 a_707_n1029.n1 a_707_n1029.t4 168.701
R15197 a_707_n1029.t0 a_707_n1029.n3 96.1553
R15198 a_707_n1029.n3 a_707_n1029.t3 65.6672
R15199 a_707_n1029.n0 a_707_n1029.t1 65.0005
R15200 a_707_n1029.n0 a_707_n1029.t2 45.0005
R15201 a_6694_n5624.t1 a_6694_n5624.t0 198.571
R15202 a_6752_2959.n3 a_6752_2959.n2 647.119
R15203 a_6752_2959.n1 a_6752_2959.t5 350.253
R15204 a_6752_2959.n2 a_6752_2959.n0 260.339
R15205 a_6752_2959.n2 a_6752_2959.n1 246.119
R15206 a_6752_2959.n1 a_6752_2959.t4 189.588
R15207 a_6752_2959.n3 a_6752_2959.t0 89.1195
R15208 a_6752_2959.n0 a_6752_2959.t3 63.3338
R15209 a_6752_2959.t2 a_6752_2959.n3 41.0422
R15210 a_6752_2959.n0 a_6752_2959.t1 31.9797
R15211 a_n3327_n9484.t1 a_n3327_n9484.n3 370.026
R15212 a_n3327_n9484.n0 a_n3327_n9484.t5 351.356
R15213 a_n3327_n9484.n1 a_n3327_n9484.t3 334.717
R15214 a_n3327_n9484.n3 a_n3327_n9484.t0 325.971
R15215 a_n3327_n9484.n1 a_n3327_n9484.t4 309.935
R15216 a_n3327_n9484.n0 a_n3327_n9484.t2 305.683
R15217 a_n3327_n9484.n2 a_n3327_n9484.n0 16.879
R15218 a_n3327_n9484.n3 a_n3327_n9484.n2 10.8867
R15219 a_n3327_n9484.n2 a_n3327_n9484.n1 9.3005
R15220 a_n9123_n9484.t1 a_n9123_n9484.n3 370.026
R15221 a_n9123_n9484.n0 a_n9123_n9484.t2 351.356
R15222 a_n9123_n9484.n1 a_n9123_n9484.t5 334.717
R15223 a_n9123_n9484.n3 a_n9123_n9484.t0 325.971
R15224 a_n9123_n9484.n1 a_n9123_n9484.t4 309.935
R15225 a_n9123_n9484.n0 a_n9123_n9484.t3 305.683
R15226 a_n9123_n9484.n2 a_n9123_n9484.n0 16.879
R15227 a_n9123_n9484.n3 a_n9123_n9484.n2 10.8867
R15228 a_n9123_n9484.n2 a_n9123_n9484.n1 9.3005
R15229 a_5342_2691.n5 a_5342_2691.n4 807.871
R15230 a_5342_2691.n2 a_5342_2691.t4 389.183
R15231 a_5342_2691.n3 a_5342_2691.n2 251.167
R15232 a_5342_2691.n3 a_5342_2691.t1 223.571
R15233 a_5342_2691.n0 a_5342_2691.t6 212.081
R15234 a_5342_2691.n1 a_5342_2691.t8 212.081
R15235 a_5342_2691.n4 a_5342_2691.n1 176.576
R15236 a_5342_2691.n2 a_5342_2691.t3 174.891
R15237 a_5342_2691.n0 a_5342_2691.t7 139.78
R15238 a_5342_2691.n1 a_5342_2691.t5 139.78
R15239 a_5342_2691.n5 a_5342_2691.t2 63.3219
R15240 a_5342_2691.t0 a_5342_2691.n5 63.3219
R15241 a_5342_2691.n1 a_5342_2691.n0 61.346
R15242 a_5342_2691.n4 a_5342_2691.n3 37.7195
R15243 auto_sampling_0.x11.Q.n6 auto_sampling_0.x11.Q.n5 289.096
R15244 auto_sampling_0.x11.Q.n2 auto_sampling_0.x11.Q.t4 230.576
R15245 auto_sampling_0.x11.Q.n1 auto_sampling_0.x11.Q.n0 185
R15246 auto_sampling_0.x11.Q.n2 auto_sampling_0.x11.Q.t5 158.275
R15247 auto_sampling_0.x11.Q.n3 auto_sampling_0.x11.Q.n2 152
R15248 auto_sampling_0.x11.Q.n4 auto_sampling_0.x11.Q.n1 31.2387
R15249 auto_sampling_0.x11.Q.n5 auto_sampling_0.x11.Q.t3 26.5955
R15250 auto_sampling_0.x11.Q.n5 auto_sampling_0.x11.Q.t2 26.5955
R15251 auto_sampling_0.x11.Q.n0 auto_sampling_0.x11.Q.t0 24.9236
R15252 auto_sampling_0.x11.Q.n0 auto_sampling_0.x11.Q.t1 24.9236
R15253 auto_sampling_0.x11.Q.n4 auto_sampling_0.x11.Q.n3 19.3721
R15254 auto_sampling_0.x11.Q auto_sampling_0.x11.Q.n4 17.7956
R15255 auto_sampling_0.x11.Q.n1 auto_sampling_0.x11.Q 10.4965
R15256 auto_sampling_0.x11.Q auto_sampling_0.x11.Q.n6 9.48653
R15257 auto_sampling_0.x11.Q.n6 auto_sampling_0.x11.Q 7.7181
R15258 auto_sampling_0.x11.Q.n3 auto_sampling_0.x11.Q 6.66717
R15259 a_7209_3557.t0 a_7209_3557.t1 94.7268
R15260 a_n305_n9724.n4 a_n305_n9724.n1 807.871
R15261 a_n305_n9724.n0 a_n305_n9724.t3 389.183
R15262 a_n305_n9724.n5 a_n305_n9724.n0 251.167
R15263 a_n305_n9724.t0 a_n305_n9724.n5 223.571
R15264 a_n305_n9724.n2 a_n305_n9724.t7 212.081
R15265 a_n305_n9724.n3 a_n305_n9724.t4 212.081
R15266 a_n305_n9724.n4 a_n305_n9724.n3 176.576
R15267 a_n305_n9724.n0 a_n305_n9724.t5 174.891
R15268 a_n305_n9724.n2 a_n305_n9724.t8 139.78
R15269 a_n305_n9724.n3 a_n305_n9724.t6 139.78
R15270 a_n305_n9724.n1 a_n305_n9724.t1 63.3219
R15271 a_n305_n9724.n1 a_n305_n9724.t2 63.3219
R15272 a_n305_n9724.n3 a_n305_n9724.n2 61.346
R15273 a_n305_n9724.n5 a_n305_n9724.n4 37.7195
R15274 a_n318_n10028.t0 a_n318_n10028.t1 126.644
R15275 DOUT[3].n3 DOUT[3].n2 585
R15276 DOUT[3].n4 DOUT[3].n3 585
R15277 DOUT[3].n1 DOUT[3].n0 185
R15278 DOUT[3] DOUT[3].n1 57.7379
R15279 DOUT[3].n3 DOUT[3].t3 26.5955
R15280 DOUT[3].n3 DOUT[3].t2 26.5955
R15281 DOUT[3].n0 DOUT[3].t1 24.9236
R15282 DOUT[3].n0 DOUT[3].t0 24.9236
R15283 DOUT[3] DOUT[3].n5 17.8924
R15284 DOUT[3].n2 DOUT[3] 10.4965
R15285 DOUT[3].n4 DOUT[3] 10.4965
R15286 DOUT[3].n2 DOUT[3] 6.9125
R15287 DOUT[3].n5 DOUT[3] 4.3525
R15288 DOUT[3].n5 DOUT[3].n4 2.5605
R15289 DOUT[3].n1 DOUT[3] 1.7925
R15290 a_7919_n1029.n1 a_7919_n1029.t2 530.01
R15291 a_7919_n1029.t1 a_7919_n1029.n5 421.021
R15292 a_7919_n1029.n0 a_7919_n1029.t5 337.142
R15293 a_7919_n1029.n3 a_7919_n1029.t0 280.223
R15294 a_7919_n1029.n4 a_7919_n1029.t7 263.173
R15295 a_7919_n1029.n4 a_7919_n1029.t4 227.826
R15296 a_7919_n1029.n0 a_7919_n1029.t6 199.762
R15297 a_7919_n1029.n2 a_7919_n1029.n1 170.81
R15298 a_7919_n1029.n2 a_7919_n1029.n0 167.321
R15299 a_7919_n1029.n5 a_7919_n1029.n4 152
R15300 a_7919_n1029.n1 a_7919_n1029.t3 141.923
R15301 a_7919_n1029.n3 a_7919_n1029.n2 10.8376
R15302 a_7919_n1029.n5 a_7919_n1029.n3 2.50485
R15303 a_8543_n663.n0 a_8543_n663.t2 1327.82
R15304 a_8543_n663.t0 a_8543_n663.n0 194.655
R15305 a_8543_n663.n0 a_8543_n663.t1 63.3219
R15306 a_5276_2717.t1 a_5276_2717.t0 94.7268
R15307 auto_sampling_0.x16.D.n5 auto_sampling_0.x16.D.n4 585
R15308 auto_sampling_0.x16.D.n4 auto_sampling_0.x16.D.n3 585
R15309 auto_sampling_0.x16.D.n2 auto_sampling_0.x16.D.t5 333.651
R15310 auto_sampling_0.x16.D.n2 auto_sampling_0.x16.D.t4 297.233
R15311 auto_sampling_0.x16.D auto_sampling_0.x16.D.n2 196.493
R15312 auto_sampling_0.x16.D.n1 auto_sampling_0.x16.D.n0 185
R15313 auto_sampling_0.x16.D auto_sampling_0.x16.D.n1 49.0339
R15314 auto_sampling_0.x16.D.n3 auto_sampling_0.x16.D 44.2533
R15315 auto_sampling_0.x16.D.n4 auto_sampling_0.x16.D.t3 26.5955
R15316 auto_sampling_0.x16.D.n4 auto_sampling_0.x16.D.t2 26.5955
R15317 auto_sampling_0.x16.D.n0 auto_sampling_0.x16.D.t0 24.9236
R15318 auto_sampling_0.x16.D.n0 auto_sampling_0.x16.D.t1 24.9236
R15319 auto_sampling_0.x16.D.n5 auto_sampling_0.x16.D 15.6165
R15320 auto_sampling_0.x16.D.n1 auto_sampling_0.x16.D 10.4965
R15321 auto_sampling_0.x16.D.n3 auto_sampling_0.x16.D 1.7925
R15322 auto_sampling_0.x16.D auto_sampling_0.x16.D.n5 1.7925
R15323 a_6439_2717.n1 a_6439_2717.n0 926.024
R15324 a_6439_2717.n0 a_6439_2717.t3 82.0838
R15325 a_6439_2717.n1 a_6439_2717.t0 63.3338
R15326 a_6439_2717.n0 a_6439_2717.t2 63.3219
R15327 a_6439_2717.n2 a_6439_2717.t1 26.3935
R15328 a_6439_2717.n3 a_6439_2717.n2 14.4005
R15329 a_6439_2717.n2 a_6439_2717.n1 3.33383
R15330 a_2915_n9484.t0 a_2915_n9484.t1 198.571
R15331 a_n949_n9650.t1 a_n949_n9650.t0 198.571
R15332 SWP[6].n0 SWP[6].t5 332.312
R15333 SWP[6].n0 SWP[6].t4 295.627
R15334 SWP[6].n4 SWP[6].n3 289.096
R15335 SWP[6] SWP[6].n0 196.004
R15336 SWP[6].n6 SWP[6].n5 185
R15337 SWP[6] SWP[6].n6 49.0339
R15338 SWP[6].n1 SWP[6] 41.1202
R15339 SWP[6].n2 SWP[6] 35.3521
R15340 SWP[6].n3 SWP[6].t2 26.5955
R15341 SWP[6].n3 SWP[6].t3 26.5955
R15342 SWP[6].n5 SWP[6].t0 24.9236
R15343 SWP[6].n5 SWP[6].t1 24.9236
R15344 SWP[6] SWP[6].n7 14.6049
R15345 SWP[6].n7 SWP[6] 13.0565
R15346 SWP[6].n2 SWP[6].n1 12.9918
R15347 SWP[6] SWP[6].n2 12.026
R15348 SWP[6].n6 SWP[6] 10.4965
R15349 SWP[6] SWP[6].n4 9.48653
R15350 SWP[6].n4 SWP[6] 7.7181
R15351 SWP[6].n7 SWP[6] 4.3525
R15352 SWP[6].n1 SWP[6] 0.0034375
R15353 a_6901_n9242.n3 a_6901_n9242.n2 647.119
R15354 a_6901_n9242.n1 a_6901_n9242.t5 350.253
R15355 a_6901_n9242.n2 a_6901_n9242.n0 260.339
R15356 a_6901_n9242.n2 a_6901_n9242.n1 246.119
R15357 a_6901_n9242.n1 a_6901_n9242.t4 189.588
R15358 a_6901_n9242.n3 a_6901_n9242.t0 89.1195
R15359 a_6901_n9242.n0 a_6901_n9242.t1 63.3338
R15360 a_6901_n9242.t3 a_6901_n9242.n3 41.0422
R15361 a_6901_n9242.n0 a_6901_n9242.t2 31.9797
R15362 a_n8773_n9650.n3 a_n8773_n9650.n2 674.338
R15363 a_n8773_n9650.n1 a_n8773_n9650.t4 332.58
R15364 a_n8773_n9650.n2 a_n8773_n9650.n0 284.012
R15365 a_n8773_n9650.n2 a_n8773_n9650.n1 253.648
R15366 a_n8773_n9650.n1 a_n8773_n9650.t5 168.701
R15367 a_n8773_n9650.t0 a_n8773_n9650.n3 96.1553
R15368 a_n8773_n9650.n3 a_n8773_n9650.t3 65.6672
R15369 a_n8773_n9650.n0 a_n8773_n9650.t1 65.0005
R15370 a_n8773_n9650.n0 a_n8773_n9650.t2 45.0005
R15371 a_n8665_n10028.n0 a_n8665_n10028.t2 1327.82
R15372 a_n8665_n10028.t0 a_n8665_n10028.n0 194.655
R15373 a_n8665_n10028.n0 a_n8665_n10028.t1 63.3219
R15374 SWP[9].n0 SWP[9].t5 333.651
R15375 SWP[9].n0 SWP[9].t4 297.233
R15376 SWP[9].n3 SWP[9].n2 289.096
R15377 SWP[9].n1 SWP[9].n0 196.493
R15378 SWP[9].n5 SWP[9].n4 185
R15379 SWP[9] SWP[9].n5 49.0339
R15380 SWP[9].n8 SWP[9].n1 39.5118
R15381 SWP[9].n7 SWP[9] 28.7841
R15382 SWP[9].n2 SWP[9].t3 26.5955
R15383 SWP[9].n2 SWP[9].t2 26.5955
R15384 SWP[9].n4 SWP[9].t1 24.9236
R15385 SWP[9].n4 SWP[9].t0 24.9236
R15386 SWP[9].n8 SWP[9].n7 18.2035
R15387 SWP[9] SWP[9].n6 14.6135
R15388 SWP[9].n6 SWP[9] 13.0565
R15389 SWP[9].n5 SWP[9] 10.4965
R15390 SWP[9] SWP[9].n3 9.48653
R15391 SWP[9].n3 SWP[9] 7.7181
R15392 SWP[9].n7 SWP[9] 4.61472
R15393 SWP[9].n6 SWP[9] 4.3525
R15394 SWP[9].n1 SWP[9] 0.24431
R15395 SWP[9] SWP[9].n8 0.0057875
R15396 a_7917_n4714.n1 a_7917_n4714.n0 926.024
R15397 a_7917_n4714.n0 a_7917_n4714.t3 82.0838
R15398 a_7917_n4714.n1 a_7917_n4714.t2 63.3338
R15399 a_7917_n4714.n0 a_7917_n4714.t1 63.3219
R15400 a_7917_n4714.t0 a_7917_n4714.n1 29.7268
R15401 a_7117_n1207.t1 a_7117_n1207.t0 198.571
R15402 a_6807_n1599.n3 a_6807_n1599.n2 674.338
R15403 a_6807_n1599.n1 a_6807_n1599.t4 332.58
R15404 a_6807_n1599.n2 a_6807_n1599.n0 284.012
R15405 a_6807_n1599.n2 a_6807_n1599.n1 253.648
R15406 a_6807_n1599.n1 a_6807_n1599.t5 168.701
R15407 a_6807_n1599.n3 a_6807_n1599.t2 96.1553
R15408 a_6807_n1599.t0 a_6807_n1599.n3 65.6672
R15409 a_6807_n1599.n0 a_6807_n1599.t3 65.0005
R15410 a_6807_n1599.n0 a_6807_n1599.t1 45.0005
R15411 a_983_n9650.t0 a_983_n9650.t1 198.571
R15412 a_3798_n5074.t1 a_3798_n5074.n3 370.026
R15413 a_3798_n5074.n0 a_3798_n5074.t5 351.356
R15414 a_3798_n5074.n1 a_3798_n5074.t4 334.717
R15415 a_3798_n5074.n3 a_3798_n5074.t0 325.971
R15416 a_3798_n5074.n1 a_3798_n5074.t2 309.935
R15417 a_3798_n5074.n0 a_3798_n5074.t3 305.683
R15418 a_3798_n5074.n2 a_3798_n5074.n0 16.879
R15419 a_3798_n5074.n3 a_3798_n5074.n2 10.8867
R15420 a_3798_n5074.n2 a_3798_n5074.n1 9.3005
R15421 a_4053_n4714.n1 a_4053_n4714.n0 926.024
R15422 a_4053_n4714.n0 a_4053_n4714.t3 82.0838
R15423 a_4053_n4714.n1 a_4053_n4714.t0 63.3338
R15424 a_4053_n4714.n0 a_4053_n4714.t2 63.3219
R15425 a_4053_n4714.t1 a_4053_n4714.n1 29.7268
R15426 a_4148_n4702.n3 a_4148_n4702.n2 674.338
R15427 a_4148_n4702.n1 a_4148_n4702.t5 332.58
R15428 a_4148_n4702.n2 a_4148_n4702.n0 284.012
R15429 a_4148_n4702.n2 a_4148_n4702.n1 253.648
R15430 a_4148_n4702.n1 a_4148_n4702.t4 168.701
R15431 a_4148_n4702.t0 a_4148_n4702.n3 96.1553
R15432 a_4148_n4702.n3 a_4148_n4702.t2 65.6672
R15433 a_4148_n4702.n0 a_4148_n4702.t1 65.0005
R15434 a_4148_n4702.n0 a_4148_n4702.t3 45.0005
R15435 auto_sampling_0.x12.D.n0 auto_sampling_0.x12.D.t3 333.651
R15436 auto_sampling_0.x12.D.n0 auto_sampling_0.x12.D.t2 297.233
R15437 auto_sampling_0.x12.D.n1 auto_sampling_0.x12.D.t1 233.815
R15438 auto_sampling_0.x12.D auto_sampling_0.x12.D.n0 196.493
R15439 auto_sampling_0.x12.D auto_sampling_0.x12.D.t0 152.889
R15440 auto_sampling_0.x12.D.n1 auto_sampling_0.x12.D 83.172
R15441 auto_sampling_0.x12.D.n2 auto_sampling_0.x12.D 2.22659
R15442 auto_sampling_0.x12.D.n2 auto_sampling_0.x12.D.n1 1.74595
R15443 auto_sampling_0.x12.D auto_sampling_0.x12.D.n2 1.55202
R15444 a_n318_n9118.t0 a_n318_n9118.t1 126.644
R15445 a_826_n5624.t0 a_826_n5624.t1 60.0005
R15446 a_1700_n5074.n1 a_1700_n5074.t3 530.01
R15447 a_1700_n5074.t1 a_1700_n5074.n5 421.021
R15448 a_1700_n5074.n0 a_1700_n5074.t6 337.142
R15449 a_1700_n5074.n3 a_1700_n5074.t0 280.223
R15450 a_1700_n5074.n4 a_1700_n5074.t7 263.173
R15451 a_1700_n5074.n4 a_1700_n5074.t4 227.826
R15452 a_1700_n5074.n0 a_1700_n5074.t2 199.762
R15453 a_1700_n5074.n2 a_1700_n5074.n1 170.81
R15454 a_1700_n5074.n2 a_1700_n5074.n0 167.321
R15455 a_1700_n5074.n5 a_1700_n5074.n4 152
R15456 a_1700_n5074.n1 a_1700_n5074.t5 141.923
R15457 a_1700_n5074.n3 a_1700_n5074.n2 10.8376
R15458 a_1700_n5074.n5 a_1700_n5074.n3 2.50485
R15459 a_2890_n4702.n0 a_2890_n4702.t0 68.3338
R15460 a_2890_n4702.n0 a_2890_n4702.t1 26.3935
R15461 a_2890_n4702.n1 a_2890_n4702.n0 14.4005
R15462 a_2766_2717.t1 a_2766_2717.t0 198.571
R15463 a_2932_2717.t0 a_2932_2717.t1 60.0005
R15464 a_n6733_n10028.t0 a_n6733_n10028.n0 1327.82
R15465 a_n6733_n10028.n0 a_n6733_n10028.t1 194.655
R15466 a_n6733_n10028.n0 a_n6733_n10028.t2 63.3219
R15467 a_4437_n1207.t0 a_4437_n1207.t1 87.1434
R15468 a_6631_3557.t1 a_6631_3557.t0 198.571
R15469 a_n1045_n9650.n3 a_n1045_n9650.n2 674.338
R15470 a_n1045_n9650.n1 a_n1045_n9650.t4 332.58
R15471 a_n1045_n9650.n2 a_n1045_n9650.n0 284.012
R15472 a_n1045_n9650.n2 a_n1045_n9650.n1 253.648
R15473 a_n1045_n9650.n1 a_n1045_n9650.t5 168.701
R15474 a_n1045_n9650.n3 a_n1045_n9650.t2 96.1553
R15475 a_n1045_n9650.t1 a_n1045_n9650.n3 65.6672
R15476 a_n1045_n9650.n0 a_n1045_n9650.t3 65.0005
R15477 a_n1045_n9650.n0 a_n1045_n9650.t0 45.0005
R15478 a_n2412_n9484.n3 a_n2412_n9484.n2 636.953
R15479 a_n2412_n9484.n1 a_n2412_n9484.t4 366.856
R15480 a_n2412_n9484.n2 a_n2412_n9484.n0 300.2
R15481 a_n2412_n9484.n2 a_n2412_n9484.n1 225.036
R15482 a_n2412_n9484.n1 a_n2412_n9484.t5 174.056
R15483 a_n2412_n9484.n0 a_n2412_n9484.t1 70.0005
R15484 a_n2412_n9484.n3 a_n2412_n9484.t3 68.0124
R15485 a_n2412_n9484.t0 a_n2412_n9484.n3 63.3219
R15486 a_n2412_n9484.n0 a_n2412_n9484.t2 61.6672
R15487 a_n7191_n9484.t1 a_n7191_n9484.n3 370.026
R15488 a_n7191_n9484.n0 a_n7191_n9484.t3 351.356
R15489 a_n7191_n9484.n1 a_n7191_n9484.t5 334.717
R15490 a_n7191_n9484.n3 a_n7191_n9484.t0 325.971
R15491 a_n7191_n9484.n1 a_n7191_n9484.t2 309.935
R15492 a_n7191_n9484.n0 a_n7191_n9484.t4 305.683
R15493 a_n7191_n9484.n2 a_n7191_n9484.n0 16.879
R15494 a_n7191_n9484.n3 a_n7191_n9484.n2 10.8867
R15495 a_n7191_n9484.n2 a_n7191_n9484.n1 9.3005
R15496 a_8575_3923.t0 a_8575_3923.n0 1327.82
R15497 a_8575_3923.n0 a_8575_3923.t1 194.655
R15498 a_8575_3923.n0 a_8575_3923.t2 63.3219
R15499 auto_sampling_0.x14.D.n5 auto_sampling_0.x14.D.n4 585
R15500 auto_sampling_0.x14.D.n4 auto_sampling_0.x14.D.n3 585
R15501 auto_sampling_0.x14.D.n2 auto_sampling_0.x14.D.t4 333.651
R15502 auto_sampling_0.x14.D.n2 auto_sampling_0.x14.D.t5 297.233
R15503 auto_sampling_0.x14.D auto_sampling_0.x14.D.n2 196.493
R15504 auto_sampling_0.x14.D.n1 auto_sampling_0.x14.D.n0 185
R15505 auto_sampling_0.x14.D auto_sampling_0.x14.D.n1 49.0339
R15506 auto_sampling_0.x14.D.n3 auto_sampling_0.x14.D 44.2533
R15507 auto_sampling_0.x14.D.n4 auto_sampling_0.x14.D.t2 26.5955
R15508 auto_sampling_0.x14.D.n4 auto_sampling_0.x14.D.t3 26.5955
R15509 auto_sampling_0.x14.D.n0 auto_sampling_0.x14.D.t0 24.9236
R15510 auto_sampling_0.x14.D.n0 auto_sampling_0.x14.D.t1 24.9236
R15511 auto_sampling_0.x14.D.n5 auto_sampling_0.x14.D 15.6165
R15512 auto_sampling_0.x14.D.n1 auto_sampling_0.x14.D 10.4965
R15513 auto_sampling_0.x14.D.n3 auto_sampling_0.x14.D 1.7925
R15514 auto_sampling_0.x14.D auto_sampling_0.x14.D.n5 1.7925
R15515 a_2575_2717.n1 a_2575_2717.n0 926.024
R15516 a_2575_2717.t0 a_2575_2717.n1 82.0838
R15517 a_2575_2717.n0 a_2575_2717.t3 63.3338
R15518 a_2575_2717.n1 a_2575_2717.t2 63.3219
R15519 a_2575_2717.n0 a_2575_2717.t1 29.7268
R15520 a_792_n9484.n1 a_792_n9484.n0 926.024
R15521 a_792_n9484.t1 a_792_n9484.n1 82.0838
R15522 a_792_n9484.n0 a_792_n9484.t0 63.3338
R15523 a_792_n9484.n1 a_792_n9484.t3 63.3219
R15524 a_792_n9484.n0 a_792_n9484.t2 29.7268
R15525 a_9342_n9118.t0 a_9342_n9118.t1 126.644
R15526 a_2289_n1029.t1 a_2289_n1029.n3 370.026
R15527 a_2289_n1029.n0 a_2289_n1029.t4 351.356
R15528 a_2289_n1029.n1 a_2289_n1029.t3 334.717
R15529 a_2289_n1029.n3 a_2289_n1029.t0 325.971
R15530 a_2289_n1029.n1 a_2289_n1029.t2 309.935
R15531 a_2289_n1029.n0 a_2289_n1029.t5 305.683
R15532 a_2289_n1029.n2 a_2289_n1029.n0 16.879
R15533 a_2289_n1029.n3 a_2289_n1029.n2 10.8867
R15534 a_2289_n1029.n2 a_2289_n1029.n1 9.3005
R15535 a_n274_3557.t0 a_n274_3557.t1 87.1434
R15536 a_4656_n9484.n1 a_4656_n9484.n0 926.024
R15537 a_4656_n9484.t1 a_4656_n9484.n1 82.0838
R15538 a_4656_n9484.n0 a_4656_n9484.t0 63.3338
R15539 a_4656_n9484.n1 a_4656_n9484.t3 63.3219
R15540 a_4656_n9484.n0 a_4656_n9484.t2 29.7268
R15541 a_1303_2717.n3 a_1303_2717.n2 636.953
R15542 a_1303_2717.n1 a_1303_2717.t5 366.856
R15543 a_1303_2717.n2 a_1303_2717.n0 300.2
R15544 a_1303_2717.n2 a_1303_2717.n1 225.036
R15545 a_1303_2717.n1 a_1303_2717.t4 174.056
R15546 a_1303_2717.n0 a_1303_2717.t1 70.0005
R15547 a_1303_2717.n3 a_1303_2717.t2 68.0124
R15548 a_1303_2717.t0 a_1303_2717.n3 63.3219
R15549 a_1303_2717.n0 a_1303_2717.t3 61.6672
R15550 a_1478_2691.n5 a_1478_2691.n4 807.871
R15551 a_1478_2691.n2 a_1478_2691.t6 389.183
R15552 a_1478_2691.n3 a_1478_2691.n2 251.167
R15553 a_1478_2691.n3 a_1478_2691.t1 223.571
R15554 a_1478_2691.n0 a_1478_2691.t3 212.081
R15555 a_1478_2691.n1 a_1478_2691.t4 212.081
R15556 a_1478_2691.n4 a_1478_2691.n1 176.576
R15557 a_1478_2691.n2 a_1478_2691.t8 174.891
R15558 a_1478_2691.n0 a_1478_2691.t5 139.78
R15559 a_1478_2691.n1 a_1478_2691.t7 139.78
R15560 a_1478_2691.n5 a_1478_2691.t2 63.3219
R15561 a_1478_2691.t0 a_1478_2691.n5 63.3219
R15562 a_1478_2691.n1 a_1478_2691.n0 61.346
R15563 a_1478_2691.n4 a_1478_2691.n3 37.7195
R15564 a_5329_3083.t0 a_5329_3083.t1 126.644
R15565 a_n5259_n10022.t1 a_n5259_n10022.n3 370.026
R15566 a_n5259_n10022.n0 a_n5259_n10022.t2 351.356
R15567 a_n5259_n10022.n1 a_n5259_n10022.t4 334.717
R15568 a_n5259_n10022.n3 a_n5259_n10022.t0 325.971
R15569 a_n5259_n10022.n1 a_n5259_n10022.t3 309.935
R15570 a_n5259_n10022.n0 a_n5259_n10022.t5 305.683
R15571 a_n5259_n10022.n2 a_n5259_n10022.n0 16.879
R15572 a_n5259_n10022.n3 a_n5259_n10022.n2 10.8867
R15573 a_n5259_n10022.n2 a_n5259_n10022.n1 9.3005
R15574 a_4366_n5106.n3 a_4366_n5106.n2 647.119
R15575 a_4366_n5106.n1 a_4366_n5106.t5 350.253
R15576 a_4366_n5106.n2 a_4366_n5106.n0 260.339
R15577 a_4366_n5106.n2 a_4366_n5106.n1 246.119
R15578 a_4366_n5106.n1 a_4366_n5106.t4 189.588
R15579 a_4366_n5106.n3 a_4366_n5106.t0 89.1195
R15580 a_4366_n5106.n0 a_4366_n5106.t3 63.3338
R15581 a_4366_n5106.t2 a_4366_n5106.n3 41.0422
R15582 a_4366_n5106.n0 a_4366_n5106.t1 31.9797
R15583 a_n1395_n9484.t1 a_n1395_n9484.n3 370.026
R15584 a_n1395_n9484.n0 a_n1395_n9484.t2 351.356
R15585 a_n1395_n9484.n1 a_n1395_n9484.t4 334.717
R15586 a_n1395_n9484.n3 a_n1395_n9484.t0 325.971
R15587 a_n1395_n9484.n1 a_n1395_n9484.t5 309.935
R15588 a_n1395_n9484.n0 a_n1395_n9484.t3 305.683
R15589 a_n1395_n9484.n2 a_n1395_n9484.n0 16.879
R15590 a_n1395_n9484.n3 a_n1395_n9484.n2 10.8867
R15591 a_n1395_n9484.n2 a_n1395_n9484.n1 9.3005
R15592 a_8118_n5624.n0 a_8118_n5624.t1 68.3338
R15593 a_8118_n5624.n0 a_8118_n5624.t0 26.3935
R15594 a_8118_n5624.n1 a_8118_n5624.n0 14.4005
R15595 a_2747_n663.n0 a_2747_n663.t2 1327.82
R15596 a_2747_n663.t0 a_2747_n663.n0 194.655
R15597 a_2747_n663.n0 a_2747_n663.t1 63.3219
R15598 a_1561_n9484.t1 a_1561_n9484.t0 94.7268
R15599 a_4789_n787.n3 a_4789_n787.n2 647.119
R15600 a_4789_n787.n1 a_4789_n787.t5 350.253
R15601 a_4789_n787.n2 a_4789_n787.n0 260.339
R15602 a_4789_n787.n2 a_4789_n787.n1 246.119
R15603 a_4789_n787.n1 a_4789_n787.t4 189.588
R15604 a_4789_n787.n3 a_4789_n787.t1 89.1195
R15605 a_4789_n787.n0 a_4789_n787.t0 63.3338
R15606 a_4789_n787.t3 a_4789_n787.n3 41.0422
R15607 a_4789_n787.n0 a_4789_n787.t2 31.9797
R15608 a_5316_n9484.n3 a_5316_n9484.n2 636.953
R15609 a_5316_n9484.n1 a_5316_n9484.t5 366.856
R15610 a_5316_n9484.n2 a_5316_n9484.n0 300.2
R15611 a_5316_n9484.n2 a_5316_n9484.n1 225.036
R15612 a_5316_n9484.n1 a_5316_n9484.t4 174.056
R15613 a_5316_n9484.n0 a_5316_n9484.t3 70.0005
R15614 a_5316_n9484.t1 a_5316_n9484.n3 68.0124
R15615 a_5316_n9484.n3 a_5316_n9484.t2 63.3219
R15616 a_5316_n9484.n0 a_5316_n9484.t0 61.6672
R15617 a_6342_n4714.t0 a_6342_n4714.t1 60.0005
R15618 SWN[2].n4 SWN[2].n3 585
R15619 SWN[2].n3 SWN[2].n2 585
R15620 SWN[2].n1 SWN[2].n0 185
R15621 SWN[2].n5 SWN[2].n1 53.3859
R15622 SWN[2].n3 SWN[2].t3 26.5955
R15623 SWN[2].n3 SWN[2].t2 26.5955
R15624 SWN[2].n0 SWN[2].t0 24.9236
R15625 SWN[2].n0 SWN[2].t1 24.9236
R15626 SWN[2] SWN[2].n5 14.6566
R15627 SWN[2] SWN[2].n4 10.4965
R15628 SWN[2].n2 SWN[2] 10.4965
R15629 SWN[2].n4 SWN[2] 6.9125
R15630 SWN[2].n2 SWN[2] 6.9125
R15631 SWN[2].n5 SWN[2] 4.3525
R15632 SWN[2].n1 SWN[2] 1.7925
R15633 a_6408_n1029.n1 a_6408_n1029.n0 926.024
R15634 a_6408_n1029.t1 a_6408_n1029.n1 82.0838
R15635 a_6408_n1029.n0 a_6408_n1029.t0 63.3338
R15636 a_6408_n1029.n1 a_6408_n1029.t3 63.3219
R15637 a_6408_n1029.n0 a_6408_n1029.t2 29.7268
R15638 SWN[4].n4 SWN[4].n3 585
R15639 SWN[4].n3 SWN[4].n2 585
R15640 SWN[4].n1 SWN[4].n0 185
R15641 SWN[4].n5 SWN[4].n1 53.3859
R15642 SWN[4].n3 SWN[4].t2 26.5955
R15643 SWN[4].n3 SWN[4].t3 26.5955
R15644 SWN[4].n0 SWN[4].t0 24.9236
R15645 SWN[4].n0 SWN[4].t1 24.9236
R15646 SWN[4] SWN[4].n5 14.676
R15647 SWN[4] SWN[4].n4 10.4965
R15648 SWN[4].n2 SWN[4] 10.4965
R15649 SWN[4].n4 SWN[4] 6.9125
R15650 SWN[4].n2 SWN[4] 6.9125
R15651 SWN[4].n5 SWN[4] 4.3525
R15652 SWN[4].n1 SWN[4] 1.7925
R15653 a_n6276_n9484.n3 a_n6276_n9484.n2 636.953
R15654 a_n6276_n9484.n1 a_n6276_n9484.t4 366.856
R15655 a_n6276_n9484.n2 a_n6276_n9484.n0 300.2
R15656 a_n6276_n9484.n2 a_n6276_n9484.n1 225.036
R15657 a_n6276_n9484.n1 a_n6276_n9484.t5 174.056
R15658 a_n6276_n9484.n0 a_n6276_n9484.t3 70.0005
R15659 a_n6276_n9484.t1 a_n6276_n9484.n3 68.0124
R15660 a_n6276_n9484.n3 a_n6276_n9484.t2 63.3219
R15661 a_n6276_n9484.n0 a_n6276_n9484.t0 61.6672
R15662 a_223_3557.n1 a_223_3557.t7 530.01
R15663 a_223_3557.t1 a_223_3557.n5 421.021
R15664 a_223_3557.n0 a_223_3557.t4 337.142
R15665 a_223_3557.n3 a_223_3557.t0 280.223
R15666 a_223_3557.n4 a_223_3557.t2 263.173
R15667 a_223_3557.n4 a_223_3557.t3 227.826
R15668 a_223_3557.n0 a_223_3557.t5 199.762
R15669 a_223_3557.n2 a_223_3557.n1 170.81
R15670 a_223_3557.n2 a_223_3557.n0 167.321
R15671 a_223_3557.n5 a_223_3557.n4 152
R15672 a_223_3557.n1 a_223_3557.t6 141.923
R15673 a_223_3557.n3 a_223_3557.n2 10.8376
R15674 a_223_3557.n5 a_223_3557.n3 2.50485
R15675 a_898_n5624.t1 a_898_n5624.t0 198.571
R15676 CF[0].n17 CF[0].n16 585
R15677 CF[0].n18 CF[0].n17 585
R15678 CF[0].n3 CF[0].t7 294.557
R15679 CF[0].n0 CF[0].t6 294.557
R15680 CF[0].n6 CF[0].t8 235.763
R15681 CF[0].n10 CF[0].t13 221.72
R15682 CF[0].n7 CF[0].t9 221.72
R15683 CF[0].n3 CF[0].t12 211.01
R15684 CF[0].n0 CF[0].t10 211.01
R15685 CF[0].n15 CF[0].n14 185
R15686 CF[0].n6 CF[0].t4 163.464
R15687 CF[0].n4 CF[0].n3 153.097
R15688 CF[0].n9 CF[0].n8 152
R15689 CF[0].n12 CF[0].n11 152
R15690 CF[0].n13 CF[0].n6 152
R15691 CF[0].n1 CF[0].n0 152
R15692 CF[0].n10 CF[0].t11 149.421
R15693 CF[0].n7 CF[0].t5 149.421
R15694 CF[0] CF[0].n21 71.8051
R15695 CF[0].n9 CF[0].n7 58.019
R15696 CF[0] CF[0].n15 57.7379
R15697 CF[0].n11 CF[0].n10 43.7375
R15698 CF[0].n21 CF[0] 36.914
R15699 CF[0].n17 CF[0].t2 26.5955
R15700 CF[0].n17 CF[0].t3 26.5955
R15701 CF[0].n14 CF[0].t0 24.9236
R15702 CF[0].n14 CF[0].t1 24.9236
R15703 CF[0] CF[0].n12 20.8005
R15704 CF[0].n11 CF[0].n6 17.8524
R15705 CF[0].n10 CF[0].n9 16.9598
R15706 CF[0].n8 CF[0] 16.3205
R15707 CF[0].n5 CF[0].n2 14.9321
R15708 CF[0].n20 CF[0].n13 14.5044
R15709 CF[0].n5 CF[0].n4 13.9063
R15710 CF[0].n20 CF[0].n19 13.8005
R15711 CF[0].n8 CF[0] 13.1205
R15712 CF[0].n16 CF[0] 10.4965
R15713 CF[0].n18 CF[0] 10.4965
R15714 CF[0].n2 CF[0] 9.32621
R15715 CF[0].n21 CF[0] 8.71425
R15716 CF[0].n12 CF[0] 8.6405
R15717 CF[0].n16 CF[0] 6.9125
R15718 CF[0].n19 CF[0] 4.3525
R15719 CF[0].n4 CF[0] 3.10907
R15720 CF[0].n19 CF[0].n18 2.5605
R15721 CF[0].n1 CF[0] 2.01193
R15722 CF[0].n15 CF[0] 1.7925
R15723 CF[0].n2 CF[0].n1 1.09764
R15724 CF[0].n13 CF[0] 0.9605
R15725 CF[0] CF[0].n20 0.923018
R15726 CF[0] CF[0].n5 0.856103
R15727 a_8301_n1207.t0 a_8301_n1207.t1 87.1434
R15728 a_9140_2717.t0 a_9140_2717.t1 94.7268
R15729 a_2779_3923.t0 a_2779_3923.n0 1327.82
R15730 a_2779_3923.n0 a_2779_3923.t1 194.655
R15731 a_2779_3923.n0 a_2779_3923.t2 63.3219
R15732 a_8461_n5258.t0 a_8461_n5258.n0 1327.82
R15733 a_8461_n5258.n0 a_8461_n5258.t2 194.655
R15734 a_8461_n5258.n0 a_8461_n5258.t1 63.3219
R15735 a_8316_n5387.n3 a_8316_n5387.n2 674.338
R15736 a_8316_n5387.n1 a_8316_n5387.t5 332.58
R15737 a_8316_n5387.n2 a_8316_n5387.n0 284.012
R15738 a_8316_n5387.n2 a_8316_n5387.n1 253.648
R15739 a_8316_n5387.n1 a_8316_n5387.t4 168.701
R15740 a_8316_n5387.n3 a_8316_n5387.t3 96.1553
R15741 a_8316_n5387.t1 a_8316_n5387.n3 65.6672
R15742 a_8316_n5387.n0 a_8316_n5387.t2 65.0005
R15743 a_8316_n5387.n0 a_8316_n5387.t0 45.0005
R15744 a_n8677_n9650.t1 a_n8677_n9650.t0 198.571
R15745 a_n8511_n9662.t0 a_n8511_n9662.t1 60.0005
R15746 SWP[3].n0 SWP[3].t4 333.651
R15747 SWP[3].n0 SWP[3].t5 297.233
R15748 SWP[3].n4 SWP[3].n3 289.096
R15749 SWP[3].n1 SWP[3].n0 196.493
R15750 SWP[3].n6 SWP[3].n5 185
R15751 SWP[3] SWP[3].n6 49.0339
R15752 SWP[3].n2 SWP[3] 47.3888
R15753 SWP[3] SWP[3].n1 39.5082
R15754 SWP[3].n3 SWP[3].t2 26.5955
R15755 SWP[3].n3 SWP[3].t3 26.5955
R15756 SWP[3].n5 SWP[3].t0 24.9236
R15757 SWP[3].n5 SWP[3].t1 24.9236
R15758 SWP[3] SWP[3].n7 14.6049
R15759 SWP[3] SWP[3].n2 14.3123
R15760 SWP[3].n7 SWP[3] 13.0565
R15761 SWP[3].n2 SWP[3] 12.0667
R15762 SWP[3].n6 SWP[3] 10.4965
R15763 SWP[3] SWP[3].n4 9.48653
R15764 SWP[3].n4 SWP[3] 7.7181
R15765 SWP[3].n7 SWP[3] 4.3525
R15766 SWP[3].n1 SWP[3] 0.24431
R15767 a_8274_n4714.t0 a_8274_n4714.t1 60.0005
R15768 a_538_n1441.n3 a_538_n1441.n2 636.953
R15769 a_538_n1441.n1 a_538_n1441.t4 366.856
R15770 a_538_n1441.n2 a_538_n1441.n0 300.2
R15771 a_538_n1441.n2 a_538_n1441.n1 225.036
R15772 a_538_n1441.n1 a_538_n1441.t5 174.056
R15773 a_538_n1441.n0 a_538_n1441.t1 70.0005
R15774 a_538_n1441.n3 a_538_n1441.t3 68.0124
R15775 a_538_n1441.t0 a_538_n1441.n3 63.3219
R15776 a_538_n1441.n0 a_538_n1441.t2 61.6672
R15777 a_4847_n9484.t1 a_4847_n9484.t0 198.571
R15778 a_4213_n5258.t0 a_4213_n5258.t1 126.644
R15779 a_2748_n1457.t1 a_2748_n1457.n3 370.026
R15780 a_2748_n1457.n0 a_2748_n1457.t3 351.356
R15781 a_2748_n1457.n1 a_2748_n1457.t4 334.717
R15782 a_2748_n1457.n3 a_2748_n1457.t0 325.971
R15783 a_2748_n1457.n1 a_2748_n1457.t2 309.935
R15784 a_2748_n1457.n0 a_2748_n1457.t5 305.683
R15785 a_2748_n1457.n2 a_2748_n1457.n0 16.879
R15786 a_2748_n1457.n3 a_2748_n1457.n2 10.8867
R15787 a_2748_n1457.n2 a_2748_n1457.n1 9.3005
R15788 a_3506_n1573.n1 a_3506_n1573.n0 926.024
R15789 a_3506_n1573.n0 a_3506_n1573.t3 82.0838
R15790 a_3506_n1573.n1 a_3506_n1573.t0 63.3338
R15791 a_3506_n1573.n0 a_3506_n1573.t2 63.3219
R15792 a_3506_n1573.n2 a_3506_n1573.t1 26.3935
R15793 a_3506_n1573.n3 a_3506_n1573.n2 14.4005
R15794 a_3506_n1573.n2 a_3506_n1573.n1 3.33383
R15795 a_8563_3557.t1 a_8563_3557.t0 198.571
R15796 a_8729_3557.t0 a_8729_3557.t1 60.0005
R15797 a_3037_n9242.n3 a_3037_n9242.n2 647.119
R15798 a_3037_n9242.n1 a_3037_n9242.t5 350.253
R15799 a_3037_n9242.n2 a_3037_n9242.n0 260.339
R15800 a_3037_n9242.n2 a_3037_n9242.n1 246.119
R15801 a_3037_n9242.n1 a_3037_n9242.t4 189.588
R15802 a_3037_n9242.n3 a_3037_n9242.t3 89.1195
R15803 a_3037_n9242.n0 a_3037_n9242.t2 63.3338
R15804 a_3037_n9242.t1 a_3037_n9242.n3 41.0422
R15805 a_3037_n9242.n0 a_3037_n9242.t0 31.9797
R15806 a_3493_n9650.n0 a_3493_n9650.t1 68.3338
R15807 a_3493_n9650.n0 a_3493_n9650.t0 26.3935
R15808 a_3493_n9650.n1 a_3493_n9650.n0 14.4005
R15809 a_2303_n10022.n1 a_2303_n10022.t5 530.01
R15810 a_2303_n10022.t1 a_2303_n10022.n5 421.021
R15811 a_2303_n10022.n0 a_2303_n10022.t3 337.142
R15812 a_2303_n10022.n3 a_2303_n10022.t0 280.223
R15813 a_2303_n10022.n4 a_2303_n10022.t7 263.173
R15814 a_2303_n10022.n4 a_2303_n10022.t6 227.826
R15815 a_2303_n10022.n0 a_2303_n10022.t2 199.762
R15816 a_2303_n10022.n2 a_2303_n10022.n1 170.81
R15817 a_2303_n10022.n2 a_2303_n10022.n0 167.321
R15818 a_2303_n10022.n5 a_2303_n10022.n4 152
R15819 a_2303_n10022.n1 a_2303_n10022.t4 141.923
R15820 a_2303_n10022.n3 a_2303_n10022.n2 10.8376
R15821 a_2303_n10022.n5 a_2303_n10022.n3 2.50485
R15822 a_5491_n9724.n5 a_5491_n9724.n4 807.871
R15823 a_5491_n9724.n2 a_5491_n9724.t3 389.183
R15824 a_5491_n9724.n3 a_5491_n9724.n2 251.167
R15825 a_5491_n9724.n3 a_5491_n9724.t1 223.571
R15826 a_5491_n9724.n0 a_5491_n9724.t4 212.081
R15827 a_5491_n9724.n1 a_5491_n9724.t5 212.081
R15828 a_5491_n9724.n4 a_5491_n9724.n1 176.576
R15829 a_5491_n9724.n2 a_5491_n9724.t6 174.891
R15830 a_5491_n9724.n0 a_5491_n9724.t7 139.78
R15831 a_5491_n9724.n1 a_5491_n9724.t8 139.78
R15832 a_5491_n9724.t0 a_5491_n9724.n5 63.3219
R15833 a_5491_n9724.n5 a_5491_n9724.t2 63.3219
R15834 a_5491_n9724.n1 a_5491_n9724.n0 61.346
R15835 a_5491_n9724.n4 a_5491_n9724.n3 37.7195
R15836 a_5478_n10028.t0 a_5478_n10028.t1 126.644
R15837 a_957_3799.n3 a_957_3799.n2 647.119
R15838 a_957_3799.n1 a_957_3799.t4 350.253
R15839 a_957_3799.n2 a_957_3799.n0 260.339
R15840 a_957_3799.n2 a_957_3799.n1 246.119
R15841 a_957_3799.n1 a_957_3799.t5 189.588
R15842 a_957_3799.n3 a_957_3799.t2 89.1195
R15843 a_957_3799.n0 a_957_3799.t3 63.3338
R15844 a_957_3799.t0 a_957_3799.n3 41.0422
R15845 a_957_3799.n0 a_957_3799.t1 31.9797
R15846 a_835_3557.t0 a_835_3557.t1 198.571
R15847 a_1001_3557.t0 a_1001_3557.t1 60.0005
R15848 a_n8046_n10028.t0 a_n8046_n10028.t1 126.644
R15849 a_n1140_n9484.n1 a_n1140_n9484.n0 926.024
R15850 a_n1140_n9484.n0 a_n1140_n9484.t3 82.0838
R15851 a_n1140_n9484.n1 a_n1140_n9484.t0 63.3338
R15852 a_n1140_n9484.n0 a_n1140_n9484.t2 63.3219
R15853 a_n1140_n9484.n2 a_n1140_n9484.t1 26.3935
R15854 a_n1140_n9484.n3 a_n1140_n9484.n2 14.4005
R15855 a_n1140_n9484.n2 a_n1140_n9484.n1 3.33383
R15856 a_803_n1029.t0 a_803_n1029.t1 198.571
R15857 a_969_n1029.t0 a_969_n1029.t1 60.0005
R15858 a_9193_3083.t0 a_9193_3083.t1 126.644
R15859 a_n5425_n9484.n1 a_n5425_n9484.t3 530.01
R15860 a_n5425_n9484.t1 a_n5425_n9484.n5 421.021
R15861 a_n5425_n9484.n0 a_n5425_n9484.t2 337.142
R15862 a_n5425_n9484.n3 a_n5425_n9484.t0 280.223
R15863 a_n5425_n9484.n4 a_n5425_n9484.t6 263.173
R15864 a_n5425_n9484.n4 a_n5425_n9484.t7 227.826
R15865 a_n5425_n9484.n0 a_n5425_n9484.t5 199.762
R15866 a_n5425_n9484.n2 a_n5425_n9484.n1 170.81
R15867 a_n5425_n9484.n2 a_n5425_n9484.n0 167.321
R15868 a_n5425_n9484.n5 a_n5425_n9484.n4 152
R15869 a_n5425_n9484.n1 a_n5425_n9484.t4 141.923
R15870 a_n5425_n9484.n3 a_n5425_n9484.n2 10.8376
R15871 a_n5425_n9484.n5 a_n5425_n9484.n3 2.50485
R15872 SWP[2].n0 SWP[2].t4 332.312
R15873 SWP[2].n0 SWP[2].t5 295.627
R15874 SWP[2].n3 SWP[2].n2 289.096
R15875 SWP[2] SWP[2].n0 196.004
R15876 SWP[2].n5 SWP[2].n4 185
R15877 SWP[2] SWP[2].n5 49.0339
R15878 SWP[2].n1 SWP[2] 44.6416
R15879 SWP[2].n2 SWP[2].t2 26.5955
R15880 SWP[2].n2 SWP[2].t3 26.5955
R15881 SWP[2].n4 SWP[2].t0 24.9236
R15882 SWP[2].n4 SWP[2].t1 24.9236
R15883 SWP[2] SWP[2].n1 21.6493
R15884 SWP[2] SWP[2].n6 14.6092
R15885 SWP[2].n6 SWP[2] 13.0565
R15886 SWP[2].n1 SWP[2] 11.7357
R15887 SWP[2].n5 SWP[2] 10.4965
R15888 SWP[2] SWP[2].n3 9.48653
R15889 SWP[2].n3 SWP[2] 7.7181
R15890 SWP[2].n6 SWP[2] 4.3525
R15891 a_n1086_3083.t0 a_n1086_3083.n0 1327.82
R15892 a_n1086_3083.n0 a_n1086_3083.t1 194.655
R15893 a_n1086_3083.n0 a_n1086_3083.t2 63.3219
R15894 a_n519_3557.t1 a_n519_3557.t0 94.7268
R15895 a_3738_n9484.t0 a_3738_n9484.t1 87.1434
R15896 a_n4235_n9650.n0 a_n4235_n9650.t1 68.3338
R15897 a_n4235_n9650.n0 a_n4235_n9650.t0 26.3935
R15898 a_n4235_n9650.n1 a_n4235_n9650.n0 14.4005
R15899 a_2735_n1029.t1 a_2735_n1029.t0 198.571
R15900 a_7261_3083.t0 a_7261_3083.t1 126.644
R15901 a_5277_3557.t1 a_5277_3557.t0 94.7268
R15902 a_n1140_n9662.n1 a_n1140_n9662.n0 926.024
R15903 a_n1140_n9662.t0 a_n1140_n9662.n1 82.0838
R15904 a_n1140_n9662.n0 a_n1140_n9662.t1 63.3338
R15905 a_n1140_n9662.n1 a_n1140_n9662.t3 63.3219
R15906 a_n1140_n9662.n0 a_n1140_n9662.t2 29.7268
R15907 a_8884_n1573.n0 a_8884_n1573.t2 1327.82
R15908 a_8884_n1573.t0 a_8884_n1573.n0 194.655
R15909 a_8884_n1573.n0 a_8884_n1573.t1 63.3219
R15910 a_n371_n9650.n0 a_n371_n9650.t0 68.3338
R15911 a_n371_n9650.n0 a_n371_n9650.t1 26.3935
R15912 a_n371_n9650.n1 a_n371_n9650.n0 14.4005
R15913 a_7248_n9484.n3 a_7248_n9484.n2 636.953
R15914 a_7248_n9484.n1 a_7248_n9484.t4 366.856
R15915 a_7248_n9484.n2 a_7248_n9484.n0 300.2
R15916 a_7248_n9484.n2 a_7248_n9484.n1 225.036
R15917 a_7248_n9484.n1 a_7248_n9484.t5 174.056
R15918 a_7248_n9484.n0 a_7248_n9484.t2 70.0005
R15919 a_7248_n9484.t1 a_7248_n9484.n3 68.0124
R15920 a_7248_n9484.n3 a_7248_n9484.t3 63.3219
R15921 a_7248_n9484.n0 a_7248_n9484.t0 61.6672
R15922 a_7410_n9118.t0 a_7410_n9118.t1 126.644
R15923 a_2767_3557.t0 a_2767_3557.t1 198.571
R15924 a_2933_3557.t0 a_2933_3557.t1 60.0005
R15925 a_4859_n9118.n0 a_4859_n9118.t1 1327.82
R15926 a_4859_n9118.t0 a_4859_n9118.n0 194.655
R15927 a_4859_n9118.n0 a_4859_n9118.t2 63.3219
R15928 a_9342_n10028.t0 a_9342_n10028.t1 126.644
R15929 a_2576_3557.n1 a_2576_3557.n0 926.024
R15930 a_2576_3557.n0 a_2576_3557.t3 82.0838
R15931 a_2576_3557.n1 a_2576_3557.t0 63.3338
R15932 a_2576_3557.n0 a_2576_3557.t2 63.3219
R15933 a_2576_3557.n2 a_2576_3557.t1 26.3935
R15934 a_2576_3557.n3 a_2576_3557.n2 14.4005
R15935 a_2576_3557.n2 a_2576_3557.n1 3.33383
R15936 a_6642_3083.t0 a_6642_3083.n0 1327.82
R15937 a_6642_3083.n0 a_6642_3083.t1 194.655
R15938 a_6642_3083.n0 a_6642_3083.t2 63.3219
R15939 a_n6167_n9484.t1 a_n6167_n9484.t0 94.7268
R15940 a_7423_n9724.n5 a_7423_n9724.n4 807.871
R15941 a_7423_n9724.n2 a_7423_n9724.t8 389.183
R15942 a_7423_n9724.n3 a_7423_n9724.n2 251.167
R15943 a_7423_n9724.n3 a_7423_n9724.t1 223.571
R15944 a_7423_n9724.n0 a_7423_n9724.t6 212.081
R15945 a_7423_n9724.n1 a_7423_n9724.t4 212.081
R15946 a_7423_n9724.n4 a_7423_n9724.n1 176.576
R15947 a_7423_n9724.n2 a_7423_n9724.t7 174.891
R15948 a_7423_n9724.n0 a_7423_n9724.t5 139.78
R15949 a_7423_n9724.n1 a_7423_n9724.t3 139.78
R15950 a_7423_n9724.t0 a_7423_n9724.n5 63.3219
R15951 a_7423_n9724.n5 a_7423_n9724.t2 63.3219
R15952 a_7423_n9724.n1 a_7423_n9724.n0 61.346
R15953 a_7423_n9724.n4 a_7423_n9724.n3 37.7195
R15954 a_5136_n1029.n3 a_5136_n1029.n2 636.953
R15955 a_5136_n1029.n1 a_5136_n1029.t5 366.856
R15956 a_5136_n1029.n2 a_5136_n1029.n0 300.2
R15957 a_5136_n1029.n2 a_5136_n1029.n1 225.036
R15958 a_5136_n1029.n1 a_5136_n1029.t4 174.056
R15959 a_5136_n1029.n0 a_5136_n1029.t1 70.0005
R15960 a_5136_n1029.n3 a_5136_n1029.t2 68.0124
R15961 a_5136_n1029.t0 a_5136_n1029.n3 63.3219
R15962 a_5136_n1029.n0 a_5136_n1029.t3 61.6672
R15963 a_5438_n1573.n1 a_5438_n1573.n0 926.024
R15964 a_5438_n1573.t1 a_5438_n1573.n1 82.0838
R15965 a_5438_n1573.n0 a_5438_n1573.t0 63.3338
R15966 a_5438_n1573.n1 a_5438_n1573.t3 63.3219
R15967 a_5438_n1573.n0 a_5438_n1573.t2 29.7268
R15968 a_7602_n9484.t0 a_7602_n9484.t1 87.1434
R15969 a_7423_n9510.n5 a_7423_n9510.n4 807.871
R15970 a_7423_n9510.n2 a_7423_n9510.t5 389.183
R15971 a_7423_n9510.n3 a_7423_n9510.n2 251.167
R15972 a_7423_n9510.n3 a_7423_n9510.t1 223.571
R15973 a_7423_n9510.n0 a_7423_n9510.t8 212.081
R15974 a_7423_n9510.n1 a_7423_n9510.t6 212.081
R15975 a_7423_n9510.n4 a_7423_n9510.n1 176.576
R15976 a_7423_n9510.n2 a_7423_n9510.t3 174.891
R15977 a_7423_n9510.n0 a_7423_n9510.t7 139.78
R15978 a_7423_n9510.n1 a_7423_n9510.t4 139.78
R15979 a_7423_n9510.t0 a_7423_n9510.n5 63.3219
R15980 a_7423_n9510.n5 a_7423_n9510.t2 63.3219
R15981 a_7423_n9510.n1 a_7423_n9510.n0 61.346
R15982 a_7423_n9510.n4 a_7423_n9510.n3 37.7195
R15983 a_1465_3083.t0 a_1465_3083.t1 126.644
R15984 a_n827_n9242.n3 a_n827_n9242.n2 647.119
R15985 a_n827_n9242.n1 a_n827_n9242.t5 350.253
R15986 a_n827_n9242.n2 a_n827_n9242.n0 260.339
R15987 a_n827_n9242.n2 a_n827_n9242.n1 246.119
R15988 a_n827_n9242.n1 a_n827_n9242.t4 189.588
R15989 a_n827_n9242.n3 a_n827_n9242.t2 89.1195
R15990 a_n827_n9242.n0 a_n827_n9242.t3 63.3338
R15991 a_n827_n9242.t1 a_n827_n9242.n3 41.0422
R15992 a_n827_n9242.n0 a_n827_n9242.t0 31.9797
R15993 a_7979_n1599.n4 a_7979_n1599.n1 807.871
R15994 a_7979_n1599.n0 a_7979_n1599.t8 389.183
R15995 a_7979_n1599.n5 a_7979_n1599.n0 251.167
R15996 a_7979_n1599.t0 a_7979_n1599.n5 223.571
R15997 a_7979_n1599.n3 a_7979_n1599.t6 212.081
R15998 a_7979_n1599.n2 a_7979_n1599.t7 212.081
R15999 a_7979_n1599.n4 a_7979_n1599.n3 176.576
R16000 a_7979_n1599.n0 a_7979_n1599.t5 174.891
R16001 a_7979_n1599.n3 a_7979_n1599.t3 139.78
R16002 a_7979_n1599.n2 a_7979_n1599.t4 139.78
R16003 a_7979_n1599.n1 a_7979_n1599.t2 63.3219
R16004 a_7979_n1599.n1 a_7979_n1599.t1 63.3219
R16005 a_7979_n1599.n3 a_7979_n1599.n2 61.346
R16006 a_7979_n1599.n5 a_7979_n1599.n4 37.5061
R16007 a_n931_3557.t0 a_n931_3557.t1 60.0005
R16008 a_n6936_n9662.n1 a_n6936_n9662.n0 926.024
R16009 a_n6936_n9662.t0 a_n6936_n9662.n1 82.0838
R16010 a_n6936_n9662.n0 a_n6936_n9662.t3 63.3338
R16011 a_n6936_n9662.n1 a_n6936_n9662.t2 63.3219
R16012 a_n6936_n9662.n0 a_n6936_n9662.t1 29.7268
R16013 a_1156_n1573.n0 a_1156_n1573.t2 1327.82
R16014 a_1156_n1573.t0 a_1156_n1573.n0 194.655
R16015 a_1156_n1573.n0 a_1156_n1573.t1 63.3219
R16016 a_5168_3557.n3 a_5168_3557.n2 636.953
R16017 a_5168_3557.n1 a_5168_3557.t5 366.856
R16018 a_5168_3557.n2 a_5168_3557.n0 300.2
R16019 a_5168_3557.n2 a_5168_3557.n1 225.036
R16020 a_5168_3557.n1 a_5168_3557.t4 174.056
R16021 a_5168_3557.n0 a_5168_3557.t3 70.0005
R16022 a_5168_3557.t0 a_5168_3557.n3 68.0124
R16023 a_5168_3557.n3 a_5168_3557.t2 63.3219
R16024 a_5168_3557.n0 a_5168_3557.t1 61.6672
R16025 a_983_n9484.t1 a_983_n9484.t0 198.571
R16026 a_1149_n9484.t0 a_1149_n9484.t1 60.0005
R16027 COMP_P.n6 COMP_P.t3 235.763
R16028 COMP_P.n1 COMP_P.t1 221.72
R16029 COMP_P.n0 COMP_P.t5 221.72
R16030 COMP_P.n6 COMP_P.t2 163.464
R16031 COMP_P.n3 COMP_P.n2 152
R16032 COMP_P.n5 COMP_P.n4 152
R16033 COMP_P.n7 COMP_P.n6 152
R16034 COMP_P.n1 COMP_P.t0 149.421
R16035 COMP_P.n0 COMP_P.t4 149.421
R16036 COMP_P.n9 COMP_P 129.843
R16037 COMP_P.n2 COMP_P.n1 58.019
R16038 COMP_P.n5 COMP_P.n0 43.7375
R16039 COMP_P.n4 COMP_P.n3 21.7605
R16040 COMP_P.n7 COMP_P 19.5205
R16041 COMP_P.n6 COMP_P.n5 17.8524
R16042 COMP_P.n2 COMP_P.n0 16.9598
R16043 COMP_P.n9 COMP_P.n8 10.747
R16044 COMP_P.n3 COMP_P 5.4405
R16045 COMP_P.n8 COMP_P 5.4405
R16046 COMP_P.n8 COMP_P.n7 4.4805
R16047 COMP_P.n4 COMP_P 2.2405
R16048 COMP_P COMP_P.n9 0.0225588
R16049 a_8520_n9484.n1 a_8520_n9484.n0 926.024
R16050 a_8520_n9484.t0 a_8520_n9484.n1 82.0838
R16051 a_8520_n9484.n0 a_8520_n9484.t1 63.3338
R16052 a_8520_n9484.n1 a_8520_n9484.t3 63.3219
R16053 a_8520_n9484.n0 a_8520_n9484.t2 29.7268
R16054 a_8615_n9484.n3 a_8615_n9484.n2 674.338
R16055 a_8615_n9484.n1 a_8615_n9484.t5 332.58
R16056 a_8615_n9484.n2 a_8615_n9484.n0 284.012
R16057 a_8615_n9484.n2 a_8615_n9484.n1 253.648
R16058 a_8615_n9484.n1 a_8615_n9484.t4 168.701
R16059 a_8615_n9484.n3 a_8615_n9484.t3 96.1553
R16060 a_8615_n9484.t1 a_8615_n9484.n3 65.6672
R16061 a_8615_n9484.n0 a_8615_n9484.t2 65.0005
R16062 a_8615_n9484.n0 a_8615_n9484.t0 45.0005
R16063 a_2745_n1207.t1 a_2745_n1207.t0 94.7268
R16064 a_4507_2717.n1 a_4507_2717.n0 926.024
R16065 a_4507_2717.t1 a_4507_2717.n1 82.0838
R16066 a_4507_2717.n0 a_4507_2717.t0 63.3338
R16067 a_4507_2717.n1 a_4507_2717.t3 63.3219
R16068 a_4507_2717.n0 a_4507_2717.t2 29.7268
R16069 a_4602_2717.n3 a_4602_2717.n2 674.338
R16070 a_4602_2717.n1 a_4602_2717.t4 332.58
R16071 a_4602_2717.n2 a_4602_2717.n0 284.012
R16072 a_4602_2717.n2 a_4602_2717.n1 253.648
R16073 a_4602_2717.n1 a_4602_2717.t5 168.701
R16074 a_4602_2717.t1 a_4602_2717.n3 96.1553
R16075 a_4602_2717.n3 a_4602_2717.t2 65.6672
R16076 a_4602_2717.n0 a_4602_2717.t0 65.0005
R16077 a_4602_2717.n0 a_4602_2717.t3 45.0005
R16078 a_5425_n9484.t1 a_5425_n9484.t0 94.7268
R16079 a_739_3557.n3 a_739_3557.n2 674.338
R16080 a_739_3557.n1 a_739_3557.t4 332.58
R16081 a_739_3557.n2 a_739_3557.n0 284.012
R16082 a_739_3557.n2 a_739_3557.n1 253.648
R16083 a_739_3557.n1 a_739_3557.t5 168.701
R16084 a_739_3557.t0 a_739_3557.n3 96.1553
R16085 a_739_3557.n3 a_739_3557.t2 65.6672
R16086 a_739_3557.n0 a_739_3557.t1 65.0005
R16087 a_739_3557.n0 a_739_3557.t3 45.0005
R16088 a_6807_n5080.t0 a_6807_n5080.t1 126.644
R16089 a_9141_3557.t1 a_9141_3557.t0 94.7268
R16090 a_4751_n9650.n3 a_4751_n9650.n2 674.338
R16091 a_4751_n9650.n1 a_4751_n9650.t5 332.58
R16092 a_4751_n9650.n2 a_4751_n9650.n0 284.012
R16093 a_4751_n9650.n2 a_4751_n9650.n1 253.648
R16094 a_4751_n9650.n1 a_4751_n9650.t4 168.701
R16095 a_4751_n9650.t0 a_4751_n9650.n3 96.1553
R16096 a_4751_n9650.n3 a_4751_n9650.t2 65.6672
R16097 a_4751_n9650.n0 a_4751_n9650.t1 65.0005
R16098 a_4751_n9650.n0 a_4751_n9650.t3 45.0005
R16099 DOUT[7].n3 DOUT[7].n2 585
R16100 DOUT[7].n4 DOUT[7].n3 585
R16101 DOUT[7].n1 DOUT[7].n0 185
R16102 DOUT[7] DOUT[7].n1 57.7379
R16103 DOUT[7].n3 DOUT[7].t3 26.5955
R16104 DOUT[7].n3 DOUT[7].t2 26.5955
R16105 DOUT[7].n0 DOUT[7].t1 24.9236
R16106 DOUT[7].n0 DOUT[7].t0 24.9236
R16107 DOUT[7] DOUT[7].n5 17.8783
R16108 DOUT[7].n2 DOUT[7] 10.4965
R16109 DOUT[7].n4 DOUT[7] 10.4965
R16110 DOUT[7].n2 DOUT[7] 6.9125
R16111 DOUT[7].n5 DOUT[7] 4.3525
R16112 DOUT[7].n5 DOUT[7].n4 2.5605
R16113 DOUT[7].n1 DOUT[7] 1.7925
R16114 DOUT[4].n3 DOUT[4].n2 585
R16115 DOUT[4].n4 DOUT[4].n3 585
R16116 DOUT[4].n1 DOUT[4].n0 185
R16117 DOUT[4] DOUT[4].n1 49.0339
R16118 DOUT[4].n3 DOUT[4].t2 26.5955
R16119 DOUT[4].n3 DOUT[4].t3 26.5955
R16120 DOUT[4].n0 DOUT[4].t0 24.9236
R16121 DOUT[4].n0 DOUT[4].t1 24.9236
R16122 DOUT[4] DOUT[4].n4 20.4383
R16123 DOUT[4].n2 DOUT[4] 15.6165
R16124 DOUT[4].n1 DOUT[4] 10.4965
R16125 DOUT[4].n4 DOUT[4] 1.7925
R16126 DOUT[4].n2 DOUT[4] 1.7925
R16127 a_7878_n5624.t0 a_7878_n5624.t1 87.1434
R16128 a_4710_3083.t0 a_4710_3083.n0 1327.82
R16129 a_4710_3083.n0 a_4710_3083.t1 194.655
R16130 a_4710_3083.n0 a_4710_3083.t2 63.3219
R16131 a_2324_n5080.t0 a_2324_n5080.n0 1327.82
R16132 a_2324_n5080.n0 a_2324_n5080.t1 194.655
R16133 a_2324_n5080.n0 a_2324_n5080.t2 63.3219
R16134 a_813_n1207.t1 a_813_n1207.t0 94.7268
R16135 a_n4801_n10028.n0 a_n4801_n10028.t1 1327.82
R16136 a_n4801_n10028.n0 a_n4801_n10028.t2 194.655
R16137 a_n4801_n10028.t0 a_n4801_n10028.n0 63.3219
R16138 a_8670_n1573.n3 a_8670_n1573.n2 647.119
R16139 a_8670_n1573.n1 a_8670_n1573.t5 350.253
R16140 a_8670_n1573.n2 a_8670_n1573.n0 260.339
R16141 a_8670_n1573.n2 a_8670_n1573.n1 246.119
R16142 a_8670_n1573.n1 a_8670_n1573.t4 189.588
R16143 a_8670_n1573.n3 a_8670_n1573.t0 89.1195
R16144 a_8670_n1573.n0 a_8670_n1573.t1 63.3338
R16145 a_8670_n1573.t3 a_8670_n1573.n3 41.0422
R16146 a_8670_n1573.n0 a_8670_n1573.t2 31.9797
R16147 a_5490_n1029.t0 a_5490_n1029.t1 87.1434
R16148 a_8265_n9484.t1 a_8265_n9484.n3 370.026
R16149 a_8265_n9484.n0 a_8265_n9484.t5 351.356
R16150 a_8265_n9484.n1 a_8265_n9484.t3 334.717
R16151 a_8265_n9484.n3 a_8265_n9484.t0 325.971
R16152 a_8265_n9484.n1 a_8265_n9484.t4 309.935
R16153 a_8265_n9484.n0 a_8265_n9484.t2 305.683
R16154 a_8265_n9484.n2 a_8265_n9484.n0 16.879
R16155 a_8265_n9484.n3 a_8265_n9484.n2 10.8867
R16156 a_8265_n9484.n2 a_8265_n9484.n1 9.3005
R16157 a_9534_n9662.t0 a_9534_n9662.t1 87.1434
R16158 a_3366_n663.t0 a_3366_n663.t1 126.644
R16159 a_573_n1207.t0 a_573_n1207.t1 87.1434
R16160 a_n232_n5074.n1 a_n232_n5074.t5 530.01
R16161 a_n232_n5074.t1 a_n232_n5074.n5 421.021
R16162 a_n232_n5074.n0 a_n232_n5074.t4 337.142
R16163 a_n232_n5074.n3 a_n232_n5074.t0 280.223
R16164 a_n232_n5074.n4 a_n232_n5074.t3 263.173
R16165 a_n232_n5074.n4 a_n232_n5074.t2 227.826
R16166 a_n232_n5074.n0 a_n232_n5074.t6 199.762
R16167 a_n232_n5074.n2 a_n232_n5074.n1 170.81
R16168 a_n232_n5074.n2 a_n232_n5074.n0 167.321
R16169 a_n232_n5074.n5 a_n232_n5074.n4 152
R16170 a_n232_n5074.n1 a_n232_n5074.t7 141.923
R16171 a_n232_n5074.n3 a_n232_n5074.n2 10.8376
R16172 a_n232_n5074.n5 a_n232_n5074.n3 2.50485
R16173 a_4636_n1573.t0 a_4636_n1573.t1 126.644
R16174 a_4821_3799.n3 a_4821_3799.n2 647.119
R16175 a_4821_3799.n1 a_4821_3799.t5 350.253
R16176 a_4821_3799.n2 a_4821_3799.n0 260.339
R16177 a_4821_3799.n2 a_4821_3799.n1 246.119
R16178 a_4821_3799.n1 a_4821_3799.t4 189.588
R16179 a_4821_3799.n3 a_4821_3799.t0 89.1195
R16180 a_4821_3799.n0 a_4821_3799.t1 63.3338
R16181 a_4821_3799.t3 a_4821_3799.n3 41.0422
R16182 a_4821_3799.n0 a_4821_3799.t2 31.9797
R16183 a_n8046_n9118.t0 a_n8046_n9118.t1 126.644
R16184 a_6622_n5624.t0 a_6622_n5624.t1 60.0005
R16185 a_3204_n1029.n3 a_3204_n1029.n2 636.953
R16186 a_3204_n1029.n1 a_3204_n1029.t5 366.856
R16187 a_3204_n1029.n2 a_3204_n1029.n0 300.2
R16188 a_3204_n1029.n2 a_3204_n1029.n1 225.036
R16189 a_3204_n1029.n1 a_3204_n1029.t4 174.056
R16190 a_3204_n1029.n0 a_3204_n1029.t1 70.0005
R16191 a_3204_n1029.n3 a_3204_n1029.t3 68.0124
R16192 a_3204_n1029.t0 a_3204_n1029.n3 63.3219
R16193 a_3204_n1029.n0 a_3204_n1029.t2 61.6672
R16194 a_3313_n1029.t0 a_3313_n1029.t1 94.7268
R16195 a_n466_3923.t0 a_n466_3923.t1 126.644
R16196 a_4762_n5624.t1 a_4762_n5624.t0 198.571
R16197 a_3398_3923.t0 a_3398_3923.t1 126.644
R16198 a_6791_n10028.n0 a_6791_n10028.t2 1327.82
R16199 a_6791_n10028.t0 a_6791_n10028.n0 194.655
R16200 a_6791_n10028.n0 a_6791_n10028.t1 63.3219
R16201 a_1151_n5258.n1 a_1151_n5258.n0 926.024
R16202 a_1151_n5258.t1 a_1151_n5258.n1 82.0838
R16203 a_1151_n5258.n0 a_1151_n5258.t0 63.3338
R16204 a_1151_n5258.n1 a_1151_n5258.t3 63.3219
R16205 a_1151_n5258.n0 a_1151_n5258.t2 29.7268
R16206 CLKSB.n1 CLKSB.t1 233.815
R16207 CLKSB CLKSB.t0 152.889
R16208 CLKSB CLKSB.n1 14.5864
R16209 CLKSB.n0 CLKSB 2.22659
R16210 CLKSB.n1 CLKSB.n0 1.74595
R16211 CLKSB.n0 CLKSB 1.55202
R16212 SWN[8].n4 SWN[8].n3 585
R16213 SWN[8].n3 SWN[8].n2 585
R16214 SWN[8].n1 SWN[8].n0 185
R16215 SWN[8].n5 SWN[8].n1 53.3859
R16216 SWN[8].n3 SWN[8].t2 26.5955
R16217 SWN[8].n3 SWN[8].t3 26.5955
R16218 SWN[8].n0 SWN[8].t0 24.9236
R16219 SWN[8].n0 SWN[8].t1 24.9236
R16220 SWN[8] SWN[8].n5 14.676
R16221 SWN[8] SWN[8].n4 10.4965
R16222 SWN[8].n2 SWN[8] 10.4965
R16223 SWN[8].n4 SWN[8] 6.9125
R16224 SWN[8].n2 SWN[8] 6.9125
R16225 SWN[8].n5 SWN[8] 4.3525
R16226 SWN[8].n1 SWN[8] 1.7925
R16227 a_n1544_2717.t1 a_n1544_2717.n3 370.026
R16228 a_n1544_2717.n0 a_n1544_2717.t3 351.356
R16229 a_n1544_2717.n1 a_n1544_2717.t2 334.717
R16230 a_n1544_2717.n3 a_n1544_2717.t0 325.971
R16231 a_n1544_2717.n1 a_n1544_2717.t5 309.935
R16232 a_n1544_2717.n0 a_n1544_2717.t4 305.683
R16233 a_n1544_2717.n2 a_n1544_2717.n0 16.879
R16234 a_n1544_2717.n3 a_n1544_2717.n2 10.8867
R16235 a_n1544_2717.n2 a_n1544_2717.n1 9.3005
R16236 a_n629_2717.n3 a_n629_2717.n2 636.953
R16237 a_n629_2717.n1 a_n629_2717.t5 366.856
R16238 a_n629_2717.n2 a_n629_2717.n0 300.2
R16239 a_n629_2717.n2 a_n629_2717.n1 225.036
R16240 a_n629_2717.n1 a_n629_2717.t4 174.056
R16241 a_n629_2717.n0 a_n629_2717.t1 70.0005
R16242 a_n629_2717.n3 a_n629_2717.t3 68.0124
R16243 a_n629_2717.t0 a_n629_2717.n3 63.3219
R16244 a_n629_2717.n0 a_n629_2717.t2 61.6672
R16245 a_6945_n9484.t0 a_6945_n9484.t1 60.0005
R16246 a_1412_2717.t0 a_1412_2717.t1 94.7268
R16247 a_n126_n9662.t0 a_n126_n9662.t1 87.1434
R16248 a_1452_n9650.n3 a_1452_n9650.n2 636.953
R16249 a_1452_n9650.n1 a_1452_n9650.t4 366.856
R16250 a_1452_n9650.n2 a_1452_n9650.n0 300.2
R16251 a_1452_n9650.n2 a_1452_n9650.n1 225.036
R16252 a_1452_n9650.n1 a_1452_n9650.t5 174.056
R16253 a_1452_n9650.n0 a_1452_n9650.t1 70.0005
R16254 a_1452_n9650.n3 a_1452_n9650.t2 68.0124
R16255 a_1452_n9650.t0 a_1452_n9650.n3 63.3219
R16256 a_1452_n9650.n0 a_1452_n9650.t3 61.6672
R16257 a_1806_n9662.t0 a_1806_n9662.t1 87.1434
R16258 a_7357_n9484.t0 a_7357_n9484.t1 94.7268
R16259 a_n4182_n10028.t0 a_n4182_n10028.t1 126.644
R16260 a_8574_3083.t0 a_8574_3083.n0 1327.82
R16261 a_8574_3083.n0 a_8574_3083.t1 194.655
R16262 a_8574_3083.n0 a_8574_3083.t2 63.3219
R16263 a_9661_n4742.t0 a_9661_n4742.t1 77.1434
R16264 DOUT[6].n3 DOUT[6].n2 585
R16265 DOUT[6].n4 DOUT[6].n3 585
R16266 DOUT[6].n1 DOUT[6].n0 185
R16267 DOUT[6] DOUT[6].n1 49.0339
R16268 DOUT[6].n3 DOUT[6].t2 26.5955
R16269 DOUT[6].n3 DOUT[6].t3 26.5955
R16270 DOUT[6].n0 DOUT[6].t0 24.9236
R16271 DOUT[6].n0 DOUT[6].t1 24.9236
R16272 DOUT[6] DOUT[6].n4 20.4368
R16273 DOUT[6].n2 DOUT[6] 15.6165
R16274 DOUT[6].n1 DOUT[6] 10.4965
R16275 DOUT[6].n4 DOUT[6] 1.7925
R16276 DOUT[6].n2 DOUT[6] 1.7925
R16277 a_n4647_n9484.t0 a_n4647_n9484.t1 60.0005
R16278 a_8711_n9484.t1 a_8711_n9484.t0 198.571
R16279 a_8877_n9484.t0 a_8877_n9484.t1 60.0005
R16280 a_n5922_n9662.t0 a_n5922_n9662.t1 87.1434
R16281 a_6315_n5258.n3 a_6315_n5258.n2 647.119
R16282 a_6315_n5258.n1 a_6315_n5258.t4 350.253
R16283 a_6315_n5258.n2 a_6315_n5258.n0 260.339
R16284 a_6315_n5258.n2 a_6315_n5258.n1 246.119
R16285 a_6315_n5258.n1 a_6315_n5258.t5 189.588
R16286 a_6315_n5258.n3 a_6315_n5258.t1 89.1195
R16287 a_6315_n5258.n0 a_6315_n5258.t0 63.3338
R16288 a_6315_n5258.t3 a_6315_n5258.n3 41.0422
R16289 a_6315_n5258.n0 a_6315_n5258.t2 31.9797
R16290 a_6568_n1573.t0 a_6568_n1573.t1 126.644
R16291 a_4833_n1029.t0 a_4833_n1029.t1 60.0005
R16292 a_n6579_n9484.t0 a_n6579_n9484.t1 60.0005
R16293 SWN[3].n4 SWN[3].n3 585
R16294 SWN[3].n3 SWN[3].n2 585
R16295 SWN[3].n1 SWN[3].n0 185
R16296 SWN[3].n5 SWN[3].n1 53.3859
R16297 SWN[3].n3 SWN[3].t3 26.5955
R16298 SWN[3].n3 SWN[3].t2 26.5955
R16299 SWN[3].n0 SWN[3].t0 24.9236
R16300 SWN[3].n0 SWN[3].t1 24.9236
R16301 SWN[3] SWN[3].n5 14.6588
R16302 SWN[3] SWN[3].n4 10.4965
R16303 SWN[3].n2 SWN[3] 10.4965
R16304 SWN[3].n4 SWN[3] 6.9125
R16305 SWN[3].n2 SWN[3] 6.9125
R16306 SWN[3].n5 SWN[3] 4.3525
R16307 SWN[3].n1 SWN[3] 1.7925
R16308 a_5245_n1029.t0 a_5245_n1029.t1 94.7268
R16309 SWN[7].n4 SWN[7].n3 585
R16310 SWN[7].n3 SWN[7].n2 585
R16311 SWN[7].n1 SWN[7].n0 185
R16312 SWN[7].n5 SWN[7].n1 53.3859
R16313 SWN[7].n3 SWN[7].t3 26.5955
R16314 SWN[7].n3 SWN[7].t2 26.5955
R16315 SWN[7].n0 SWN[7].t1 24.9236
R16316 SWN[7].n0 SWN[7].t0 24.9236
R16317 SWN[7] SWN[7].n5 14.6803
R16318 SWN[7] SWN[7].n4 10.4965
R16319 SWN[7].n2 SWN[7] 10.4965
R16320 SWN[7].n4 SWN[7] 6.9125
R16321 SWN[7].n2 SWN[7] 6.9125
R16322 SWN[7].n5 SWN[7] 4.3525
R16323 SWN[7].n1 SWN[7] 1.7925
R16324 a_6599_n1029.t0 a_6599_n1029.t1 198.571
R16325 a_6765_n1029.t0 a_6765_n1029.t1 60.0005
R16326 a_5167_2717.n3 a_5167_2717.n2 636.953
R16327 a_5167_2717.n1 a_5167_2717.t4 366.856
R16328 a_5167_2717.n2 a_5167_2717.n0 300.2
R16329 a_5167_2717.n2 a_5167_2717.n1 225.036
R16330 a_5167_2717.n1 a_5167_2717.t5 174.056
R16331 a_5167_2717.n0 a_5167_2717.t2 70.0005
R16332 a_5167_2717.t0 a_5167_2717.n3 68.0124
R16333 a_5167_2717.n3 a_5167_2717.t3 63.3219
R16334 a_5167_2717.n0 a_5167_2717.t1 61.6672
R16335 a_6176_n4702.t0 a_6176_n4702.t1 198.571
R16336 a_6529_n5258.t0 a_6529_n5258.n0 1327.82
R16337 a_6529_n5258.n0 a_6529_n5258.t2 194.655
R16338 a_6529_n5258.n0 a_6529_n5258.t1 63.3219
R16339 a_4698_2717.t1 a_4698_2717.t0 198.571
R16340 a_n2058_n9484.t0 a_n2058_n9484.t1 87.1434
R16341 a_n2881_n9484.t1 a_n2881_n9484.t0 198.571
R16342 a_4014_n5624.t0 a_4014_n5624.t1 87.1434
R16343 a_n6745_n9484.t0 a_n6745_n9484.t1 198.571
R16344 a_2927_n10028.n0 a_2927_n10028.t1 1327.82
R16345 a_2927_n10028.n0 a_2927_n10028.t2 194.655
R16346 a_2927_n10028.t0 a_2927_n10028.n0 63.3219
R16347 a_4244_n4702.t1 a_4244_n4702.t0 198.571
R16348 a_4410_n4714.t0 a_4410_n4714.t1 60.0005
R16349 a_n2869_n9118.n0 a_n2869_n9118.t2 1327.82
R16350 a_n2869_n9118.t0 a_n2869_n9118.n0 194.655
R16351 a_n2869_n9118.n0 a_n2869_n9118.t1 63.3219
R16352 a_5185_n1207.t1 a_5185_n1207.t0 198.571
R16353 a_189_n4714.n1 a_189_n4714.n0 926.024
R16354 a_189_n4714.t0 a_189_n4714.n1 82.0838
R16355 a_189_n4714.n0 a_189_n4714.t1 63.3338
R16356 a_189_n4714.n1 a_189_n4714.t3 63.3219
R16357 a_189_n4714.n0 a_189_n4714.t2 29.7268
R16358 a_n4235_n9484.t0 a_n4235_n9484.t1 94.7268
R16359 a_4656_n9662.n1 a_4656_n9662.n0 926.024
R16360 a_4656_n9662.t1 a_4656_n9662.n1 82.0838
R16361 a_4656_n9662.n0 a_4656_n9662.t0 63.3338
R16362 a_4656_n9662.n1 a_4656_n9662.t3 63.3219
R16363 a_4656_n9662.n0 a_4656_n9662.t2 29.7268
R16364 a_n1045_n9484.n3 a_n1045_n9484.n2 674.338
R16365 a_n1045_n9484.n1 a_n1045_n9484.t5 332.58
R16366 a_n1045_n9484.n2 a_n1045_n9484.n0 284.012
R16367 a_n1045_n9484.n2 a_n1045_n9484.n1 253.648
R16368 a_n1045_n9484.n1 a_n1045_n9484.t4 168.701
R16369 a_n1045_n9484.t0 a_n1045_n9484.n3 96.1553
R16370 a_n1045_n9484.n3 a_n1045_n9484.t3 65.6672
R16371 a_n1045_n9484.n0 a_n1045_n9484.t1 65.0005
R16372 a_n1045_n9484.n0 a_n1045_n9484.t2 45.0005
R16373 a_6796_2717.t0 a_6796_2717.t1 60.0005
R16374 a_6186_n5624.n0 a_6186_n5624.t0 68.3338
R16375 a_6186_n5624.n0 a_6186_n5624.t1 26.3935
R16376 a_6186_n5624.n1 a_6186_n5624.n0 14.4005
R16377 a_5521_2717.t0 a_5521_2717.t1 87.1434
R16378 a_9289_n9650.n0 a_9289_n9650.t0 68.3338
R16379 a_9289_n9650.n0 a_9289_n9650.t1 26.3935
R16380 a_9289_n9650.n1 a_9289_n9650.n0 14.4005
R16381 a_n3990_n9484.t0 a_n3990_n9484.t1 87.1434
R16382 a_1614_n10028.t0 a_1614_n10028.t1 126.644
R16383 a_5946_n5624.t0 a_5946_n5624.t1 87.1434
R16384 a_6228_n5482.n1 a_6228_n5482.t6 530.01
R16385 a_6228_n5482.t1 a_6228_n5482.n5 421.021
R16386 a_6228_n5482.n0 a_6228_n5482.t2 337.171
R16387 a_6228_n5482.n3 a_6228_n5482.t0 280.223
R16388 a_6228_n5482.n4 a_6228_n5482.t5 263.173
R16389 a_6228_n5482.n4 a_6228_n5482.t7 227.826
R16390 a_6228_n5482.n0 a_6228_n5482.t4 199.762
R16391 a_6228_n5482.n2 a_6228_n5482.n1 170.81
R16392 a_6228_n5482.n2 a_6228_n5482.n0 167.321
R16393 a_6228_n5482.n5 a_6228_n5482.n4 152
R16394 a_6228_n5482.n1 a_6228_n5482.t3 141.923
R16395 a_6228_n5482.n3 a_6228_n5482.n2 10.8376
R16396 a_6228_n5482.n5 a_6228_n5482.n3 2.50485
R16397 a_6369_n1207.t0 a_6369_n1207.t1 87.1434
R16398 a_n5004_n9484.n1 a_n5004_n9484.n0 926.024
R16399 a_n5004_n9484.t0 a_n5004_n9484.n1 82.0838
R16400 a_n5004_n9484.n0 a_n5004_n9484.t3 63.3338
R16401 a_n5004_n9484.n1 a_n5004_n9484.t2 63.3219
R16402 a_n5004_n9484.n0 a_n5004_n9484.t1 29.7268
R16403 a_4820_2959.n3 a_4820_2959.n2 647.119
R16404 a_4820_2959.n1 a_4820_2959.t5 350.253
R16405 a_4820_2959.n2 a_4820_2959.n0 260.339
R16406 a_4820_2959.n2 a_4820_2959.n1 246.119
R16407 a_4820_2959.n1 a_4820_2959.t4 189.588
R16408 a_4820_2959.n3 a_4820_2959.t0 89.1195
R16409 a_4820_2959.n0 a_4820_2959.t1 63.3338
R16410 a_4820_2959.t3 a_4820_2959.n3 41.0422
R16411 a_4820_2959.n0 a_4820_2959.t2 31.9797
R16412 a_2281_n5258.t0 a_2281_n5258.t1 126.644
R16413 a_3344_2717.t0 a_3344_2717.t1 94.7268
R16414 a_n6745_n9650.t1 a_n6745_n9650.t0 198.571
R16415 a_4699_3557.t1 a_4699_3557.t0 198.571
R16416 a_1561_n9650.n0 a_1561_n9650.t1 68.3338
R16417 a_1561_n9650.n0 a_1561_n9650.t0 26.3935
R16418 a_1561_n9650.n1 a_1561_n9650.n0 14.4005
R16419 a_9487_n4848.n2 a_9487_n4848.n0 672.948
R16420 a_9487_n4848.t0 a_9487_n4848.n2 314.563
R16421 a_9487_n4848.n1 a_9487_n4848.t4 236.18
R16422 a_9487_n4848.n1 a_9487_n4848.t3 163.881
R16423 a_9487_n4848.n2 a_9487_n4848.n1 152
R16424 a_9487_n4848.n0 a_9487_n4848.t1 63.3219
R16425 a_9487_n4848.n0 a_9487_n4848.t2 63.3219
R16426 a_5013_n9484.t0 a_5013_n9484.t1 60.0005
R16427 SWP[0].n0 SWP[0].t4 332.312
R16428 SWP[0].n0 SWP[0].t5 295.627
R16429 SWP[0].n3 SWP[0].n2 289.096
R16430 SWP[0] SWP[0].n0 196.004
R16431 SWP[0].n5 SWP[0].n4 185
R16432 SWP[0].n1 SWP[0] 49.3509
R16433 SWP[0] SWP[0].n5 49.0339
R16434 SWP[0].n2 SWP[0].t2 26.5955
R16435 SWP[0].n2 SWP[0].t3 26.5955
R16436 SWP[0] SWP[0].n1 26.3678
R16437 SWP[0].n4 SWP[0].t0 24.9236
R16438 SWP[0].n4 SWP[0].t1 24.9236
R16439 SWP[0] SWP[0].n6 14.5963
R16440 SWP[0].n6 SWP[0] 13.0565
R16441 SWP[0].n1 SWP[0] 11.211
R16442 SWP[0].n5 SWP[0] 10.4965
R16443 SWP[0] SWP[0].n3 9.48653
R16444 SWP[0].n3 SWP[0] 7.7181
R16445 SWP[0].n6 SWP[0] 4.3525
R16446 a_7045_n1207.t0 a_7045_n1207.t1 60.0005
R16447 a_n949_n9484.t0 a_n949_n9484.t1 198.571
R16448 a_9385_2717.t0 a_9385_2717.t1 87.1434
R16449 a_6952_n1573.n0 a_6952_n1573.t2 1327.82
R16450 a_6952_n1573.t0 a_6952_n1573.n0 194.655
R16451 a_6952_n1573.n0 a_6952_n1573.t1 63.3219
R16452 a_8541_n1207.t1 a_8541_n1207.t0 94.7268
R16453 a_2927_n9118.n0 a_2927_n9118.t1 1327.82
R16454 a_2927_n9118.n0 a_2927_n9118.t2 194.655
R16455 a_2927_n9118.t0 a_2927_n9118.n0 63.3219
R16456 a_7496_n5074.n1 a_7496_n5074.t2 530.01
R16457 a_7496_n5074.t1 a_7496_n5074.n5 421.021
R16458 a_7496_n5074.n0 a_7496_n5074.t5 337.142
R16459 a_7496_n5074.n3 a_7496_n5074.t0 280.223
R16460 a_7496_n5074.n4 a_7496_n5074.t6 263.173
R16461 a_7496_n5074.n4 a_7496_n5074.t4 227.826
R16462 a_7496_n5074.n0 a_7496_n5074.t3 199.762
R16463 a_7496_n5074.n2 a_7496_n5074.n1 170.81
R16464 a_7496_n5074.n2 a_7496_n5074.n0 167.321
R16465 a_7496_n5074.n5 a_7496_n5074.n4 152
R16466 a_7496_n5074.n1 a_7496_n5074.t7 141.923
R16467 a_7496_n5074.n3 a_7496_n5074.n2 10.8376
R16468 a_7496_n5074.n5 a_7496_n5074.n3 2.50485
R16469 a_8120_n5080.t0 a_8120_n5080.n0 1327.82
R16470 a_8120_n5080.n0 a_8120_n5080.t1 194.655
R16471 a_8120_n5080.n0 a_8120_n5080.t2 63.3219
R16472 a_5670_n9484.t0 a_5670_n9484.t1 87.1434
R16473 a_n275_2717.t0 a_n275_2717.t1 87.1434
R16474 a_6797_3557.t0 a_6797_3557.t1 60.0005
R16475 a_5522_3557.t0 a_5522_3557.t1 87.1434
R16476 a_2724_n9662.n1 a_2724_n9662.n0 926.024
R16477 a_2724_n9662.t0 a_2724_n9662.n1 82.0838
R16478 a_2724_n9662.n0 a_2724_n9662.t3 63.3338
R16479 a_2724_n9662.n1 a_2724_n9662.t2 63.3219
R16480 a_2724_n9662.n0 a_2724_n9662.t1 29.7268
R16481 a_8977_n1207.t0 a_8977_n1207.t1 60.0005
R16482 a_9049_n1207.t1 a_9049_n1207.t0 198.571
R16483 a_3493_n9484.t1 a_3493_n9484.t0 94.7268
R16484 a_4822_n4702.n0 a_4822_n4702.t0 68.3338
R16485 a_4822_n4702.n0 a_4822_n4702.t1 26.3935
R16486 a_4822_n4702.n1 a_4822_n4702.n0 14.4005
R16487 a_7602_n9662.t0 a_7602_n9662.t1 87.1434
R16488 a_3345_3557.t1 a_3345_3557.t0 94.7268
R16489 a_n2715_n9484.t0 a_n2715_n9484.t1 60.0005
R16490 a_4690_n5624.t0 a_4690_n5624.t1 60.0005
R16491 a_9386_3557.t0 a_9386_3557.t1 87.1434
R16492 a_2901_n1029.t0 a_2901_n1029.t1 60.0005
R16493 a_n937_n9118.n0 a_n937_n9118.t2 1327.82
R16494 a_n937_n9118.n0 a_n937_n9118.t1 194.655
R16495 a_n937_n9118.t0 a_n937_n9118.n0 63.3219
R16496 a_4875_n5080.t0 a_4875_n5080.t1 126.644
R16497 a_2704_n1573.t0 a_2704_n1573.t1 126.644
R16498 a_5067_n4714.t0 a_5067_n4714.t1 87.1434
R16499 a_n4813_n9650.t1 a_n4813_n9650.t0 198.571
R16500 a_8877_n9662.t0 a_8877_n9662.t1 60.0005
R16501 a_n6114_n9118.t0 a_n6114_n9118.t1 126.644
R16502 a_2082_n5624.t0 a_2082_n5624.t1 87.1434
R16503 a_n6579_n9662.t0 a_n6579_n9662.t1 60.0005
R16504 a_7410_n10028.t0 a_7410_n10028.t1 126.644
R16505 a_6609_n1207.t1 a_6609_n1207.t0 94.7268
R16506 a_5478_n9118.t0 a_5478_n9118.t1 126.644
R16507 a_n2303_n9484.t0 a_n2303_n9484.t1 94.7268
R16508 a_4254_n5624.n0 a_4254_n5624.t1 68.3338
R16509 a_4254_n5624.n0 a_4254_n5624.t0 26.3935
R16510 a_4254_n5624.n1 a_4254_n5624.n0 14.4005
R16511 a_3081_n9484.t0 a_3081_n9484.t1 60.0005
R16512 a_3589_2717.t0 a_3589_2717.t1 87.1434
R16513 a_5113_n1207.t0 a_5113_n1207.t1 60.0005
R16514 a_n7854_n9484.t0 a_n7854_n9484.t1 87.1434
R16515 a_2943_n5080.t0 a_2943_n5080.t1 126.644
R16516 a_n783_n9484.t0 a_n783_n9484.t1 60.0005
R16517 a_9109_n1029.t1 a_9109_n1029.t0 94.7268
R16518 a_5013_n9662.t0 a_5013_n9662.t1 60.0005
R16519 a_4847_n9650.t1 a_4847_n9650.t0 198.571
R16520 a_n8677_n9484.t1 a_n8677_n9484.t0 198.571
C0 CF[5] CF[4] 10.218201f
C1 CF[5] SWN[6] 0.061496f
C2 VSSD SWN[3] 3.60764f
C3 CF[6] SWP[4] 0.067225f
C4 CF[8] SWP[1] 0.065113f
C5 auto_sampling_0.x7.Q EN 0.022065f
C6 CF[5] COMP_N 0.062035f
C7 out_latch_0.FINAL CKO 0.222681f
C8 out_latch_0.FINAL SWP[4] 0.089194f
C9 out_latch_0.FINAL DOUT[0] 0.173136f
C10 CF[6] SWN[4] 0.128503f
C11 out_latch_0.FINAL DOUT[7] 0.171243f
C12 CF[7] SWP[8] 0.062091f
C13 CKO SWP[1] 0.038863f
C14 CF[9] SWP[3] 0.071213f
C15 SWP[1] SWP[4] 0.127316f
C16 cdac_ctrl_0.x1.X CF[1] 0.03374f
C17 SWP[1] DOUT[0] 0.086605f
C18 SWP[3] SWP[0] 0.369772f
C19 auto_sampling_0.x5.D EN 0.022065f
C20 CLKSB DOUT[2] 0.075355f
C21 CLKSB DOUT[5] 0.075489f
C22 CF[9] SWN[9] 0.075326f
C23 CF[7] SWN[2] 0.131673f
C24 SWP[0] SWN[9] 5.70956f
C25 CF[4] SWP[3] 0.102408f
C26 SWP[5] SWN[8] 0.061785f
C27 SWP[3] SWN[6] 0.061504f
C28 SWP[1] SWN[4] 0.065886f
C29 cdac_ctrl_0.x1.X CF[5] 0.03374f
C30 cdac_ctrl_0.x2.X VDDD 13.660901f
C31 cdac_ctrl_0.x2.X SWN[0] 0.077566f
C32 cdac_ctrl_0.x2.X CLKS 0.655767f
C33 CF[4] SWN[9] 0.07529f
C34 VDDD CF[8] 1.19473f
C35 SWP[3] COMP_N 0.112017f
C36 CKO DOUT[8] 0.136361f
C37 SWN[7] SWN[8] 8.93889f
C38 SWN[6] SWN[9] 0.062245f
C39 CF[8] SWN[0] 0.450475f
C40 VSSD CF[6] 4.2129f
C41 CLKS CF[8] 0.184685f
C42 CF[3] SWP[5] 0.06747f
C43 SWP[6] COMP_P 0.106289f
C44 DOUT[2] DOUT[6] 0.050572f
C45 DOUT[0] DOUT[8] 0.05229f
C46 DOUT[7] DOUT[8] 16.0942f
C47 DOUT[5] DOUT[6] 14.9485f
C48 SWP[9] COMP_P 0.106279f
C49 DOUT[1] DOUT[2] 12.0577f
C50 DOUT[3] DOUT[4] 12.347301f
C51 DOUT[1] DOUT[5] 0.057777f
C52 COMP_N SWN[9] 0.062035f
C53 VDDD CKO 6.1211f
C54 out_latch_0.FINAL VSSD 14.2655f
C55 CF[3] SWN[7] 0.062015f
C56 VDDD SWP[4] 0.72212f
C57 CLKS CKO 0.549538f
C58 VDDD DOUT[0] 1.01385f
C59 CF[2] SWP[2] 0.068288f
C60 VDDD DOUT[7] 0.894441f
C61 COMP_P SWN[3] 0.062287f
C62 CF[2] DOUT[9] 0.031889f
C63 CF[2] SWP[7] 0.062625f
C64 SWP[8] SWN[2] 0.067874f
C65 SWP[6] SWN[1] 0.065124f
C66 SWP[4] SWN[0] 0.075119f
C67 CLKS DOUT[0] 0.308894f
C68 SWP[9] SWN[1] 0.065124f
C69 CLKS SWP[4] 0.120302f
C70 CLKS DOUT[7] 0.305978f
C71 VSSD SWP[1] 4.83543f
C72 auto_sampling_0.x11.D EN 0.029189f
C73 CF[0] DOUT[9] 0.161343f
C74 CF[0] SWP[2] 0.075652f
C75 CF[0] SWP[7] 0.069989f
C76 cdac_ctrl_0.x1.X SWP[3] 0.083576f
C77 VDDD SWN[4] 0.413667f
C78 CF[2] SWN[5] 0.064173f
C79 SWN[0] SWN[4] 0.075469f
C80 SWN[1] SWN[3] 0.066474f
C81 CF[1] SWP[6] 0.067837f
C82 CLKS SWN[4] 0.024253f
C83 CF[1] SWP[9] 0.075687f
C84 auto_sampling_0.x12.D VDDD 3.31755f
C85 CF[0] SWN[5] 0.071538f
C86 EN SWP[0] 0.098973f
C87 CF[1] SWN[3] 0.065379f
C88 CF[5] SWP[6] 0.067886f
C89 VSSD DOUT[8] 3.4192f
C90 CF[5] SWP[9] 0.075825f
C91 out_latch_0.FINAL CLKSB 0.179085f
C92 VDDD VSSD 1.84148p
C93 CF[5] SWN[3] 0.127707f
C94 CF[6] COMP_P 0.058086f
C95 VSSD SWN[0] 6.34788f
C96 VSSD CLKS 45.3641f
C97 CLK CF[8] 0.211173f
C98 cdac_ctrl_0.x2.X SWN[8] 0.07755f
C99 out_latch_0.FINAL DOUT[6] 0.171245f
C100 CF[8] SWN[8] 0.061784f
C101 out_latch_0.FINAL DOUT[1] 0.1711f
C102 CF[6] SWN[1] 0.12732f
C103 CLK CKO 0.178011f
C104 auto_sampling_0.x22.A VDDD 1.03914f
C105 CF[9] SWP[0] 0.072959f
C106 SWP[1] COMP_P 0.107116f
C107 SWP[3] DOUT[2] 0.084169f
C108 CLK DOUT[0] 0.144134f
C109 SWP[3] SWP[6] 0.136932f
C110 CLK DOUT[7] 0.142691f
C111 SWP[5] SWP[2] 0.383692f
C112 cdac_ctrl_0.x2.X CF[3] 0.074929f
C113 SWP[5] SWP[7] 0.13303f
C114 SWP[3] SWP[9] 0.136546f
C115 SWP[1] DOUT[1] 0.011518f
C116 CLKSB DOUT[8] 0.075904f
C117 CF[8] CF[3] 0.126634f
C118 CF[6] CF[1] 0.12516f
C119 CF[9] CF[4] 0.140036f
C120 CF[7] CF[2] 0.127417f
C121 CF[9] SWN[6] 0.121634f
C122 SWP[6] SWN[9] 0.075428f
C123 CF[4] SWP[0] 0.072959f
C124 SWP[4] SWN[8] 0.061798f
C125 SWP[2] SWN[7] 0.062085f
C126 SWP[0] SWN[6] 0.061583f
C127 SWP[9] SWN[9] 0.182717f
C128 SWP[7] SWN[7] 0.070414f
C129 SWP[5] SWN[5] 0.072572f
C130 SWP[1] SWN[1] 0.073523f
C131 SWP[3] SWN[3] 0.073755f
C132 VDDD CLKSB 0.830232f
C133 CF[7] CF[0] 0.141229f
C134 CF[9] COMP_N 0.062035f
C135 auto_sampling_0.x12.D CLK 1.56089f
C136 CLKS CLKSB 11.3385f
C137 SWP[0] COMP_N 0.11219f
C138 CF[4] SWN[6] 0.061492f
C139 SWN[3] SWN[9] 0.065524f
C140 SWN[5] SWN[7] 0.066052f
C141 SWN[4] SWN[8] 0.066242f
C142 CF[6] CF[5] 10.6877f
C143 CF[3] SWP[4] 0.067118f
C144 auto_sampling_0.x12.D auto_sampling_0.x14.D 0.012731f
C145 DOUT[6] DOUT[8] 0.053038f
C146 CF[1] SWP[1] 0.065061f
C147 auto_sampling_0.x12.D auto_sampling_0.x11.Q 0.081966f
C148 DOUT[1] DOUT[8] 0.051693f
C149 CF[4] COMP_N 0.062035f
C150 COMP_N SWN[6] 0.062092f
C151 CF[3] SWN[4] 0.065879f
C152 VDDD COMP_P 0.556762f
C153 VDDD DOUT[6] 0.941062f
C154 CF[2] SWP[8] 0.061875f
C155 VDDD DOUT[1] 0.902635f
C156 COMP_P SWN[0] 5.70012f
C157 CLKS COMP_P 0.077648f
C158 CLKS DOUT[6] 0.305633f
C159 CF[5] SWP[1] 0.065113f
C160 CLKS DOUT[1] 0.305226f
C161 VSSD CLK 11.72f
C162 CF[0] SWP[8] 0.06924f
C163 cdac_ctrl_0.x1.X CF[9] 0.03374f
C164 cdac_ctrl_0.x1.X SWP[0] 0.083359f
C165 auto_sampling_0.x14.D VSSD 0.314301f
C166 CF[2] SWN[2] 0.067907f
C167 VDDD SWN[1] 0.373055f
C168 VSSD auto_sampling_0.x11.Q 0.351674f
C169 VSSD SWN[8] 2.36657f
C170 SWN[0] SWN[1] 15.4865f
C171 CLKS SWN[1] 0.01099f
C172 CF[6] SWP[3] 0.071145f
C173 cdac_ctrl_0.x1.X CF[4] 0.03374f
C174 CF[0] SWN[2] 0.075261f
C175 auto_sampling_0.x22.A CLK 0.189895f
C176 VDDD CF[1] 1.18878f
C177 EN DOUT[2] 0.299589f
C178 EN SWP[6] 0.076129f
C179 EN DOUT[5] 0.346286f
C180 VSSD CF[3] 5.06919f
C181 CF[6] SWN[9] 0.075305f
C182 CF[1] SWN[0] 0.789812f
C183 EN SWP[9] 0.100588f
C184 VDDD auto_sampling_0.x2.D 0.706808f
C185 CLKS CF[1] 0.236104f
C186 auto_sampling_0.x12.D auto_sampling_0.x15.D 0.012731f
C187 out_latch_0.FINAL SWP[3] 0.089175f
C188 CF[7] SWP[5] 0.067673f
C189 SWP[1] SWP[3] 0.130009f
C190 CLK CLKSB 5.78473f
C191 VDDD CF[5] 1.64383f
C192 CF[7] SWN[7] 0.06205f
C193 CF[5] SWN[0] 0.263737f
C194 CLKS CF[5] 0.238311f
C195 CF[8] SWP[2] 0.06835f
C196 SWP[1] SWN[9] 0.075877f
C197 CF[8] SWP[7] 0.094389f
C198 cdac_ctrl_0.x2.X SWN[5] 0.077721f
C199 auto_sampling_0.x15.D VSSD 0.315204f
C200 CKO DOUT[9] 0.181724f
C201 CKO SWP[2] 0.109854f
C202 CF[8] SWN[5] 0.125877f
C203 CKO SWP[7] 0.107342f
C204 CF[9] SWP[6] 0.068258f
C205 SWP[0] DOUT[2] 0.016951f
C206 SWP[2] SWP[4] 0.133771f
C207 CF[9] SWP[9] 5.71272f
C208 SWP[0] SWP[6] 0.139557f
C209 DOUT[7] DOUT[9] 0.073107f
C210 SWP[5] SWP[8] 0.132342f
C211 CLK DOUT[6] 0.142592f
C212 SWP[5] DOUT[4] 0.08397f
C213 DOUT[9] DOUT[0] 0.072233f
C214 SWP[7] SWP[4] 0.406981f
C215 SWP[9] SWP[0] 0.139468f
C216 SWP[5] DOUT[3] 0.013729f
C217 CLK DOUT[1] 0.142459f
C218 auto_sampling_0.x23.A auto_sampling_0.x24.A 0.391541f
C219 VDDD auto_sampling_0.x3.D 0.706808f
C220 auto_sampling_0.x12.D auto_sampling_0.x16.D 0.012731f
C221 CF[4] SWP[6] 0.067837f
C222 COMP_P SWN[8] 0.062035f
C223 CF[9] SWN[3] 0.127707f
C224 SWP[8] SWN[7] 0.062015f
C225 SWP[6] SWN[6] 0.069867f
C226 SWP[2] SWN[4] 0.065874f
C227 CF[4] SWP[9] 0.075782f
C228 SWP[4] SWN[5] 0.064173f
C229 VDDD SWP[3] 0.767483f
C230 SWP[0] SWN[3] 0.065392f
C231 SWP[9] SWN[6] 0.061468f
C232 SWP[7] SWN[4] 0.065851f
C233 SWP[5] SWN[2] 0.067874f
C234 SWP[3] SWN[0] 0.075119f
C235 CLKS SWP[3] 0.11927f
C236 SWP[6] COMP_N 0.111992f
C237 VDDD SWN[9] 0.455023f
C238 SWP[9] COMP_N 0.11198f
C239 CF[4] SWN[3] 0.57484f
C240 CF[3] COMP_P 0.058086f
C241 SWN[2] SWN[7] 0.068104f
C242 SWN[4] SWN[5] 10.4834f
C243 SWN[0] SWN[9] 0.075167f
C244 SWN[1] SWN[8] 0.065236f
C245 SWN[3] SWN[6] 0.066037f
C246 CLK CF[1] 0.130496f
C247 auto_sampling_0.x2.D CLK 0.104376f
C248 out_latch_0.FINAL EN 5.89978f
C249 COMP_N SWN[3] 0.062192f
C250 VDDD auto_sampling_0.x7.Q 0.706849f
C251 auto_sampling_0.x16.D VSSD 0.315204f
C252 CF[1] SWN[8] 0.061748f
C253 CF[3] SWN[1] 0.12732f
C254 EN SWP[1] 0.035003f
C255 VSSD SWP[2] 4.64915f
C256 CLK CF[5] 0.211098f
C257 VSSD DOUT[9] 6.4308f
C258 VSSD SWP[7] 3.30316f
C259 cdac_ctrl_0.x1.X SWP[6] 0.083749f
C260 cdac_ctrl_0.x2.X CF[7] 0.074929f
C261 CF[1] CF[3] 0.131478f
C262 VDDD auto_sampling_0.x5.D 0.706808f
C263 CF[5] SWN[8] 0.061757f
C264 auto_sampling_0.x12.D auto_sampling_0.x21.D 0.015303f
C265 CF[8] CF[7] 10.5645f
C266 CF[9] CF[6] 0.141621f
C267 VSSD SWN[5] 3.12581f
C268 CF[6] SWP[0] 0.072959f
C269 CF[0] CF[2] 0.145681f
C270 EN DOUT[8] 0.308662f
C271 CF[5] CF[3] 0.140947f
C272 CF[6] CF[4] 0.126922f
C273 CF[6] SWN[6] 0.061503f
C274 out_latch_0.FINAL SWP[0] 0.089329f
C275 CF[7] SWP[4] 0.06727f
C276 CF[9] SWP[1] 0.065113f
C277 auto_sampling_0.x3.D CLK 0.104379f
C278 VDDD EN 12.683001f
C279 SWP[1] SWP[0] 13.7247f
C280 CF[6] COMP_N 0.062035f
C281 auto_sampling_0.x21.D VSSD 0.315204f
C282 CLKSB DOUT[9] 0.076663f
C283 EN CLKS 0.298169f
C284 CF[7] SWN[4] 0.128503f
C285 CF[8] SWP[8] 0.062276f
C286 CF[4] SWP[1] 0.065113f
C287 SWP[1] SWN[6] 0.061539f
C288 SWP[3] SWN[8] 0.06182f
C289 out_latch_0.FINAL COMP_N 1.31352f
C290 cdac_ctrl_0.x2.X SWN[2] 0.077619f
C291 VDDD auto_sampling_0.x11.D 0.70687f
C292 SWN[8] SWN[9] 8.06844f
C293 SWP[1] COMP_N 0.112722f
C294 CKO DOUT[4] 0.210053f
C295 CKO SWP[8] 0.125201f
C296 auto_sampling_0.x7.Q CLK 0.104376f
C297 CF[8] SWN[2] 0.131673f
C298 CKO DOUT[3] 0.19924f
C299 CF[3] SWP[3] 0.071065f
C300 SWP[4] SWP[8] 0.131511f
C301 SWP[2] COMP_P 0.106384f
C302 SWP[7] COMP_P 0.10628f
C303 DOUT[0] DOUT[4] 0.062486f
C304 DOUT[9] DOUT[6] 0.072237f
C305 DOUT[7] DOUT[4] 0.050845f
C306 SWP[7] DOUT[6] 0.08358f
C307 DOUT[5] DOUT[2] 0.05807f
C308 SWP[9] SWP[6] 0.431255f
C309 DOUT[3] DOUT[0] 0.060198f
C310 DOUT[1] DOUT[9] 0.071677f
C311 DOUT[3] DOUT[7] 0.050571f
C312 cdac_ctrl_0.x1.X CF[6] 0.033738f
C313 VDDD CF[9] 1.16911f
C314 CF[3] SWN[9] 0.07529f
C315 VDDD SWP[0] 0.681865f
C316 VSSD CF[7] 4.28593f
C317 COMP_P SWN[5] 0.062143f
C318 SWP[8] SWN[4] 0.065851f
C319 CF[9] SWN[0] 1.72371f
C320 SWP[4] SWN[2] 0.067874f
C321 CLKS CF[9] 0.184498f
C322 SWP[6] SWN[3] 0.065356f
C323 SWP[2] SWN[1] 0.065124f
C324 CF[2] SWP[5] 0.06747f
C325 SWP[0] SWN[0] 0.083518f
C326 SWP[7] SWN[1] 0.065124f
C327 auto_sampling_0.x5.D CLK 0.104376f
C328 SWP[9] SWN[3] 0.065356f
C329 CLKS SWP[0] 0.10256f
C330 CF[0] SWP[5] 0.074835f
C331 VDDD CF[4] 1.45528f
C332 VDDD SWN[6] 0.471939f
C333 cdac_ctrl_0.x1.X SWP[1] 0.083508f
C334 CF[2] SWN[7] 0.062015f
C335 CF[4] SWN[0] 0.242352f
C336 CLKS CF[4] 0.183231f
C337 SWN[1] SWN[5] 0.065448f
C338 SWN[2] SWN[4] 0.069424f
C339 SWN[0] SWN[6] 0.075271f
C340 CF[1] DOUT[9] 0.059657f
C341 CF[1] SWP[2] 0.068288f
C342 CLKS SWN[6] 0.022102f
C343 CF[1] SWP[7] 0.062625f
C344 VDDD COMP_N 2.09563f
C345 CF[0] SWN[7] 0.069379f
C346 COMP_N SWN[0] 0.063172f
C347 CLKS COMP_N 0.062062f
C348 CF[1] SWN[5] 0.064173f
C349 CLK EN 15.6896f
C350 CF[5] SWP[2] 0.06835f
C351 VSSD SWP[8] 3.0427f
C352 CF[5] SWP[7] 0.062693f
C353 VSSD DOUT[4] 3.36149f
C354 VSSD DOUT[3] 3.34726f
C355 auto_sampling_0.x12.D auto_sampling_0.x21.Q 0.643519f
C356 auto_sampling_0.x14.D EN 0.025516f
C357 auto_sampling_0.x11.Q EN 0.010534f
C358 CF[5] SWN[5] 0.064207f
C359 CF[6] SWP[6] 0.067906f
C360 VSSD SWN[2] 3.98568f
C361 auto_sampling_0.x11.D CLK 0.075486f
C362 CF[6] SWP[9] 0.075909f
C363 cdac_ctrl_0.x1.X VDDD 13.6628f
C364 cdac_ctrl_0.x1.X CLKS 0.842598f
C365 out_latch_0.FINAL DOUT[2] 0.171142f
C366 out_latch_0.FINAL SWP[6] 0.089201f
C367 out_latch_0.FINAL DOUT[5] 0.171175f
C368 VSSD auto_sampling_0.x21.Q 2.338f
C369 CF[6] SWN[3] 0.127707f
C370 out_latch_0.FINAL SWP[9] 0.089111f
C371 CF[7] COMP_P 0.058086f
C372 CLK CF[9] 0.221334f
C373 SWP[1] SWP[6] 0.126979f
C374 SWP[3] SWP[2] 10.666901f
C375 SWP[3] SWP[7] 0.1367f
C376 SWP[1] SWP[9] 0.126871f
C377 CLKSB DOUT[4] 0.075452f
C378 CLKSB DOUT[3] 0.075423f
C379 CF[9] SWN[8] 0.360998f
C380 CF[7] SWN[1] 0.12732f
C381 CLK CF[4] 0.214221f
C382 SWP[2] SWN[9] 0.075597f
C383 SWP[0] SWN[8] 0.062251f
C384 auto_sampling_0.x22.A auto_sampling_0.x21.Q 0.016637f
C385 SWP[7] SWN[9] 0.075415f
C386 SWP[5] SWN[7] 0.062041f
C387 SWP[3] SWN[5] 0.064199f
C388 SWP[1] SWN[3] 0.065379f
C389 auto_sampling_0.x15.D EN 0.025516f
C390 auto_sampling_0.x23.A VSSD 0.575926f
C391 cdac_ctrl_0.x2.X CF[2] 0.074929f
C392 CF[4] SWN[8] 0.061748f
C393 CF[9] CF[3] 0.139944f
C394 CF[7] CF[1] 0.127325f
C395 CF[8] CF[2] 0.126543f
C396 SWN[5] SWN[9] 0.0646f
C397 SWN[6] SWN[8] 0.063299f
C398 CF[3] SWP[0] 0.072959f
C399 cdac_ctrl_0.x2.X CF[0] 0.110249f
C400 SWP[6] DOUT[8] 0.016637f
C401 SWP[8] COMP_P 0.106912f
C402 DOUT[4] DOUT[6] 0.051655f
C403 DOUT[2] DOUT[8] 0.051735f
C404 SWP[9] DOUT[8] 0.087888f
C405 DOUT[5] DOUT[8] 0.052227f
C406 DOUT[3] DOUT[6] 0.050858f
C407 DOUT[1] DOUT[4] 0.062129f
C408 CF[8] CF[0] 0.140406f
C409 DOUT[1] DOUT[3] 0.060353f
C410 COMP_N SWN[8] 0.062035f
C411 auto_sampling_0.x22.A auto_sampling_0.x23.A 0.149102f
C412 CF[3] CF[4] 12.4648f
C413 CF[3] SWN[6] 0.061468f
C414 VDDD SWP[6] 0.772231f
C415 CF[7] CF[5] 0.13116f
C416 VDDD DOUT[2] 0.942008f
C417 CF[2] SWP[4] 0.067118f
C418 VDDD DOUT[5] 0.881634f
C419 COMP_P SWN[2] 0.062503f
C420 VDDD SWP[9] 1.41577f
C421 SWP[8] SWN[1] 0.065124f
C422 SWP[6] SWN[0] 0.075119f
C423 CLKS SWP[6] 0.119813f
C424 SWP[9] SWN[0] 0.075119f
C425 CLKS DOUT[2] 0.305361f
C426 CLKS SWP[9] 0.100725f
C427 CLKS DOUT[5] 0.30545f
C428 CF[3] COMP_N 0.062035f
C429 CF[0] SWP[4] 0.074483f
C430 CF[0] DOUT[7] 0.020562f
C431 VDDD SWN[3] 0.397183f
C432 CF[2] SWN[4] 0.065874f
C433 CF[1] SWP[8] 0.061875f
C434 SWN[0] SWN[3] 0.075747f
C435 SWN[1] SWN[2] 12.197901f
C436 CLKS SWN[3] 0.02465f
C437 CF[6] SWP[1] 0.065113f
C438 auto_sampling_0.x16.D EN 0.025516f
C439 CF[0] SWN[4] 0.073215f
C440 EN SWP[2] 0.076264f
C441 EN DOUT[9] 0.238119f
C442 EN SWP[7] 0.086174f
C443 CF[1] SWN[2] 0.067901f
C444 CF[5] SWP[8] 0.06197f
C445 out_latch_0.FINAL SWP[1] 0.090696f
C446 CF[7] SWP[3] 0.071145f
C447 cdac_ctrl_0.x1.X CF[3] 0.03374f
C448 CF[7] SWN[9] 0.075315f
C449 CF[5] SWN[2] 0.131673f
C450 VSSD CF[2] 5.4997f
C451 CF[8] SWP[5] 0.067699f
C452 VSSD CF[0] 12.5597f
C453 cdac_ctrl_0.x2.X SWN[7] 0.077679f
C454 out_latch_0.FINAL DOUT[8] 0.171346f
C455 VDDD CF[6] 1.25811f
C456 CF[8] SWN[7] 0.401462f
C457 CF[6] SWN[0] 0.295933f
C458 CLKS CF[6] 0.237953f
C459 CKO SWP[5] 0.121231f
C460 CF[9] SWP[2] 0.068399f
C461 auto_sampling_0.x21.D EN 0.035599f
C462 CF[9] SWP[7] 0.063312f
C463 CLK DOUT[2] 0.142459f
C464 SWP[0] SWP[2] 0.142057f
C465 SWP[3] SWP[8] 0.137681f
C466 SWP[5] SWP[4] 10.7404f
C467 SWP[7] SWP[0] 0.139518f
C468 auto_sampling_0.x24.A VSSD 0.940294f
C469 CLK DOUT[5] 0.142557f
C470 out_latch_0.FINAL VDDD 3.97736f
C471 out_latch_0.FINAL CLKS 7.49005f
C472 CF[4] SWP[2] 0.06835f
C473 CF[9] SWN[5] 0.125877f
C474 SWP[8] SWN[9] 0.080982f
C475 SWP[6] SWN[8] 0.061773f
C476 SWP[2] SWN[6] 0.061517f
C477 CF[4] SWP[7] 0.062675f
C478 VDDD SWP[1] 0.749414f
C479 SWP[4] SWN[7] 0.062051f
C480 SWP[0] SWN[5] 0.064245f
C481 SWP[9] SWN[8] 0.061748f
C482 SWP[7] SWN[6] 0.061468f
C483 SWP[5] SWN[4] 0.065851f
C484 SWP[1] SWN[0] 0.075119f
C485 SWP[3] SWN[2] 0.067874f
C486 CLKS SWP[1] 0.103972f
C487 SWP[2] COMP_N 0.112047f
C488 CF[4] SWN[5] 0.064201f
C489 SWP[7] COMP_N 0.11198f
C490 SWN[4] SWN[7] 0.066554f
C491 SWN[2] SWN[9] 0.067993f
C492 SWN[5] SWN[6] 10.927099f
C493 SWN[3] SWN[8] 0.065598f
C494 CF[3] SWP[6] 0.067837f
C495 CF[3] SWP[9] 0.075755f
C496 COMP_N SWN[5] 0.062113f
C497 CF[3] SWN[3] 0.06539f
C498 VDDD DOUT[8] 0.957086f
C499 CF[2] COMP_P 0.058086f
C500 CLKS DOUT[8] 0.306859f
C501 VSSD SWP[5] 3.91254f
C502 CF[0] COMP_P 0.065349f
C503 CF[0] DOUT[6] 0.01178f
C504 cdac_ctrl_0.x1.X SWP[2] 0.08353f
C505 cdac_ctrl_0.x1.X SWP[7] 0.083769f
C506 CF[2] SWN[1] 0.670422f
C507 VDDD SWN[0] 0.367454f
C508 VDDD CLKS 9.31742f
C509 VSSD SWN[7] 2.60283f
C510 CLKS SWN[0] 0.010852f
C511 CLK CF[6] 0.112587f
C512 CF[0] SWN[1] 0.072516f
C513 cdac_ctrl_0.x2.X CF[8] 0.074945f
C514 CF[1] CF[2] 14.7825f
C515 EN SWP[8] 0.073685f
C516 EN DOUT[4] 0.318518f
C517 EN DOUT[3] 0.305539f
C518 CF[6] SWN[8] 0.061773f
C519 CF[9] CF[7] 0.143272f
C520 out_latch_0.FINAL CLK 5.81852f
C521 CF[7] SWP[0] 0.072959f
C522 CF[0] CF[1] 15.699f
C523 CF[5] CF[2] 0.139008f
C524 CF[6] CF[3] 0.125728f
C525 CF[7] CF[4] 0.127981f
C526 CF[7] SWN[6] 0.440553f
C527 CF[8] SWP[4] 0.067293f
C528 SWP[1] SWN[8] 0.061954f
C529 CF[5] CF[0] 0.198987f
C530 CF[7] COMP_N 0.062035f
C531 auto_sampling_0.x21.Q EN 0.494011f
C532 cdac_ctrl_0.x2.X SWN[4] 0.077679f
C533 CKO SWP[4] 0.112234f
C534 CKO DOUT[0] 5.37292f
C535 CF[8] SWN[4] 0.128503f
C536 CKO DOUT[7] 0.182985f
C537 CF[9] SWP[8] 0.094521f
C538 CF[3] SWP[1] 0.065113f
C539 CLK DOUT[8] 0.144029f
C540 SWP[2] SWP[6] 0.132239f
C541 SWP[0] SWP[8] 0.140578f
C542 DOUT[9] DOUT[2] 0.071717f
C543 SWP[7] SWP[6] 9.0391f
C544 SWP[5] COMP_P 0.106296f
C545 DOUT[7] DOUT[0] 0.050959f
C546 SWP[9] SWP[2] 0.132059f
C547 DOUT[5] DOUT[9] 0.071959f
C548 SWP[7] SWP[9] 0.162747f
C549 SWP[7] DOUT[5] 0.013729f
C550 CF[4] SWP[8] 0.061944f
C551 COMP_P SWN[7] 0.062091f
C552 SWP[8] SWN[6] 0.061468f
C553 CF[9] SWN[2] 0.131673f
C554 VDDD CLK 6.42539f
C555 SWP[6] SWN[5] 0.064173f
C556 SWP[4] SWN[4] 0.07425f
C557 SWP[2] SWN[3] 0.065356f
C558 CF[2] SWP[3] 0.071065f
C559 SWP[0] SWN[2] 0.067899f
C560 SWP[9] SWN[5] 0.064173f
C561 SWP[7] SWN[3] 0.065356f
C562 SWP[5] SWN[1] 0.065124f
C563 CLK CLKS 12.391099f
C564 cdac_ctrl_0.x1.X CF[7] 0.033738f
C565 auto_sampling_0.x14.D VDDD 0.705926f
C566 SWP[8] COMP_N 0.112617f
C567 VDDD auto_sampling_0.x11.Q 0.327961f
C568 CF[0] SWP[3] 0.078429f
C569 cdac_ctrl_0.x2.X VSSD 2.56323f
C570 VDDD SWN[8] 0.616893f
C571 CF[2] SWN[9] 0.07529f
C572 CF[4] SWN[2] 0.131673f
C573 SWN[3] SWN[5] 0.066853f
C574 SWN[1] SWN[7] 0.065274f
C575 SWN[0] SWN[8] 0.075203f
C576 SWN[2] SWN[6] 0.068233f
C577 CLKS SWN[8] 0.015293f
C578 VSSD CF[8] 4.29059f
C579 CF[1] SWP[5] 0.06747f
C580 CF[0] SWN[9] 0.099405f
C581 COMP_N SWN[2] 0.062288f
C582 VDDD CF[3] 1.26851f
C583 CF[1] SWN[7] 0.062015f
C584 VSSD CKO 7.58383f
C585 CF[3] SWN[0] 0.227324f
C586 CLKS CF[3] 0.183528f
C587 VSSD SWP[4] 4.13822f
C588 VSSD DOUT[0] 4.56258f
C589 CF[5] SWP[5] 0.06747f
C590 VSSD DOUT[7] 3.50706f
C591 cdac_ctrl_0.x1.X SWP[8] 0.082755f
C592 CF[5] SWN[7] 0.062039f
C593 VSSD SWN[4] 3.40309f
C594 CF[6] SWP[2] 0.06835f
C595 CF[6] SWP[7] 0.06272f
C596 auto_sampling_0.x12.D VSSD 2.51502f
C597 auto_sampling_0.x15.D VDDD 0.705036f
C598 out_latch_0.FINAL SWP[2] 0.089276f
C599 out_latch_0.FINAL DOUT[9] 0.192516f
C600 CF[6] SWN[5] 0.483326f
C601 out_latch_0.FINAL SWP[7] 0.089097f
C602 CF[7] SWP[6] 0.099394f
C603 CF[7] SWP[9] 0.07608f
C604 CLKSB CKO 0.093675f
C605 SWP[1] SWP[2] 12.5587f
C606 SWP[3] SWP[5] 0.138867f
C607 SWP[1] SWP[7] 0.126919f
C608 CLKSB DOUT[0] 0.076126f
C609 CLKSB DOUT[7] 0.075667f
C610 auto_sampling_0.x12.D auto_sampling_0.x22.A 0.042649f
C611 auto_sampling_0.x14.D CLK 0.100077f
C612 CF[7] SWN[3] 0.127707f
C613 CF[8] COMP_P 0.058086f
C614 SWP[3] SWN[7] 0.062064f
C615 SWP[5] SWN[9] 0.075442f
C616 SWP[1] SWN[5] 0.064222f
C617 cdac_ctrl_0.x2.X SWN[1] 0.07758f
C618 CKO DOUT[6] 0.188171f
C619 SWN[7] SWN[9] 0.063876f
C620 CF[8] SWN[1] 0.12732f
C621 CKO DOUT[1] 0.186066f
C622 auto_sampling_0.x24.A EN 0.014923f
C623 CLK CF[3] 0.213638f
C624 SWP[6] SWP[8] 0.134089f
C625 SWP[4] COMP_P 0.106307f
C626 DOUT[2] DOUT[4] 0.062987f
C627 SWP[4] DOUT[6] 0.016885f
C628 DOUT[9] DOUT[8] 15.940799f
C629 DOUT[0] DOUT[6] 0.051001f
C630 SWP[9] SWP[8] 8.24617f
C631 DOUT[7] DOUT[6] 15.3517f
C632 DOUT[5] DOUT[4] 11.5867f
C633 DOUT[3] DOUT[2] 11.553f
C634 DOUT[1] DOUT[0] 10.5082f
C635 auto_sampling_0.x16.D VDDD 0.705036f
C636 auto_sampling_0.x22.A VSSD 0.987372f
C637 DOUT[3] DOUT[5] 0.058899f
C638 DOUT[1] DOUT[7] 0.050371f
C639 cdac_ctrl_0.x2.X CF[1] 0.074929f
C640 CF[3] SWN[8] 0.061748f
C641 CF[8] CF[1] 0.126486f
C642 CF[9] CF[2] 0.139888f
C643 VDDD DOUT[9] 1.00964f
C644 VDDD SWP[2] 0.69293f
C645 SWP[8] SWN[3] 0.065356f
C646 VDDD SWP[7] 0.903703f
C647 COMP_P SWN[4] 0.062193f
C648 CF[2] SWP[0] 0.072959f
C649 SWP[4] SWN[1] 0.065124f
C650 SWP[6] SWN[2] 0.067874f
C651 SWP[2] SWN[0] 0.075119f
C652 SWP[7] SWN[0] 0.075119f
C653 CLKS SWP[2] 0.11853f
C654 SWP[9] SWN[2] 0.067874f
C655 CLKS DOUT[9] 5.95988f
C656 CLKS SWP[7] 0.117436f
C657 CF[9] CF[0] 0.15375f
C658 cdac_ctrl_0.x2.X CF[5] 0.074929f
C659 VSSD CLKSB 6.695509f
C660 CF[0] SWP[0] 0.080306f
C661 CF[2] CF[4] 0.142645f
C662 VDDD SWN[5] 0.440646f
C663 auto_sampling_0.x15.D CLK 0.100077f
C664 CF[2] SWN[6] 0.061468f
C665 CF[8] CF[5] 0.128226f
C666 CF[7] CF[6] 10.533099f
C667 CF[1] SWP[4] 0.067118f
C668 SWN[2] SWN[3] 12.177799f
C669 SWN[1] SWN[4] 0.065729f
C670 SWN[0] SWN[5] 0.075333f
C671 CLKS SWN[5] 0.023781f
C672 CF[0] CF[4] 0.153926f
C673 CF[0] SWN[6] 0.068833f
C674 CF[2] COMP_N 0.062035f
C675 EN SWP[5] 0.120944f
C676 CF[1] SWN[4] 0.065851f
C677 CF[0] COMP_N 0.070024f
C678 CF[5] SWP[4] 0.098488f
C679 VSSD COMP_P 6.17072f
C680 VSSD DOUT[6] 3.24308f
C681 VSSD DOUT[1] 3.13349f
C682 CF[7] SWP[1] 0.065113f
C683 auto_sampling_0.x21.D VDDD 0.705114f
C684 CF[5] SWN[4] 0.532142f
C685 CF[6] SWP[8] 0.062014f
C686 VSSD SWN[1] 4.04712f
C687 CF[8] SWP[3] 0.071193f
C688 cdac_ctrl_0.x1.X CF[2] 0.03374f
C689 auto_sampling_0.x16.D CLK 0.100077f
C690 out_latch_0.FINAL SWP[8] 0.107681f
C691 out_latch_0.FINAL DOUT[4] 0.171142f
C692 VSSD CF[1] 5.91701f
C693 CF[8] SWN[9] 0.07532f
C694 cdac_ctrl_0.x1.X CF[0] 0.056157f
C695 CF[6] SWN[2] 0.131673f
C696 out_latch_0.FINAL DOUT[3] 0.1711f
C697 CKO SWP[3] 0.104337f
C698 CF[9] SWP[5] 0.067743f
C699 VSSD auto_sampling_0.x2.D 0.311297f
C700 SWP[1] SWP[8] 0.127971f
C701 SWP[3] SWP[4] 9.93085f
C702 SWP[5] SWP[0] 0.139621f
C703 CLK DOUT[9] 0.155057f
C704 CLKSB DOUT[6] 0.075548f
C705 CLKSB DOUT[1] 0.075355f
C706 VDDD CF[7] 1.23618f
C707 VSSD CF[5] 4.739f
C708 CF[9] SWN[7] 0.122547f
C709 SWP[4] SWN[9] 0.075464f
C710 CF[7] SWN[0] 0.349351f
C711 SWP[2] SWN[8] 0.061861f
C712 SWP[0] SWN[7] 0.062225f
C713 CLKS CF[7] 0.185021f
C714 CF[4] SWP[5] 0.06747f
C715 SWP[7] SWN[8] 0.061748f
C716 SWP[3] SWN[4] 0.065851f
C717 SWP[5] SWN[6] 0.061468f
C718 SWP[1] SWN[2] 0.067874f
C719 CF[4] SWN[7] 0.062018f
C720 SWP[5] COMP_N 0.111991f
C721 SWN[5] SWN[8] 0.064959f
C722 SWN[6] SWN[7] 9.79241f
C723 SWN[4] SWN[9] 0.066099f
C724 CF[3] SWP[2] 0.099613f
C725 CF[3] DOUT[9] 0.016477f
C726 DOUT[4] DOUT[8] 0.05193f
C727 CF[3] SWP[7] 0.062625f
C728 DOUT[3] DOUT[8] 0.051804f
C729 DOUT[1] DOUT[6] 0.050439f
C730 COMP_N SWN[7] 0.062035f
C731 auto_sampling_0.x21.D CLK 0.07367f
C732 CF[3] SWN[5] 0.064197f
C733 VDDD SWP[8] 0.616847f
C734 VDDD DOUT[4] 0.937925f
C735 CF[2] SWP[6] 0.067837f
C736 VDDD DOUT[3] 0.894027f
C737 COMP_P SWN[1] 0.06318f
C738 SWP[8] SWN[0] 0.075119f
C739 VSSD auto_sampling_0.x3.D 0.311297f
C740 CF[2] SWP[9] 0.075735f
C741 CLKS SWP[8] 0.151374f
C742 CLKS DOUT[4] 0.305433f
C743 CLKS DOUT[3] 0.305338f
C744 VSSD SWP[3] 4.58346f
C745 CF[0] SWP[6] 0.075202f
C746 CF[0] SWP[9] 0.100166f
C747 VDDD SWN[2] 0.38389f
C748 cdac_ctrl_0.x1.X SWP[5] 0.08366f
C749 CF[2] SWN[3] 0.065384f
C750 CF[1] COMP_P 0.058086f
C751 SWN[0] SWN[2] 0.076646f
C752 VSSD SWN[9] 2.91841f
C753 CLKS SWN[2] 0.011042f
C754 CF[0] SWN[3] 0.072721f
C755 EN CKO 11.690901f
C756 VDDD auto_sampling_0.x21.Q 1.31897f
C757 EN SWP[4] 0.138573f
C758 EN DOUT[7] 0.299028f
C759 VSSD auto_sampling_0.x7.Q 0.311296f
C760 EN DOUT[0] 0.420831f
C761 CF[1] SWN[1] 0.065158f
C762 CF[5] COMP_P 0.058086f
C763 CLK CF[7] 0.210105f
C764 cdac_ctrl_0.x2.X CF[9] 0.073724f
C765 CF[5] SWN[1] 0.12732f
C766 CF[7] SWN[8] 0.061778f
C767 CF[9] CF[8] 10.9965f
C768 VSSD auto_sampling_0.x5.D 0.311297f
C769 auto_sampling_0.x12.D EN 1.94373f
C770 CF[8] SWP[0] 0.072959f
C771 auto_sampling_0.x23.A VDDD 0.517614f
C772 cdac_ctrl_0.x2.X CF[4] 0.074929f
C773 cdac_ctrl_0.x2.X SWN[6] 0.077716f
C774 CF[7] CF[3] 0.127597f
C775 CF[8] CF[4] 0.126807f
C776 CF[5] CF[1] 0.138208f
C777 CF[6] CF[2] 0.12533f
C778 CKO SWP[0] 0.021811f
C779 CF[8] SWN[6] 0.121634f
C780 CF[9] SWP[4] 0.067319f
C781 SWP[0] SWP[4] 0.139916f
C782 CLK DOUT[4] 0.142522f
C783 SWP[5] SWP[6] 8.585019f
C784 SWP[3] COMP_P 0.106335f
C785 CF[6] CF[0] 0.139154f
C786 SWP[7] SWP[2] 0.132136f
C787 SWP[5] SWP[9] 0.131001f
C788 CLK DOUT[3] 0.142459f
C789 SWP[3] DOUT[1] 0.013499f
C790 CF[8] COMP_N 0.062035f
C791 VSSD EN 37.9877f
C792 CF[4] SWP[4] 0.067118f
C793 COMP_P SWN[9] 0.062035f
C794 SWP[6] SWN[7] 0.062015f
C795 SWP[8] SWN[8] 0.070147f
C796 CF[9] SWN[4] 0.128503f
C797 SWP[2] SWN[5] 0.064209f
C798 SWP[4] SWN[6] 0.061493f
C799 SWP[9] SWN[7] 0.062015f
C800 CF[2] SWP[1] 0.096376f
C801 out_latch_0.FINAL CF[0] 0.067782f
C802 SWP[0] SWN[4] 0.0659f
C803 SWP[5] SWN[3] 0.065356f
C804 SWP[7] SWN[5] 0.064173f
C805 SWP[3] SWN[1] 0.065124f
C806 SWP[4] COMP_N 0.112004f
C807 CF[0] SWP[1] 0.072426f
C808 CF[4] SWN[4] 0.065885f
C809 SWN[3] SWN[7] 0.065736f
C810 SWN[1] SWN[9] 0.065208f
C811 VSSD auto_sampling_0.x11.D 0.311297f
C812 CF[3] SWP[8] 0.061924f
C813 SWN[2] SWN[8] 0.068035f
C814 SWN[4] SWN[6] 0.067463f
C815 auto_sampling_0.x22.A EN 0.147456f
C816 auto_sampling_0.x21.Q CLK 0.330595f
C817 cdac_ctrl_0.x1.X cdac_ctrl_0.x2.X 0.149159f
C818 CF[1] SWP[3] 0.071065f
C819 cdac_ctrl_0.x1.X CF[8] 0.03374f
C820 COMP_N SWN[4] 0.062143f
C821 CF[1] SWN[9] 0.07529f
C822 CF[3] SWN[2] 0.624398f
C823 VSSD CF[9] 6.09196f
C824 EN CLKSB 0.266704f
C825 VSSD SWP[0] 5.97717f
C826 CF[5] SWP[3] 0.071145f
C827 CF[0] DOUT[8] 0.0309f
C828 cdac_ctrl_0.x1.X SWP[4] 0.083633f
C829 VDDD CF[2] 1.21872f
C830 CF[5] SWN[9] 0.07529f
C831 VSSD CF[4] 4.93523f
C832 CF[2] SWN[0] 0.215004f
C833 VSSD SWN[6] 2.80751f
C834 CLKS CF[2] 0.183547f
C835 CF[6] SWP[5] 0.098919f
C836 VDDD CF[0] 1.30465f
C837 CF[0] SWN[0] 0.07764f
C838 CLKS CF[0] 0.153453f
C839 VSSD COMP_N 7.01361f
C840 EN DOUT[6] 0.317304f
C841 CF[6] SWN[7] 0.062043f
C842 EN DOUT[1] 0.318453f
C843 out_latch_0.FINAL SWP[5] 0.089103f
C844 CF[7] SWP[2] 0.06835f
C845 CF[7] SWP[7] 0.06276f
C846 auto_sampling_0.x24.A VDDD 0.839441f
C847 auto_sampling_0.x24.A CLKS 1.0051f
C848 SWP[1] SWP[5] 0.127098f
C849 CLKSB CF[9] 0.021519f
C850 CF[7] SWN[5] 0.125877f
C851 CF[8] SWP[6] 0.068175f
C852 CF[8] SWP[9] 0.076645f
C853 SWP[3] SWN[9] 0.075507f
C854 SWP[1] SWN[7] 0.062127f
C855 cdac_ctrl_0.x1.X VSSD 2.5607f
C856 cdac_ctrl_0.x2.X SWN[3] 0.077653f
C857 auto_sampling_0.x2.D EN 0.022065f
C858 CKO SWP[6] 0.107451f
C859 CKO DOUT[2] 0.195589f
C860 CF[8] SWN[3] 0.127707f
C861 CKO DOUT[5] 0.19774f
C862 CF[9] COMP_P 0.058086f
C863 CKO SWP[9] 0.070518f
C864 SWP[0] COMP_P 3.58746f
C865 SWP[4] SWP[6] 0.132285f
C866 SWP[2] SWP[8] 0.133168f
C867 DOUT[9] DOUT[4] 0.071825f
C868 SWP[2] DOUT[4] 0.016885f
C869 DOUT[0] DOUT[2] 0.058703f
C870 SWP[7] SWP[8] 8.21088f
C871 DOUT[7] DOUT[2] 0.050442f
C872 SWP[9] SWP[4] 0.130312f
C873 DOUT[5] DOUT[0] 0.058281f
C874 DOUT[3] DOUT[9] 0.071758f
C875 DOUT[5] DOUT[7] 0.051706f
C876 SWP[9] DOUT[7] 0.013729f
C877 CF[4] COMP_P 0.058086f
C878 COMP_P SWN[6] 0.062113f
C879 CF[9] SWN[1] 0.12732f
C880 SWP[8] SWN[5] 0.064173f
C881 SWP[4] SWN[3] 0.065356f
C882 CLK CF[2] 0.214219f
C883 VDDD SWP[5] 0.800498f
C884 SWP[6] SWN[4] 0.065851f
C885 SWP[0] SWN[1] 0.065124f
C886 SWP[2] SWN[2] 0.076273f
C887 SWP[7] SWN[2] 0.067874f
C888 SWP[9] SWN[4] 0.065851f
C889 SWP[5] SWN[0] 0.075119f
C890 CLKS SWP[5] 0.119526f
C891 COMP_P COMP_N 14.6546f
C892 VDDD SWN[7] 0.523563f
C893 CF[2] SWN[8] 0.061748f
C894 CF[4] SWN[1] 0.12732f
C895 CF[9] CF[1] 0.139852f
C896 SWN[0] SWN[7] 0.075232f
C897 SWN[2] SWN[5] 0.068495f
C898 SWN[3] SWN[4] 11.9787f
C899 SWN[1] SWN[6] 0.065338f
C900 CF[1] SWP[0] 0.104222f
C901 CLKS SWN[7] 0.019522f
C902 CF[0] SWN[8] 0.069113f
C903 COMP_N SWN[1] 0.062504f
C904 cdac_ctrl_0.x2.X CF[6] 0.074929f
C905 CF[2] CF[3] 13.2592f
C906 auto_sampling_0.x3.D EN 0.022065f
C907 CF[1] CF[4] 0.140692f
C908 CF[1] SWN[6] 0.061468f
C909 CF[8] CF[6] 0.130113f
C910 CF[9] CF[5] 0.140889f
C911 EN SWP[3] 0.083646f
C912 CF[5] SWP[0] 0.072959f
C913 VSSD SWP[6] 3.65574f
C914 VSSD DOUT[2] 3.07273f
C915 VSSD DOUT[5] 3.52092f
C916 CF[0] CF[3] 0.14365f
C917 VSSD SWP[9] 3.46966f
C918 CF[1] COMP_N 0.062035f
C919 SWN[9] VSUBS 16.62187f
C920 SWN[8] VSUBS 19.239046f
C921 SWN[7] VSUBS 21.13418f
C922 SWN[6] VSUBS 23.326672f
C923 SWN[5] VSUBS 24.334776f
C924 SWN[4] VSUBS 25.73887f
C925 SWN[3] VSUBS 27.637457f
C926 SWN[2] VSUBS 28.250862f
C927 SWN[1] VSUBS 31.536314f
C928 SWN[0] VSUBS 27.532963f
C929 COMP_N VSUBS 26.89369f
C930 COMP_P VSUBS 22.358158f
C931 DOUT[8] VSUBS 35.194984f
C932 SWP[8] VSUBS 10.736039f
C933 DOUT[6] VSUBS 33.385292f
C934 SWP[6] VSUBS 12.020971f
C935 DOUT[4] VSUBS 27.203848f
C936 SWP[4] VSUBS 14.228902f
C937 DOUT[2] VSUBS 26.695694f
C938 SWP[2] VSUBS 17.3826f
C939 DOUT[0] VSUBS 11.400654f
C940 SWP[0] VSUBS 18.106451f
C941 DOUT[9] VSUBS 29.805141f
C942 DOUT[7] VSUBS 34.965485f
C943 DOUT[5] VSUBS 29.957102f
C944 DOUT[3] VSUBS 27.15759f
C945 DOUT[1] VSUBS 25.599648f
C946 SWP[9] VSUBS 8.792482f
C947 SWP[7] VSUBS 12.98088f
C948 SWP[5] VSUBS 14.641512f
C949 SWP[3] VSUBS 15.891117f
C950 SWP[1] VSUBS 18.41134f
C951 CKO VSUBS 23.727255f
C952 CF[4] VSUBS 10.060575f
C953 CF[3] VSUBS 12.659018f
C954 CF[2] VSUBS 13.942185f
C955 CF[1] VSUBS 15.25297f
C956 CF[0] VSUBS 14.019162f
C957 CF[5] VSUBS 10.319805f
C958 CF[6] VSUBS 9.773911f
C959 CF[7] VSUBS 9.877414f
C960 CF[8] VSUBS 10.182673f
C961 CF[9] VSUBS 9.259317f
C962 CLKSB VSUBS 24.190775f
C963 CLKS VSUBS 26.954609f
C964 EN VSUBS 21.428263f
C965 CLK VSUBS 11.937539f
C966 VSSD VSUBS 53.26668f
C967 VDDD VSUBS 2.162678p
C968 cdac_ctrl_0.x2.X VSUBS 3.867246f
C969 cdac_ctrl_0.x1.X VSUBS 1.165286f
C970 out_latch_0.FINAL VSUBS 19.667854f
C971 auto_sampling_0.x24.A VSUBS 0.270258f
C972 auto_sampling_0.x23.A VSUBS 0.135663f
C973 auto_sampling_0.x21.D VSUBS 0.037498f
C974 auto_sampling_0.x16.D VSUBS 0.036085f
C975 auto_sampling_0.x15.D VSUBS 0.036085f
C976 auto_sampling_0.x14.D VSUBS 0.036085f
C977 auto_sampling_0.x22.A VSUBS 0.346459f
C978 auto_sampling_0.x12.D VSUBS 2.398725f
C979 auto_sampling_0.x11.Q VSUBS 0.040444f
C980 auto_sampling_0.x11.D VSUBS 0.038006f
C981 auto_sampling_0.x5.D VSUBS 0.036593f
C982 auto_sampling_0.x3.D VSUBS 0.036593f
C983 auto_sampling_0.x2.D VSUBS 0.036593f
C984 auto_sampling_0.x7.Q VSUBS 0.038006f
C985 auto_sampling_0.x21.Q VSUBS 2.790778f
C986 SWP[0].t5 VSUBS 0.028191f
C987 SWP[0].t4 VSUBS 0.031052f
C988 SWP[0].n0 VSUBS 0.088928f
C989 SWP[0].n1 VSUBS 10.8617f
C990 SWP[0].t2 VSUBS 0.022556f
C991 SWP[0].t3 VSUBS 0.022556f
C992 SWP[0].n2 VSUBS 0.045158f
C993 SWP[0].t0 VSUBS 0.014661f
C994 SWP[0].t1 VSUBS 0.014661f
C995 SWP[0].n4 VSUBS 0.029323f
C996 SWP[0].n5 VSUBS 0.039587f
C997 SWP[0].n6 VSUBS 0.032253f
C998 SWN[7].t1 VSUBS 0.015217f
C999 SWN[7].t0 VSUBS 0.015217f
C1000 SWN[7].n0 VSUBS 0.030435f
C1001 SWN[7].n1 VSUBS 0.036328f
C1002 SWN[7].t3 VSUBS 0.023411f
C1003 SWN[7].n2 VSUBS 0.01474f
C1004 SWN[7].t2 VSUBS 0.023411f
C1005 SWN[7].n3 VSUBS 0.046823f
C1006 SWN[7].n4 VSUBS 0.01474f
C1007 SWN[7].n5 VSUBS 0.056814f
C1008 SWN[3].t0 VSUBS 0.016376f
C1009 SWN[3].t1 VSUBS 0.016376f
C1010 SWN[3].n0 VSUBS 0.032753f
C1011 SWN[3].n1 VSUBS 0.039095f
C1012 SWN[3].t3 VSUBS 0.025195f
C1013 SWN[3].n2 VSUBS 0.015863f
C1014 SWN[3].t2 VSUBS 0.025195f
C1015 SWN[3].n3 VSUBS 0.050389f
C1016 SWN[3].n4 VSUBS 0.015863f
C1017 SWN[3].n5 VSUBS 0.060771f
C1018 DOUT[6].t2 VSUBS 0.028854f
C1019 DOUT[6].t3 VSUBS 0.028854f
C1020 DOUT[6].t0 VSUBS 0.018755f
C1021 DOUT[6].t1 VSUBS 0.018755f
C1022 DOUT[6].n0 VSUBS 0.03751f
C1023 DOUT[6].n1 VSUBS 0.05064f
C1024 DOUT[6].n2 VSUBS 0.018167f
C1025 DOUT[6].n3 VSUBS 0.057707f
C1026 DOUT[6].n4 VSUBS 0.056583f
C1027 SWN[8].t0 VSUBS 0.014635f
C1028 SWN[8].t1 VSUBS 0.014635f
C1029 SWN[8].n0 VSUBS 0.029271f
C1030 SWN[8].n1 VSUBS 0.034938f
C1031 SWN[8].t2 VSUBS 0.022516f
C1032 SWN[8].n2 VSUBS 0.014177f
C1033 SWN[8].t3 VSUBS 0.022516f
C1034 SWN[8].n3 VSUBS 0.045032f
C1035 SWN[8].n4 VSUBS 0.014177f
C1036 SWN[8].n5 VSUBS 0.054575f
C1037 CLKSB.t1 VSUBS 0.085247f
C1038 CLKSB.t0 VSUBS 0.056057f
C1039 CLKSB.n1 VSUBS 0.125716f
C1040 DOUT[4].t2 VSUBS 0.024779f
C1041 DOUT[4].t3 VSUBS 0.024779f
C1042 DOUT[4].t0 VSUBS 0.016106f
C1043 DOUT[4].t1 VSUBS 0.016106f
C1044 DOUT[4].n0 VSUBS 0.032213f
C1045 DOUT[4].n1 VSUBS 0.043489f
C1046 DOUT[4].n2 VSUBS 0.015601f
C1047 DOUT[4].n3 VSUBS 0.049558f
C1048 DOUT[4].n4 VSUBS 0.04863f
C1049 DOUT[7].t3 VSUBS 0.029144f
C1050 DOUT[7].t2 VSUBS 0.029144f
C1051 DOUT[7].t1 VSUBS 0.018944f
C1052 DOUT[7].t0 VSUBS 0.018944f
C1053 DOUT[7].n0 VSUBS 0.037888f
C1054 DOUT[7].n1 VSUBS 0.048673f
C1055 DOUT[7].n2 VSUBS 0.01835f
C1056 DOUT[7].n3 VSUBS 0.058288f
C1057 DOUT[7].n4 VSUBS 0.013763f
C1058 DOUT[7].n5 VSUBS 0.052318f
C1059 COMP_P.t3 VSUBS 0.046729f
C1060 COMP_P.t2 VSUBS 0.029138f
C1061 COMP_P.t5 VSUBS 0.044596f
C1062 COMP_P.t4 VSUBS 0.026664f
C1063 COMP_P.n0 VSUBS 0.055105f
C1064 COMP_P.t1 VSUBS 0.044596f
C1065 COMP_P.t0 VSUBS 0.026664f
C1066 COMP_P.n1 VSUBS 0.062683f
C1067 COMP_P.n2 VSUBS 0.023576f
C1068 COMP_P.n3 VSUBS 0.017672f
C1069 COMP_P.n4 VSUBS 0.015593f
C1070 COMP_P.n5 VSUBS 0.019366f
C1071 COMP_P.n6 VSUBS 0.084594f
C1072 COMP_P.n7 VSUBS 0.015593f
C1073 COMP_P.n8 VSUBS 0.018494f
C1074 COMP_P.n9 VSUBS 7.70172f
C1075 SWP[2].t5 VSUBS 0.029202f
C1076 SWP[2].t4 VSUBS 0.032166f
C1077 SWP[2].n0 VSUBS 0.092117f
C1078 SWP[2].n1 VSUBS 10.4396f
C1079 SWP[2].t2 VSUBS 0.023365f
C1080 SWP[2].t3 VSUBS 0.023365f
C1081 SWP[2].n2 VSUBS 0.046778f
C1082 SWP[2].t0 VSUBS 0.015187f
C1083 SWP[2].t1 VSUBS 0.015187f
C1084 SWP[2].n4 VSUBS 0.030374f
C1085 SWP[2].n5 VSUBS 0.041007f
C1086 SWP[2].n6 VSUBS 0.033605f
C1087 SWP[3].t5 VSUBS 0.027439f
C1088 SWP[3].t4 VSUBS 0.030205f
C1089 SWP[3].n0 VSUBS 0.086794f
C1090 SWP[3].n1 VSUBS 0.187773f
C1091 SWP[3].n2 VSUBS 9.11291f
C1092 SWP[3].t2 VSUBS 0.021846f
C1093 SWP[3].t3 VSUBS 0.021846f
C1094 SWP[3].n3 VSUBS 0.043738f
C1095 SWP[3].t0 VSUBS 0.0142f
C1096 SWP[3].t1 VSUBS 0.0142f
C1097 SWP[3].n5 VSUBS 0.0284f
C1098 SWP[3].n6 VSUBS 0.038342f
C1099 SWP[3].n7 VSUBS 0.03136f
C1100 CF[0].t6 VSUBS 0.030873f
C1101 CF[0].t10 VSUBS 0.020655f
C1102 CF[0].n0 VSUBS 0.056416f
C1103 CF[0].n2 VSUBS 0.037059f
C1104 CF[0].t12 VSUBS 0.020655f
C1105 CF[0].t7 VSUBS 0.030873f
C1106 CF[0].n3 VSUBS 0.056557f
C1107 CF[0].n4 VSUBS 0.038671f
C1108 CF[0].n5 VSUBS 0.335907f
C1109 CF[0].t4 VSUBS 0.019745f
C1110 CF[0].t8 VSUBS 0.031665f
C1111 CF[0].n6 VSUBS 0.057323f
C1112 CF[0].t11 VSUBS 0.018068f
C1113 CF[0].t13 VSUBS 0.030219f
C1114 CF[0].t5 VSUBS 0.018068f
C1115 CF[0].t9 VSUBS 0.030219f
C1116 CF[0].n7 VSUBS 0.042476f
C1117 CF[0].n8 VSUBS 0.012961f
C1118 CF[0].n9 VSUBS 0.015976f
C1119 CF[0].n10 VSUBS 0.037341f
C1120 CF[0].n11 VSUBS 0.013123f
C1121 CF[0].n12 VSUBS 0.012961f
C1122 CF[0].n13 VSUBS 0.02104f
C1123 CF[0].t2 VSUBS 0.019019f
C1124 CF[0].t3 VSUBS 0.019019f
C1125 CF[0].t0 VSUBS 0.012362f
C1126 CF[0].t1 VSUBS 0.012362f
C1127 CF[0].n14 VSUBS 0.024725f
C1128 CF[0].n15 VSUBS 0.031764f
C1129 CF[0].n16 VSUBS 0.011975f
C1130 CF[0].n17 VSUBS 0.038038f
C1131 CF[0].n19 VSUBS 0.013355f
C1132 CF[0].n20 VSUBS 0.261496f
C1133 CF[0].n21 VSUBS 15.410099f
C1134 SWN[4].t0 VSUBS 0.015956f
C1135 SWN[4].t1 VSUBS 0.015956f
C1136 SWN[4].n0 VSUBS 0.031912f
C1137 SWN[4].n1 VSUBS 0.038091f
C1138 SWN[4].t2 VSUBS 0.024548f
C1139 SWN[4].n2 VSUBS 0.015456f
C1140 SWN[4].t3 VSUBS 0.024548f
C1141 SWN[4].n3 VSUBS 0.049096f
C1142 SWN[4].n4 VSUBS 0.015456f
C1143 SWN[4].n5 VSUBS 0.0595f
C1144 SWN[2].t0 VSUBS 0.016023f
C1145 SWN[2].t1 VSUBS 0.016023f
C1146 SWN[2].n0 VSUBS 0.032046f
C1147 SWN[2].n1 VSUBS 0.03825f
C1148 SWN[2].t3 VSUBS 0.02465f
C1149 SWN[2].n2 VSUBS 0.015521f
C1150 SWN[2].t2 VSUBS 0.02465f
C1151 SWN[2].n3 VSUBS 0.049301f
C1152 SWN[2].n4 VSUBS 0.015521f
C1153 SWN[2].n5 VSUBS 0.059422f
C1154 auto_sampling_0.x12.D.t0 VSUBS 0.037889f
C1155 auto_sampling_0.x12.D.t1 VSUBS 0.057618f
C1156 auto_sampling_0.x12.D.t2 VSUBS 0.019246f
C1157 auto_sampling_0.x12.D.t3 VSUBS 0.021187f
C1158 auto_sampling_0.x12.D.n0 VSUBS 0.06088f
C1159 auto_sampling_0.x12.D.n1 VSUBS 3.42496f
C1160 SWP[9].t4 VSUBS 0.023657f
C1161 SWP[9].t5 VSUBS 0.026042f
C1162 SWP[9].n0 VSUBS 0.07483f
C1163 SWP[9].n1 VSUBS 0.161191f
C1164 SWP[9].t3 VSUBS 0.018835f
C1165 SWP[9].t2 VSUBS 0.018835f
C1166 SWP[9].n2 VSUBS 0.037709f
C1167 SWP[9].t1 VSUBS 0.012243f
C1168 SWP[9].t0 VSUBS 0.012243f
C1169 SWP[9].n4 VSUBS 0.024485f
C1170 SWP[9].n5 VSUBS 0.033057f
C1171 SWP[9].n6 VSUBS 0.027143f
C1172 SWP[9].n7 VSUBS 6.98011f
C1173 SWP[9].n8 VSUBS 1.39271f
C1174 SWP[6].t4 VSUBS 0.026304f
C1175 SWP[6].t5 VSUBS 0.028974f
C1176 SWP[6].n0 VSUBS 0.082977f
C1177 SWP[6].n1 VSUBS 1.11681f
C1178 SWP[6].n2 VSUBS 8.08604f
C1179 SWP[6].t2 VSUBS 0.021046f
C1180 SWP[6].t3 VSUBS 0.021046f
C1181 SWP[6].n3 VSUBS 0.042136f
C1182 SWP[6].t0 VSUBS 0.01368f
C1183 SWP[6].t1 VSUBS 0.01368f
C1184 SWP[6].n5 VSUBS 0.02736f
C1185 SWP[6].n6 VSUBS 0.036938f
C1186 SWP[6].n7 VSUBS 0.030212f
C1187 DOUT[3].t3 VSUBS 0.025116f
C1188 DOUT[3].t2 VSUBS 0.025116f
C1189 DOUT[3].t1 VSUBS 0.016325f
C1190 DOUT[3].t0 VSUBS 0.016325f
C1191 DOUT[3].n0 VSUBS 0.03265f
C1192 DOUT[3].n1 VSUBS 0.041945f
C1193 DOUT[3].n2 VSUBS 0.015814f
C1194 DOUT[3].n3 VSUBS 0.050231f
C1195 DOUT[3].n4 VSUBS 0.01186f
C1196 DOUT[3].n5 VSUBS 0.045475f
C1197 SWP[5].t5 VSUBS 0.027442f
C1198 SWP[5].t4 VSUBS 0.030208f
C1199 SWP[5].n0 VSUBS 0.086804f
C1200 SWP[5].n1 VSUBS 0.186906f
C1201 SWP[5].n2 VSUBS 8.313429f
C1202 SWP[5].t2 VSUBS 0.021849f
C1203 SWP[5].t3 VSUBS 0.021849f
C1204 SWP[5].n3 VSUBS 0.043742f
C1205 SWP[5].t0 VSUBS 0.014202f
C1206 SWP[5].t1 VSUBS 0.014202f
C1207 SWP[5].n5 VSUBS 0.028403f
C1208 SWP[5].n6 VSUBS 0.038346f
C1209 SWP[5].n7 VSUBS 0.031547f
C1210 CF[2].t7 VSUBS 0.040655f
C1211 CF[2].t9 VSUBS 0.0272f
C1212 CF[2].n0 VSUBS 0.074291f
C1213 CF[2].n2 VSUBS 0.048801f
C1214 CF[2].t4 VSUBS 0.0272f
C1215 CF[2].t5 VSUBS 0.040655f
C1216 CF[2].n3 VSUBS 0.074478f
C1217 CF[2].n4 VSUBS 0.050924f
C1218 CF[2].n5 VSUBS 0.439652f
C1219 CF[2].t3 VSUBS 0.025046f
C1220 CF[2].t2 VSUBS 0.025046f
C1221 CF[2].t1 VSUBS 0.01628f
C1222 CF[2].t0 VSUBS 0.01628f
C1223 CF[2].n6 VSUBS 0.032559f
C1224 CF[2].n7 VSUBS 0.041828f
C1225 CF[2].n8 VSUBS 0.015769f
C1226 CF[2].n9 VSUBS 0.050091f
C1227 CF[2].n10 VSUBS 0.011827f
C1228 CF[2].n11 VSUBS 0.02511f
C1229 CF[2].t8 VSUBS 0.031302f
C1230 CF[2].t6 VSUBS 0.03448f
C1231 CF[2].n12 VSUBS 0.098744f
C1232 CF[2].n13 VSUBS 0.414451f
C1233 CF[2].n14 VSUBS 18.5024f
C1234 COMP_N.t2 VSUBS 0.02258f
C1235 COMP_N.t4 VSUBS 0.036211f
C1236 COMP_N.t3 VSUBS 0.020662f
C1237 COMP_N.t0 VSUBS 0.034558f
C1238 COMP_N.n0 VSUBS 0.042702f
C1239 COMP_N.t1 VSUBS 0.020662f
C1240 COMP_N.t5 VSUBS 0.034558f
C1241 COMP_N.n1 VSUBS 0.048574f
C1242 COMP_N.n2 VSUBS 0.01827f
C1243 COMP_N.n3 VSUBS 0.013694f
C1244 COMP_N.n4 VSUBS 0.012083f
C1245 COMP_N.n5 VSUBS 0.015007f
C1246 COMP_N.n6 VSUBS 0.065553f
C1247 COMP_N.n7 VSUBS 0.012083f
C1248 COMP_N.n8 VSUBS 0.014724f
C1249 CF[6].t4 VSUBS 0.03711f
C1250 CF[6].t5 VSUBS 0.024829f
C1251 CF[6].n0 VSUBS 0.067813f
C1252 CF[6].n2 VSUBS 0.044546f
C1253 CF[6].t7 VSUBS 0.024829f
C1254 CF[6].t9 VSUBS 0.03711f
C1255 CF[6].n3 VSUBS 0.067983f
C1256 CF[6].n4 VSUBS 0.046483f
C1257 CF[6].n5 VSUBS 0.401315f
C1258 CF[6].t6 VSUBS 0.028714f
C1259 CF[6].t8 VSUBS 0.031609f
C1260 CF[6].n6 VSUBS 0.090828f
C1261 CF[6].n7 VSUBS 0.178888f
C1262 CF[6].t2 VSUBS 0.022862f
C1263 CF[6].t3 VSUBS 0.022862f
C1264 CF[6].t0 VSUBS 0.01486f
C1265 CF[6].t1 VSUBS 0.01486f
C1266 CF[6].n8 VSUBS 0.02972f
C1267 CF[6].n9 VSUBS 0.040124f
C1268 CF[6].n10 VSUBS 0.014394f
C1269 CF[6].n11 VSUBS 0.045723f
C1270 CF[6].n12 VSUBS 0.028354f
C1271 CF[6].n13 VSUBS 0.358367f
C1272 CF[6].n14 VSUBS 14.4044f
C1273 SWN[0].t0 VSUBS 0.014309f
C1274 SWN[0].t1 VSUBS 0.014309f
C1275 SWN[0].n0 VSUBS 0.028618f
C1276 SWN[0].n1 VSUBS 0.034159f
C1277 SWN[0].t2 VSUBS 0.022014f
C1278 SWN[0].n2 VSUBS 0.013861f
C1279 SWN[0].t3 VSUBS 0.022014f
C1280 SWN[0].n3 VSUBS 0.044028f
C1281 SWN[0].n4 VSUBS 0.013861f
C1282 SWN[0].n5 VSUBS 0.052875f
C1283 DOUT[1].t2 VSUBS 0.025103f
C1284 DOUT[1].t3 VSUBS 0.025103f
C1285 DOUT[1].t1 VSUBS 0.016317f
C1286 DOUT[1].t0 VSUBS 0.016317f
C1287 DOUT[1].n0 VSUBS 0.032634f
C1288 DOUT[1].n1 VSUBS 0.041925f
C1289 DOUT[1].n2 VSUBS 0.015806f
C1290 DOUT[1].n3 VSUBS 0.050207f
C1291 DOUT[1].n4 VSUBS 0.011854f
C1292 DOUT[1].n5 VSUBS 0.045322f
C1293 CF[1].t6 VSUBS 0.041687f
C1294 CF[1].t9 VSUBS 0.027891f
C1295 CF[1].n0 VSUBS 0.076177f
C1296 CF[1].n2 VSUBS 0.05004f
C1297 CF[1].t5 VSUBS 0.027891f
C1298 CF[1].t8 VSUBS 0.041687f
C1299 CF[1].n3 VSUBS 0.076368f
C1300 CF[1].n4 VSUBS 0.052217f
C1301 CF[1].n5 VSUBS 0.450261f
C1302 CF[1].t2 VSUBS 0.025681f
C1303 CF[1].t3 VSUBS 0.025681f
C1304 CF[1].t1 VSUBS 0.016693f
C1305 CF[1].t0 VSUBS 0.016693f
C1306 CF[1].n6 VSUBS 0.033386f
C1307 CF[1].n7 VSUBS 0.04289f
C1308 CF[1].n8 VSUBS 0.01617f
C1309 CF[1].n9 VSUBS 0.051362f
C1310 CF[1].n10 VSUBS 0.012127f
C1311 CF[1].n11 VSUBS 0.025747f
C1312 CF[1].t4 VSUBS 0.032097f
C1313 CF[1].t7 VSUBS 0.035355f
C1314 CF[1].n12 VSUBS 0.10125f
C1315 CF[1].n13 VSUBS 0.422498f
C1316 CF[1].n14 VSUBS 19.9386f
C1317 SWN[6].t0 VSUBS 0.015943f
C1318 SWN[6].t1 VSUBS 0.015943f
C1319 SWN[6].n0 VSUBS 0.031886f
C1320 SWN[6].n1 VSUBS 0.038061f
C1321 SWN[6].t2 VSUBS 0.024528f
C1322 SWN[6].n2 VSUBS 0.015444f
C1323 SWN[6].t3 VSUBS 0.024528f
C1324 SWN[6].n3 VSUBS 0.049056f
C1325 SWN[6].n4 VSUBS 0.015444f
C1326 SWN[6].n5 VSUBS 0.059452f
C1327 DOUT[2].t3 VSUBS 0.025708f
C1328 DOUT[2].t2 VSUBS 0.025708f
C1329 DOUT[2].t0 VSUBS 0.01671f
C1330 DOUT[2].t1 VSUBS 0.01671f
C1331 DOUT[2].n0 VSUBS 0.03342f
C1332 DOUT[2].n1 VSUBS 0.045119f
C1333 DOUT[2].n2 VSUBS 0.016186f
C1334 DOUT[2].n3 VSUBS 0.051416f
C1335 DOUT[2].n4 VSUBS 0.050286f
C1336 DOUT[8].t3 VSUBS 0.029043f
C1337 DOUT[8].t2 VSUBS 0.029043f
C1338 DOUT[8].t1 VSUBS 0.018878f
C1339 DOUT[8].t0 VSUBS 0.018878f
C1340 DOUT[8].n0 VSUBS 0.037755f
C1341 DOUT[8].n1 VSUBS 0.050972f
C1342 DOUT[8].n2 VSUBS 0.018286f
C1343 DOUT[8].n3 VSUBS 0.058085f
C1344 DOUT[8].n4 VSUBS 0.056998f
C1345 CF[7].t8 VSUBS 0.037065f
C1346 CF[7].t4 VSUBS 0.024798f
C1347 CF[7].n0 VSUBS 0.067731f
C1348 CF[7].n2 VSUBS 0.044491f
C1349 CF[7].t6 VSUBS 0.024798f
C1350 CF[7].t7 VSUBS 0.037065f
C1351 CF[7].n3 VSUBS 0.0679f
C1352 CF[7].n4 VSUBS 0.046427f
C1353 CF[7].n5 VSUBS 0.402787f
C1354 CF[7].t5 VSUBS 0.028679f
C1355 CF[7].t9 VSUBS 0.03157f
C1356 CF[7].n6 VSUBS 0.090717f
C1357 CF[7].n7 VSUBS 0.17867f
C1358 CF[7].t3 VSUBS 0.022834f
C1359 CF[7].t2 VSUBS 0.022834f
C1360 CF[7].t1 VSUBS 0.014842f
C1361 CF[7].t0 VSUBS 0.014842f
C1362 CF[7].n8 VSUBS 0.029684f
C1363 CF[7].n9 VSUBS 0.040075f
C1364 CF[7].n10 VSUBS 0.014377f
C1365 CF[7].n11 VSUBS 0.045667f
C1366 CF[7].n12 VSUBS 0.02832f
C1367 CF[7].n13 VSUBS 0.360568f
C1368 CF[7].n14 VSUBS 14.316f
C1369 SWP[1].t5 VSUBS 0.031381f
C1370 SWP[1].t4 VSUBS 0.034545f
C1371 SWP[1].n0 VSUBS 0.099264f
C1372 SWP[1].n1 VSUBS 0.214821f
C1373 SWP[1].n2 VSUBS 1.21344f
C1374 SWP[1].n3 VSUBS 11.3398f
C1375 SWP[1].t2 VSUBS 0.024985f
C1376 SWP[1].t3 VSUBS 0.024985f
C1377 SWP[1].n4 VSUBS 0.050022f
C1378 SWP[1].t0 VSUBS 0.01624f
C1379 SWP[1].t1 VSUBS 0.01624f
C1380 SWP[1].n6 VSUBS 0.032481f
C1381 SWP[1].n7 VSUBS 0.043851f
C1382 SWP[1].n8 VSUBS 0.035866f
C1383 DOUT[9].t3 VSUBS 0.02248f
C1384 DOUT[9].t2 VSUBS 0.02248f
C1385 DOUT[9].t1 VSUBS 0.014612f
C1386 DOUT[9].t0 VSUBS 0.014612f
C1387 DOUT[9].n0 VSUBS 0.029224f
C1388 DOUT[9].n1 VSUBS 0.037544f
C1389 DOUT[9].n2 VSUBS 0.014154f
C1390 DOUT[9].n3 VSUBS 0.044961f
C1391 DOUT[9].n4 VSUBS 0.010616f
C1392 DOUT[9].n5 VSUBS 0.040432f
C1393 SWN[9].t1 VSUBS 0.013344f
C1394 SWN[9].t0 VSUBS 0.013344f
C1395 SWN[9].n0 VSUBS 0.026689f
C1396 SWN[9].n1 VSUBS 0.031856f
C1397 SWN[9].t2 VSUBS 0.02053f
C1398 SWN[9].n2 VSUBS 0.012926f
C1399 SWN[9].t3 VSUBS 0.02053f
C1400 SWN[9].n3 VSUBS 0.04106f
C1401 SWN[9].n4 VSUBS 0.012926f
C1402 SWN[9].n5 VSUBS 0.049639f
C1403 cdac_ctrl_0.x1.X.t0 VSUBS 0.022994f
C1404 cdac_ctrl_0.x1.X.t1 VSUBS 0.022994f
C1405 cdac_ctrl_0.x1.X.n0 VSUBS 0.048313f
C1406 cdac_ctrl_0.x1.X.t6 VSUBS 0.022994f
C1407 cdac_ctrl_0.x1.X.t7 VSUBS 0.022994f
C1408 cdac_ctrl_0.x1.X.n1 VSUBS 0.048313f
C1409 cdac_ctrl_0.x1.X.t4 VSUBS 0.022994f
C1410 cdac_ctrl_0.x1.X.t5 VSUBS 0.022994f
C1411 cdac_ctrl_0.x1.X.n2 VSUBS 0.068982f
C1412 cdac_ctrl_0.x1.X.n3 VSUBS 0.180042f
C1413 cdac_ctrl_0.x1.X.n4 VSUBS 0.107706f
C1414 cdac_ctrl_0.x1.X.t26 VSUBS 0.044432f
C1415 cdac_ctrl_0.x1.X.t30 VSUBS 0.048911f
C1416 cdac_ctrl_0.x1.X.n5 VSUBS 0.140546f
C1417 cdac_ctrl_0.x1.X.n6 VSUBS 0.357279f
C1418 cdac_ctrl_0.x1.X.t23 VSUBS 0.044432f
C1419 cdac_ctrl_0.x1.X.t18 VSUBS 0.048911f
C1420 cdac_ctrl_0.x1.X.n7 VSUBS 0.140546f
C1421 cdac_ctrl_0.x1.X.n8 VSUBS 0.262654f
C1422 cdac_ctrl_0.x1.X.n9 VSUBS 1.34877f
C1423 cdac_ctrl_0.x1.X.t34 VSUBS 0.044432f
C1424 cdac_ctrl_0.x1.X.t27 VSUBS 0.048911f
C1425 cdac_ctrl_0.x1.X.n10 VSUBS 0.140546f
C1426 cdac_ctrl_0.x1.X.n11 VSUBS 0.2628f
C1427 cdac_ctrl_0.x1.X.n12 VSUBS 0.930269f
C1428 cdac_ctrl_0.x1.X.t19 VSUBS 0.044432f
C1429 cdac_ctrl_0.x1.X.t24 VSUBS 0.048911f
C1430 cdac_ctrl_0.x1.X.n13 VSUBS 0.140546f
C1431 cdac_ctrl_0.x1.X.n14 VSUBS 0.2628f
C1432 cdac_ctrl_0.x1.X.n15 VSUBS 0.930269f
C1433 cdac_ctrl_0.x1.X.t20 VSUBS 0.044432f
C1434 cdac_ctrl_0.x1.X.t31 VSUBS 0.048911f
C1435 cdac_ctrl_0.x1.X.n16 VSUBS 0.140546f
C1436 cdac_ctrl_0.x1.X.n17 VSUBS 0.262654f
C1437 cdac_ctrl_0.x1.X.n18 VSUBS 0.930402f
C1438 cdac_ctrl_0.x1.X.t25 VSUBS 0.044432f
C1439 cdac_ctrl_0.x1.X.t21 VSUBS 0.048911f
C1440 cdac_ctrl_0.x1.X.n19 VSUBS 0.140546f
C1441 cdac_ctrl_0.x1.X.n20 VSUBS 0.262654f
C1442 cdac_ctrl_0.x1.X.n21 VSUBS 0.930402f
C1443 cdac_ctrl_0.x1.X.t17 VSUBS 0.044432f
C1444 cdac_ctrl_0.x1.X.t16 VSUBS 0.048911f
C1445 cdac_ctrl_0.x1.X.n22 VSUBS 0.140546f
C1446 cdac_ctrl_0.x1.X.n23 VSUBS 0.262654f
C1447 cdac_ctrl_0.x1.X.n24 VSUBS 0.930402f
C1448 cdac_ctrl_0.x1.X.t35 VSUBS 0.044432f
C1449 cdac_ctrl_0.x1.X.t33 VSUBS 0.048911f
C1450 cdac_ctrl_0.x1.X.n25 VSUBS 0.140546f
C1451 cdac_ctrl_0.x1.X.n26 VSUBS 0.262654f
C1452 cdac_ctrl_0.x1.X.n27 VSUBS 0.930402f
C1453 cdac_ctrl_0.x1.X.t32 VSUBS 0.044432f
C1454 cdac_ctrl_0.x1.X.t29 VSUBS 0.048911f
C1455 cdac_ctrl_0.x1.X.n28 VSUBS 0.140546f
C1456 cdac_ctrl_0.x1.X.n29 VSUBS 0.262654f
C1457 cdac_ctrl_0.x1.X.n30 VSUBS 0.930402f
C1458 cdac_ctrl_0.x1.X.t28 VSUBS 0.044432f
C1459 cdac_ctrl_0.x1.X.t22 VSUBS 0.048911f
C1460 cdac_ctrl_0.x1.X.n31 VSUBS 0.140546f
C1461 cdac_ctrl_0.x1.X.n32 VSUBS 0.262654f
C1462 cdac_ctrl_0.x1.X.n33 VSUBS 0.774864f
C1463 cdac_ctrl_0.x1.X.t10 VSUBS 0.035376f
C1464 cdac_ctrl_0.x1.X.t11 VSUBS 0.035376f
C1465 cdac_ctrl_0.x1.X.n34 VSUBS 0.070779f
C1466 cdac_ctrl_0.x1.X.n35 VSUBS 0.040461f
C1467 cdac_ctrl_0.x1.X.t8 VSUBS 0.035376f
C1468 cdac_ctrl_0.x1.X.t9 VSUBS 0.035376f
C1469 cdac_ctrl_0.x1.X.n36 VSUBS 0.075444f
C1470 cdac_ctrl_0.x1.X.t12 VSUBS 0.035376f
C1471 cdac_ctrl_0.x1.X.t13 VSUBS 0.035376f
C1472 cdac_ctrl_0.x1.X.n37 VSUBS 0.095016f
C1473 cdac_ctrl_0.x1.X.t14 VSUBS 0.035376f
C1474 cdac_ctrl_0.x1.X.t15 VSUBS 0.035376f
C1475 cdac_ctrl_0.x1.X.n38 VSUBS 0.075444f
C1476 cdac_ctrl_0.x1.X.n39 VSUBS 0.242333f
C1477 cdac_ctrl_0.x1.X.n40 VSUBS 0.138302f
C1478 cdac_ctrl_0.x1.X.n41 VSUBS 0.065904f
C1479 cdac_ctrl_0.x1.X.n42 VSUBS 0.052552f
C1480 cdac_ctrl_0.x1.X.t2 VSUBS 0.022994f
C1481 cdac_ctrl_0.x1.X.t3 VSUBS 0.022994f
C1482 cdac_ctrl_0.x1.X.n43 VSUBS 0.048633f
C1483 SWP[7].t5 VSUBS 0.026474f
C1484 SWP[7].t4 VSUBS 0.029143f
C1485 SWP[7].n0 VSUBS 0.083743f
C1486 SWP[7].n1 VSUBS 0.180337f
C1487 SWP[7].n2 VSUBS 7.26299f
C1488 SWP[7].t2 VSUBS 0.021078f
C1489 SWP[7].t3 VSUBS 0.021078f
C1490 SWP[7].n3 VSUBS 0.0422f
C1491 SWP[7].t0 VSUBS 0.013701f
C1492 SWP[7].t1 VSUBS 0.013701f
C1493 SWP[7].n5 VSUBS 0.027402f
C1494 SWP[7].n6 VSUBS 0.036994f
C1495 SWP[7].n7 VSUBS 0.030375f
C1496 CKO.t1 VSUBS 0.050079f
C1497 CKO.n0 VSUBS 0.046875f
C1498 CKO.n1 VSUBS 0.015479f
C1499 CKO.t0 VSUBS 0.03518f
C1500 CKO.n2 VSUBS 0.10708f
C1501 CKO.n3 VSUBS 0.023413f
C1502 CKO.t3 VSUBS 0.127897f
C1503 CKO.n4 VSUBS 0.019566f
C1504 CKO.t2 VSUBS 0.050079f
C1505 CKO.n5 VSUBS 0.057729f
C1506 CKO.n6 VSUBS 0.016572f
C1507 CKO.n7 VSUBS 0.021893f
C1508 CKO.n8 VSUBS 0.201803f
C1509 CKO.t12 VSUBS 0.032805f
C1510 CKO.t18 VSUBS 0.021948f
C1511 CKO.n9 VSUBS 0.059947f
C1512 CKO.n10 VSUBS 0.017814f
C1513 CKO.n11 VSUBS 0.424933f
C1514 CKO.t20 VSUBS 0.032805f
C1515 CKO.t22 VSUBS 0.021948f
C1516 CKO.n12 VSUBS 0.059947f
C1517 CKO.n13 VSUBS 0.017814f
C1518 CKO.n14 VSUBS 0.750505f
C1519 CKO.t7 VSUBS 0.032805f
C1520 CKO.t15 VSUBS 0.021948f
C1521 CKO.n15 VSUBS 0.059947f
C1522 CKO.n16 VSUBS 0.017814f
C1523 CKO.n17 VSUBS 0.591523f
C1524 CKO.t14 VSUBS 0.032805f
C1525 CKO.t19 VSUBS 0.021948f
C1526 CKO.n18 VSUBS 0.059947f
C1527 CKO.n19 VSUBS 0.017814f
C1528 CKO.t6 VSUBS 0.032805f
C1529 CKO.t11 VSUBS 0.021948f
C1530 CKO.n20 VSUBS 0.059947f
C1531 CKO.n21 VSUBS 0.017814f
C1532 CKO.n22 VSUBS 0.850694f
C1533 CKO.n23 VSUBS 0.444397f
C1534 CKO.t21 VSUBS 0.021948f
C1535 CKO.t23 VSUBS 0.032805f
C1536 CKO.n24 VSUBS 0.060631f
C1537 CKO.n25 VSUBS 0.12969f
C1538 CKO.t5 VSUBS 0.021948f
C1539 CKO.t9 VSUBS 0.032805f
C1540 CKO.n26 VSUBS 0.060631f
C1541 CKO.n27 VSUBS 0.026953f
C1542 CKO.n28 VSUBS 0.904004f
C1543 CKO.n29 VSUBS 0.444401f
C1544 CKO.t4 VSUBS 0.021948f
C1545 CKO.t8 VSUBS 0.032805f
C1546 CKO.n30 VSUBS 0.060631f
C1547 CKO.n31 VSUBS 0.026953f
C1548 CKO.n32 VSUBS 0.534278f
C1549 CKO.t10 VSUBS 0.021948f
C1550 CKO.t16 VSUBS 0.032805f
C1551 CKO.n33 VSUBS 0.060631f
C1552 CKO.n34 VSUBS 0.026953f
C1553 CKO.n35 VSUBS 0.750505f
C1554 CKO.t13 VSUBS 0.021948f
C1555 CKO.t17 VSUBS 0.032805f
C1556 CKO.n36 VSUBS 0.060631f
C1557 CKO.n37 VSUBS 0.026953f
C1558 CKO.n38 VSUBS 0.462439f
C1559 SWN[5].t0 VSUBS 0.015826f
C1560 SWN[5].t1 VSUBS 0.015826f
C1561 SWN[5].n0 VSUBS 0.031653f
C1562 SWN[5].n1 VSUBS 0.037782f
C1563 SWN[5].t2 VSUBS 0.024348f
C1564 SWN[5].n2 VSUBS 0.01533f
C1565 SWN[5].t3 VSUBS 0.024348f
C1566 SWN[5].n3 VSUBS 0.048697f
C1567 SWN[5].n4 VSUBS 0.01533f
C1568 SWN[5].n5 VSUBS 0.059016f
C1569 SWP[8].t4 VSUBS 0.026341f
C1570 SWP[8].t5 VSUBS 0.029015f
C1571 SWP[8].n0 VSUBS 0.083094f
C1572 SWP[8].n1 VSUBS 1.17334f
C1573 SWP[8].n2 VSUBS 7.50078f
C1574 SWP[8].t3 VSUBS 0.021076f
C1575 SWP[8].t1 VSUBS 0.021076f
C1576 SWP[8].n3 VSUBS 0.042195f
C1577 SWP[8].t2 VSUBS 0.013699f
C1578 SWP[8].t0 VSUBS 0.013699f
C1579 SWP[8].n5 VSUBS 0.027399f
C1580 SWP[8].n6 VSUBS 0.03699f
C1581 SWP[8].n7 VSUBS 0.030254f
C1582 SWN[1].t1 VSUBS 0.017155f
C1583 SWN[1].t0 VSUBS 0.017155f
C1584 SWN[1].n0 VSUBS 0.03431f
C1585 SWN[1].n1 VSUBS 0.040953f
C1586 SWN[1].t2 VSUBS 0.026392f
C1587 SWN[1].n2 VSUBS 0.016617f
C1588 SWN[1].t3 VSUBS 0.026392f
C1589 SWN[1].n3 VSUBS 0.052785f
C1590 SWN[1].n4 VSUBS 0.016617f
C1591 SWN[1].n5 VSUBS 0.06397f
C1592 auto_sampling_0.x21.Q.n1 VSUBS 0.010663f
C1593 auto_sampling_0.x21.Q.n2 VSUBS 0.012164f
C1594 auto_sampling_0.x21.Q.n4 VSUBS 0.02379f
C1595 auto_sampling_0.x21.Q.n5 VSUBS 1.3832f
C1596 DOUT[5].t3 VSUBS 0.026244f
C1597 DOUT[5].t2 VSUBS 0.026244f
C1598 DOUT[5].t1 VSUBS 0.017059f
C1599 DOUT[5].t0 VSUBS 0.017059f
C1600 DOUT[5].n0 VSUBS 0.034118f
C1601 DOUT[5].n1 VSUBS 0.04383f
C1602 DOUT[5].n2 VSUBS 0.016524f
C1603 DOUT[5].n3 VSUBS 0.052489f
C1604 DOUT[5].n4 VSUBS 0.012393f
C1605 DOUT[5].n5 VSUBS 0.047382f
C1606 SWP[4].t5 VSUBS 0.02799f
C1607 SWP[4].t4 VSUBS 0.030831f
C1608 SWP[4].n0 VSUBS 0.088294f
C1609 SWP[4].n1 VSUBS 1.10548f
C1610 SWP[4].n2 VSUBS 9.28035f
C1611 SWP[4].t2 VSUBS 0.022395f
C1612 SWP[4].t3 VSUBS 0.022395f
C1613 SWP[4].n3 VSUBS 0.044836f
C1614 SWP[4].t0 VSUBS 0.014557f
C1615 SWP[4].t1 VSUBS 0.014557f
C1616 SWP[4].n5 VSUBS 0.029114f
C1617 SWP[4].n6 VSUBS 0.039305f
C1618 SWP[4].n7 VSUBS 0.032148f
C1619 CF[9].t5 VSUBS 0.033044f
C1620 CF[9].t7 VSUBS 0.022108f
C1621 CF[9].n0 VSUBS 0.060382f
C1622 CF[9].n2 VSUBS 0.039665f
C1623 CF[9].t9 VSUBS 0.022108f
C1624 CF[9].t4 VSUBS 0.033044f
C1625 CF[9].n3 VSUBS 0.060534f
C1626 CF[9].n4 VSUBS 0.04139f
C1627 CF[9].n5 VSUBS 0.35865f
C1628 CF[9].t8 VSUBS 0.025568f
C1629 CF[9].t6 VSUBS 0.028145f
C1630 CF[9].n6 VSUBS 0.080875f
C1631 CF[9].n7 VSUBS 0.159286f
C1632 CF[9].t2 VSUBS 0.020356f
C1633 CF[9].t3 VSUBS 0.020356f
C1634 CF[9].t0 VSUBS 0.013232f
C1635 CF[9].t1 VSUBS 0.013232f
C1636 CF[9].n8 VSUBS 0.026463f
C1637 CF[9].n9 VSUBS 0.035727f
C1638 CF[9].n10 VSUBS 0.012817f
C1639 CF[9].n11 VSUBS 0.040713f
C1640 CF[9].n12 VSUBS 0.025438f
C1641 CF[9].n13 VSUBS 0.325177f
C1642 CF[9].n14 VSUBS 12.6286f
C1643 CF[3].t9 VSUBS 0.039629f
C1644 CF[3].t4 VSUBS 0.026514f
C1645 CF[3].n0 VSUBS 0.072417f
C1646 CF[3].n2 VSUBS 0.04757f
C1647 CF[3].t6 VSUBS 0.026514f
C1648 CF[3].t7 VSUBS 0.039629f
C1649 CF[3].n3 VSUBS 0.072598f
C1650 CF[3].n4 VSUBS 0.049639f
C1651 CF[3].n5 VSUBS 0.430132f
C1652 CF[3].t2 VSUBS 0.024413f
C1653 CF[3].t3 VSUBS 0.024413f
C1654 CF[3].t1 VSUBS 0.015869f
C1655 CF[3].t0 VSUBS 0.015869f
C1656 CF[3].n6 VSUBS 0.031738f
C1657 CF[3].n7 VSUBS 0.040773f
C1658 CF[3].n8 VSUBS 0.015372f
C1659 CF[3].n9 VSUBS 0.048827f
C1660 CF[3].n10 VSUBS 0.011529f
C1661 CF[3].n11 VSUBS 0.024476f
C1662 CF[3].t8 VSUBS 0.030512f
C1663 CF[3].t5 VSUBS 0.033609f
C1664 CF[3].n12 VSUBS 0.096252f
C1665 CF[3].n13 VSUBS 0.403523f
C1666 CF[3].n14 VSUBS 17.1092f
C1667 CF[8].t9 VSUBS 0.037662f
C1668 CF[8].t5 VSUBS 0.025198f
C1669 CF[8].n0 VSUBS 0.068823f
C1670 CF[8].n2 VSUBS 0.045209f
C1671 CF[8].t8 VSUBS 0.025198f
C1672 CF[8].t4 VSUBS 0.037662f
C1673 CF[8].n3 VSUBS 0.068995f
C1674 CF[8].n4 VSUBS 0.047175f
C1675 CF[8].n5 VSUBS 0.408285f
C1676 CF[8].t7 VSUBS 0.029142f
C1677 CF[8].t6 VSUBS 0.032079f
C1678 CF[8].n6 VSUBS 0.09218f
C1679 CF[8].n7 VSUBS 0.18155f
C1680 CF[8].t0 VSUBS 0.023202f
C1681 CF[8].t2 VSUBS 0.023202f
C1682 CF[8].t1 VSUBS 0.015081f
C1683 CF[8].t3 VSUBS 0.015081f
C1684 CF[8].n8 VSUBS 0.030162f
C1685 CF[8].n9 VSUBS 0.040721f
C1686 CF[8].n10 VSUBS 0.014609f
C1687 CF[8].n11 VSUBS 0.046404f
C1688 CF[8].n12 VSUBS 0.028776f
C1689 CF[8].n13 VSUBS 0.366382f
C1690 CF[8].n14 VSUBS 14.4899f
C1691 CF[4].t7 VSUBS 0.037633f
C1692 CF[4].t9 VSUBS 0.025178f
C1693 CF[4].n0 VSUBS 0.068769f
C1694 CF[4].n2 VSUBS 0.045173f
C1695 CF[4].t4 VSUBS 0.025178f
C1696 CF[4].t8 VSUBS 0.037633f
C1697 CF[4].n3 VSUBS 0.068941f
C1698 CF[4].n4 VSUBS 0.047138f
C1699 CF[4].n5 VSUBS 0.40946f
C1700 CF[4].t2 VSUBS 0.023184f
C1701 CF[4].t3 VSUBS 0.023184f
C1702 CF[4].t0 VSUBS 0.015069f
C1703 CF[4].t1 VSUBS 0.015069f
C1704 CF[4].n6 VSUBS 0.030139f
C1705 CF[4].n7 VSUBS 0.038719f
C1706 CF[4].n8 VSUBS 0.014597f
C1707 CF[4].n9 VSUBS 0.046367f
C1708 CF[4].n10 VSUBS 0.010948f
C1709 CF[4].n11 VSUBS 0.023493f
C1710 CF[4].t6 VSUBS 0.028975f
C1711 CF[4].t5 VSUBS 0.031916f
C1712 CF[4].n12 VSUBS 0.091404f
C1713 CF[4].n13 VSUBS 0.383391f
C1714 CF[4].n14 VSUBS 1.11424f
C1715 CF[4].n15 VSUBS 15.3714f
C1716 CF[5].t7 VSUBS 0.036489f
C1717 CF[5].t8 VSUBS 0.024413f
C1718 CF[5].n0 VSUBS 0.066678f
C1719 CF[5].n2 VSUBS 0.0438f
C1720 CF[5].t4 VSUBS 0.024413f
C1721 CF[5].t6 VSUBS 0.036489f
C1722 CF[5].n3 VSUBS 0.066845f
C1723 CF[5].n4 VSUBS 0.045705f
C1724 CF[5].n5 VSUBS 0.395563f
C1725 CF[5].t5 VSUBS 0.028094f
C1726 CF[5].t9 VSUBS 0.030946f
C1727 CF[5].n6 VSUBS 0.088625f
C1728 CF[5].t2 VSUBS 0.022479f
C1729 CF[5].t3 VSUBS 0.022479f
C1730 CF[5].t0 VSUBS 0.014611f
C1731 CF[5].t1 VSUBS 0.014611f
C1732 CF[5].n7 VSUBS 0.029223f
C1733 CF[5].n8 VSUBS 0.039452f
C1734 CF[5].n9 VSUBS 0.014153f
C1735 CF[5].n10 VSUBS 0.044958f
C1736 CF[5].n11 VSUBS 0.022197f
C1737 CF[5].n12 VSUBS 0.392725f
C1738 CF[5].n13 VSUBS 14.2556f
C1739 EN.t34 VSUBS 0.018406f
C1740 EN.t89 VSUBS 0.043122f
C1741 EN.n0 VSUBS 0.07648f
C1742 EN.n1 VSUBS 0.085792f
C1743 EN.n2 VSUBS 0.107342f
C1744 EN.t50 VSUBS 0.02364f
C1745 EN.t69 VSUBS 0.037535f
C1746 EN.n3 VSUBS 0.073218f
C1747 EN.n4 VSUBS 0.01581f
C1748 EN.n5 VSUBS 0.012134f
C1749 EN.n6 VSUBS 0.028806f
C1750 EN.n7 VSUBS 0.030818f
C1751 EN.n8 VSUBS 0.288981f
C1752 EN.t25 VSUBS 0.018406f
C1753 EN.t86 VSUBS 0.043122f
C1754 EN.n9 VSUBS 0.07648f
C1755 EN.n10 VSUBS 0.085792f
C1756 EN.n11 VSUBS 0.107342f
C1757 EN.t70 VSUBS 0.02364f
C1758 EN.t84 VSUBS 0.037535f
C1759 EN.n12 VSUBS 0.073218f
C1760 EN.n13 VSUBS 0.01581f
C1761 EN.n14 VSUBS 0.012134f
C1762 EN.n15 VSUBS 0.028806f
C1763 EN.n16 VSUBS 0.030818f
C1764 EN.n17 VSUBS 0.033883f
C1765 EN.n18 VSUBS 1.23519f
C1766 EN.t53 VSUBS 0.018406f
C1767 EN.t17 VSUBS 0.043122f
C1768 EN.n19 VSUBS 0.07648f
C1769 EN.n20 VSUBS 0.085792f
C1770 EN.n21 VSUBS 0.107342f
C1771 EN.t83 VSUBS 0.02364f
C1772 EN.t5 VSUBS 0.037535f
C1773 EN.n22 VSUBS 0.073218f
C1774 EN.n23 VSUBS 0.01581f
C1775 EN.n24 VSUBS 0.012134f
C1776 EN.n25 VSUBS 0.028806f
C1777 EN.n26 VSUBS 0.030818f
C1778 EN.n27 VSUBS 0.033883f
C1779 EN.n28 VSUBS 0.54049f
C1780 EN.t52 VSUBS 0.043122f
C1781 EN.t45 VSUBS 0.018406f
C1782 EN.n29 VSUBS 0.076571f
C1783 EN.n30 VSUBS 0.104561f
C1784 EN.n31 VSUBS 0.033029f
C1785 EN.t87 VSUBS 0.037535f
C1786 EN.t40 VSUBS 0.02364f
C1787 EN.n32 VSUBS 0.073218f
C1788 EN.n33 VSUBS 0.038803f
C1789 EN.n34 VSUBS 0.031253f
C1790 EN.n35 VSUBS 0.012879f
C1791 EN.n37 VSUBS 0.652055f
C1792 EN.t48 VSUBS 0.043122f
C1793 EN.t41 VSUBS 0.018406f
C1794 EN.n38 VSUBS 0.076571f
C1795 EN.n39 VSUBS 0.104561f
C1796 EN.n40 VSUBS 0.033029f
C1797 EN.t6 VSUBS 0.037535f
C1798 EN.t55 VSUBS 0.02364f
C1799 EN.n41 VSUBS 0.073218f
C1800 EN.n42 VSUBS 0.038803f
C1801 EN.n43 VSUBS 0.031253f
C1802 EN.n44 VSUBS 0.012879f
C1803 EN.n47 VSUBS 1.3874f
C1804 EN.t31 VSUBS 0.043122f
C1805 EN.t21 VSUBS 0.018406f
C1806 EN.n48 VSUBS 0.076571f
C1807 EN.n49 VSUBS 0.104561f
C1808 EN.n50 VSUBS 0.033029f
C1809 EN.t63 VSUBS 0.037535f
C1810 EN.t12 VSUBS 0.02364f
C1811 EN.n51 VSUBS 0.073218f
C1812 EN.n52 VSUBS 0.038803f
C1813 EN.n53 VSUBS 0.031253f
C1814 EN.n54 VSUBS 0.012879f
C1815 EN.n56 VSUBS 0.263108f
C1816 EN.t29 VSUBS 0.043122f
C1817 EN.t19 VSUBS 0.018406f
C1818 EN.n57 VSUBS 0.076571f
C1819 EN.n58 VSUBS 0.104561f
C1820 EN.n59 VSUBS 0.033029f
C1821 EN.t30 VSUBS 0.037535f
C1822 EN.t76 VSUBS 0.02364f
C1823 EN.n60 VSUBS 0.073218f
C1824 EN.n61 VSUBS 0.038803f
C1825 EN.n62 VSUBS 0.031253f
C1826 EN.n63 VSUBS 0.012879f
C1827 EN.n66 VSUBS 1.23519f
C1828 EN.t0 VSUBS 0.043122f
C1829 EN.t66 VSUBS 0.018406f
C1830 EN.n67 VSUBS 0.076571f
C1831 EN.n68 VSUBS 0.104561f
C1832 EN.n69 VSUBS 0.033029f
C1833 EN.t1 VSUBS 0.037535f
C1834 EN.t49 VSUBS 0.02364f
C1835 EN.n70 VSUBS 0.073218f
C1836 EN.n71 VSUBS 0.038803f
C1837 EN.n72 VSUBS 0.031253f
C1838 EN.n73 VSUBS 0.012879f
C1839 EN.n76 VSUBS 0.708607f
C1840 EN.n77 VSUBS 0.771176f
C1841 EN.n78 VSUBS 0.755362f
C1842 EN.t80 VSUBS 0.018406f
C1843 EN.t46 VSUBS 0.043122f
C1844 EN.n79 VSUBS 0.07648f
C1845 EN.n80 VSUBS 0.085792f
C1846 EN.n81 VSUBS 0.107342f
C1847 EN.t15 VSUBS 0.02364f
C1848 EN.t36 VSUBS 0.037535f
C1849 EN.n82 VSUBS 0.073218f
C1850 EN.n83 VSUBS 0.01581f
C1851 EN.n84 VSUBS 0.012134f
C1852 EN.n85 VSUBS 0.028806f
C1853 EN.n86 VSUBS 0.030818f
C1854 EN.n87 VSUBS 0.033883f
C1855 EN.n88 VSUBS 0.935018f
C1856 EN.t8 VSUBS 0.018406f
C1857 EN.t72 VSUBS 0.043122f
C1858 EN.n89 VSUBS 0.07648f
C1859 EN.n90 VSUBS 0.085792f
C1860 EN.n91 VSUBS 0.107342f
C1861 EN.t9 VSUBS 0.02364f
C1862 EN.t28 VSUBS 0.037535f
C1863 EN.n92 VSUBS 0.073218f
C1864 EN.n93 VSUBS 0.01581f
C1865 EN.n94 VSUBS 0.012134f
C1866 EN.n95 VSUBS 0.028806f
C1867 EN.n96 VSUBS 0.030818f
C1868 EN.n97 VSUBS 0.033883f
C1869 EN.n98 VSUBS 0.961349f
C1870 EN.n99 VSUBS 0.023332f
C1871 EN.t7 VSUBS 0.037535f
C1872 EN.t85 VSUBS 0.02364f
C1873 EN.n100 VSUBS 0.073218f
C1874 EN.n101 VSUBS 0.01581f
C1875 EN.n102 VSUBS 0.012361f
C1876 EN.t35 VSUBS 0.043122f
C1877 EN.t68 VSUBS 0.018406f
C1878 EN.n103 VSUBS 0.07648f
C1879 EN.n104 VSUBS 0.085792f
C1880 EN.n105 VSUBS 0.107342f
C1881 EN.n106 VSUBS 0.054606f
C1882 EN.n107 VSUBS 0.023332f
C1883 EN.t44 VSUBS 0.037535f
C1884 EN.t24 VSUBS 0.02364f
C1885 EN.n108 VSUBS 0.073218f
C1886 EN.n109 VSUBS 0.01581f
C1887 EN.n110 VSUBS 0.012361f
C1888 EN.t10 VSUBS 0.043122f
C1889 EN.t37 VSUBS 0.018406f
C1890 EN.n111 VSUBS 0.07648f
C1891 EN.n112 VSUBS 0.085792f
C1892 EN.n113 VSUBS 0.107342f
C1893 EN.n114 VSUBS 0.320495f
C1894 EN.n115 VSUBS 0.023332f
C1895 EN.t47 VSUBS 0.037535f
C1896 EN.t27 VSUBS 0.02364f
C1897 EN.n116 VSUBS 0.073218f
C1898 EN.n117 VSUBS 0.01581f
C1899 EN.n118 VSUBS 0.012361f
C1900 EN.t4 VSUBS 0.043122f
C1901 EN.t42 VSUBS 0.018406f
C1902 EN.n119 VSUBS 0.07648f
C1903 EN.n120 VSUBS 0.085792f
C1904 EN.n121 VSUBS 0.107342f
C1905 EN.n122 VSUBS 0.054606f
C1906 EN.n123 VSUBS 1.26967f
C1907 EN.n124 VSUBS 0.023332f
C1908 EN.t39 VSUBS 0.037535f
C1909 EN.t18 VSUBS 0.02364f
C1910 EN.n125 VSUBS 0.073218f
C1911 EN.n126 VSUBS 0.01581f
C1912 EN.n127 VSUBS 0.012361f
C1913 EN.t38 VSUBS 0.043122f
C1914 EN.t71 VSUBS 0.018406f
C1915 EN.n128 VSUBS 0.07648f
C1916 EN.n129 VSUBS 0.085792f
C1917 EN.n130 VSUBS 0.107342f
C1918 EN.n131 VSUBS 0.054606f
C1919 EN.n132 VSUBS 1.00988f
C1920 EN.n133 VSUBS 0.023332f
C1921 EN.t2 VSUBS 0.037535f
C1922 EN.t82 VSUBS 0.02364f
C1923 EN.n134 VSUBS 0.073218f
C1924 EN.n135 VSUBS 0.01581f
C1925 EN.n136 VSUBS 0.012361f
C1926 EN.t75 VSUBS 0.043122f
C1927 EN.t13 VSUBS 0.018406f
C1928 EN.n137 VSUBS 0.07648f
C1929 EN.n138 VSUBS 0.085792f
C1930 EN.n139 VSUBS 0.107342f
C1931 EN.n140 VSUBS 0.054606f
C1932 EN.n141 VSUBS 1.00988f
C1933 EN.n142 VSUBS 0.023332f
C1934 EN.t43 VSUBS 0.037535f
C1935 EN.t22 VSUBS 0.02364f
C1936 EN.n143 VSUBS 0.073218f
C1937 EN.n144 VSUBS 0.01581f
C1938 EN.n145 VSUBS 0.012361f
C1939 EN.t65 VSUBS 0.043122f
C1940 EN.t77 VSUBS 0.018406f
C1941 EN.n146 VSUBS 0.07648f
C1942 EN.n147 VSUBS 0.085792f
C1943 EN.n148 VSUBS 0.107342f
C1944 EN.n149 VSUBS 0.054606f
C1945 EN.n150 VSUBS 1.00766f
C1946 EN.n151 VSUBS 0.914236f
C1947 EN.n152 VSUBS 0.023332f
C1948 EN.t51 VSUBS 0.043122f
C1949 EN.t57 VSUBS 0.018406f
C1950 EN.n153 VSUBS 0.07648f
C1951 EN.n154 VSUBS 0.085792f
C1952 EN.n155 VSUBS 0.107342f
C1953 EN.t26 VSUBS 0.037535f
C1954 EN.t79 VSUBS 0.02364f
C1955 EN.n156 VSUBS 0.073218f
C1956 EN.n157 VSUBS 0.01581f
C1957 EN.n158 VSUBS 0.012134f
C1958 EN.n159 VSUBS 0.028795f
C1959 EN.n160 VSUBS 0.031128f
C1960 EN.n161 VSUBS 0.027646f
C1961 EN.n162 VSUBS 0.914236f
C1962 EN.n163 VSUBS 0.023332f
C1963 EN.t58 VSUBS 0.043122f
C1964 EN.t67 VSUBS 0.018406f
C1965 EN.n164 VSUBS 0.07648f
C1966 EN.n165 VSUBS 0.085792f
C1967 EN.n166 VSUBS 0.107342f
C1968 EN.t59 VSUBS 0.037535f
C1969 EN.t14 VSUBS 0.02364f
C1970 EN.n167 VSUBS 0.073218f
C1971 EN.n168 VSUBS 0.01581f
C1972 EN.n169 VSUBS 0.012134f
C1973 EN.n170 VSUBS 0.028795f
C1974 EN.n171 VSUBS 0.031128f
C1975 EN.n172 VSUBS 0.027646f
C1976 EN.n173 VSUBS 1.00766f
C1977 EN.n174 VSUBS 0.023332f
C1978 EN.t88 VSUBS 0.043122f
C1979 EN.t3 VSUBS 0.018406f
C1980 EN.n175 VSUBS 0.07648f
C1981 EN.n176 VSUBS 0.085792f
C1982 EN.n177 VSUBS 0.107342f
C1983 EN.t20 VSUBS 0.037535f
C1984 EN.t73 VSUBS 0.02364f
C1985 EN.n178 VSUBS 0.073218f
C1986 EN.n179 VSUBS 0.01581f
C1987 EN.n180 VSUBS 0.012134f
C1988 EN.n181 VSUBS 0.028795f
C1989 EN.n182 VSUBS 0.031128f
C1990 EN.n183 VSUBS 0.027646f
C1991 EN.n184 VSUBS 1.00988f
C1992 EN.n185 VSUBS 0.023332f
C1993 EN.t56 VSUBS 0.043122f
C1994 EN.t60 VSUBS 0.018406f
C1995 EN.n186 VSUBS 0.07648f
C1996 EN.n187 VSUBS 0.085792f
C1997 EN.n188 VSUBS 0.107342f
C1998 EN.t32 VSUBS 0.037535f
C1999 EN.t81 VSUBS 0.02364f
C2000 EN.n189 VSUBS 0.073218f
C2001 EN.n190 VSUBS 0.01581f
C2002 EN.n191 VSUBS 0.012134f
C2003 EN.n192 VSUBS 0.028795f
C2004 EN.n193 VSUBS 0.031128f
C2005 EN.n194 VSUBS 0.027646f
C2006 EN.n195 VSUBS 1.00988f
C2007 EN.n196 VSUBS 0.023332f
C2008 EN.t23 VSUBS 0.043122f
C2009 EN.t33 VSUBS 0.018406f
C2010 EN.n197 VSUBS 0.07648f
C2011 EN.n198 VSUBS 0.085792f
C2012 EN.n199 VSUBS 0.107342f
C2013 EN.t62 VSUBS 0.037535f
C2014 EN.t16 VSUBS 0.02364f
C2015 EN.n200 VSUBS 0.073218f
C2016 EN.n201 VSUBS 0.01581f
C2017 EN.n202 VSUBS 0.012134f
C2018 EN.n203 VSUBS 0.028795f
C2019 EN.n204 VSUBS 0.031128f
C2020 EN.n205 VSUBS 0.027646f
C2021 EN.n206 VSUBS 1.00988f
C2022 EN.n207 VSUBS 0.023332f
C2023 EN.t78 VSUBS 0.043122f
C2024 EN.t74 VSUBS 0.018406f
C2025 EN.n208 VSUBS 0.07648f
C2026 EN.n209 VSUBS 0.085792f
C2027 EN.n210 VSUBS 0.107342f
C2028 EN.t11 VSUBS 0.037535f
C2029 EN.t61 VSUBS 0.02364f
C2030 EN.n211 VSUBS 0.073218f
C2031 EN.n212 VSUBS 0.01581f
C2032 EN.n213 VSUBS 0.012134f
C2033 EN.n214 VSUBS 0.028795f
C2034 EN.n215 VSUBS 0.031128f
C2035 EN.n216 VSUBS 0.027646f
C2036 EN.n217 VSUBS 1.01423f
C2037 EN.n218 VSUBS 3.90286f
C2038 EN.n219 VSUBS 5.98024f
C2039 EN.t64 VSUBS 0.0337f
C2040 EN.t54 VSUBS 0.037097f
C2041 EN.n220 VSUBS 0.106598f
C2042 EN.n221 VSUBS 0.215797f
C2043 EN.n222 VSUBS 21.9615f
C2044 DOUT[0].t2 VSUBS 0.020845f
C2045 DOUT[0].t3 VSUBS 0.020845f
C2046 DOUT[0].t1 VSUBS 0.013549f
C2047 DOUT[0].t0 VSUBS 0.013549f
C2048 DOUT[0].n0 VSUBS 0.027098f
C2049 DOUT[0].n1 VSUBS 0.036584f
C2050 DOUT[0].n2 VSUBS 0.013124f
C2051 DOUT[0].n3 VSUBS 0.041689f
C2052 DOUT[0].n4 VSUBS 0.043854f
C2053 DOUT[0].n5 VSUBS 9.764151f
C2054 CLK.t10 VSUBS 0.042487f
C2055 CLK.t17 VSUBS 0.028426f
C2056 CLK.n0 VSUBS 0.07764f
C2057 CLK.n1 VSUBS 0.023072f
C2058 CLK.t27 VSUBS 0.042487f
C2059 CLK.t35 VSUBS 0.028426f
C2060 CLK.n2 VSUBS 0.07764f
C2061 CLK.n3 VSUBS 0.023072f
C2062 CLK.n4 VSUBS 1.3595f
C2063 CLK.t3 VSUBS 0.042487f
C2064 CLK.t6 VSUBS 0.028426f
C2065 CLK.n5 VSUBS 0.07764f
C2066 CLK.n6 VSUBS 0.023072f
C2067 CLK.n7 VSUBS 0.974052f
C2068 CLK.t25 VSUBS 0.042487f
C2069 CLK.t4 VSUBS 0.028426f
C2070 CLK.n8 VSUBS 0.07764f
C2071 CLK.n9 VSUBS 0.023072f
C2072 CLK.n10 VSUBS 0.497086f
C2073 CLK.t7 VSUBS 0.028426f
C2074 CLK.t12 VSUBS 0.042487f
C2075 CLK.n11 VSUBS 0.078526f
C2076 CLK.n12 VSUBS 0.034907f
C2077 CLK.n13 VSUBS 0.547362f
C2078 CLK.t5 VSUBS 0.028426f
C2079 CLK.t8 VSUBS 0.042487f
C2080 CLK.n14 VSUBS 0.078526f
C2081 CLK.n15 VSUBS 0.034907f
C2082 CLK.n16 VSUBS 0.972006f
C2083 CLK.t14 VSUBS 0.028426f
C2084 CLK.t19 VSUBS 0.042487f
C2085 CLK.n17 VSUBS 0.078526f
C2086 CLK.n18 VSUBS 0.034907f
C2087 CLK.n19 VSUBS 0.972006f
C2088 CLK.t40 VSUBS 0.028426f
C2089 CLK.t2 VSUBS 0.042487f
C2090 CLK.n20 VSUBS 0.078526f
C2091 CLK.n21 VSUBS 0.034907f
C2092 CLK.n22 VSUBS 0.959365f
C2093 CLK.t34 VSUBS 0.028426f
C2094 CLK.t0 VSUBS 0.042487f
C2095 CLK.n23 VSUBS 0.078526f
C2096 CLK.n24 VSUBS 0.035292f
C2097 CLK.n25 VSUBS 0.729637f
C2098 CLK.n26 VSUBS 0.663742f
C2099 CLK.t13 VSUBS 0.042487f
C2100 CLK.t18 VSUBS 0.028426f
C2101 CLK.n27 VSUBS 0.07764f
C2102 CLK.n28 VSUBS 0.023072f
C2103 CLK.n29 VSUBS 0.538245f
C2104 CLK.t32 VSUBS 0.042487f
C2105 CLK.t29 VSUBS 0.028426f
C2106 CLK.n30 VSUBS 0.07764f
C2107 CLK.n31 VSUBS 0.023072f
C2108 CLK.t16 VSUBS 0.042487f
C2109 CLK.t15 VSUBS 0.028426f
C2110 CLK.n32 VSUBS 0.07764f
C2111 CLK.n33 VSUBS 0.023072f
C2112 CLK.n34 VSUBS 1.44588f
C2113 CLK.t23 VSUBS 0.042487f
C2114 CLK.t21 VSUBS 0.028426f
C2115 CLK.n35 VSUBS 0.07764f
C2116 CLK.n36 VSUBS 0.023072f
C2117 CLK.n37 VSUBS 1.01744f
C2118 CLK.t37 VSUBS 0.042487f
C2119 CLK.t36 VSUBS 0.028426f
C2120 CLK.n38 VSUBS 0.07764f
C2121 CLK.n39 VSUBS 0.023072f
C2122 CLK.n40 VSUBS 1.01744f
C2123 CLK.t33 VSUBS 0.042487f
C2124 CLK.t30 VSUBS 0.028426f
C2125 CLK.n41 VSUBS 0.07764f
C2126 CLK.n42 VSUBS 0.023072f
C2127 CLK.n43 VSUBS 1.01528f
C2128 CLK.t38 VSUBS 0.042487f
C2129 CLK.t42 VSUBS 0.028426f
C2130 CLK.n44 VSUBS 0.07764f
C2131 CLK.n45 VSUBS 0.023072f
C2132 CLK.t20 VSUBS 0.042487f
C2133 CLK.t22 VSUBS 0.028426f
C2134 CLK.n46 VSUBS 0.07764f
C2135 CLK.n47 VSUBS 0.023072f
C2136 CLK.n48 VSUBS 1.44592f
C2137 CLK.t24 VSUBS 0.042487f
C2138 CLK.t26 VSUBS 0.028426f
C2139 CLK.n49 VSUBS 0.07764f
C2140 CLK.n50 VSUBS 0.023072f
C2141 CLK.n51 VSUBS 1.01817f
C2142 CLK.t41 VSUBS 0.042487f
C2143 CLK.t1 VSUBS 0.028426f
C2144 CLK.n52 VSUBS 0.07764f
C2145 CLK.n53 VSUBS 0.023072f
C2146 CLK.n54 VSUBS 1.01678f
C2147 CLK.t39 VSUBS 0.042487f
C2148 CLK.t43 VSUBS 0.028426f
C2149 CLK.n55 VSUBS 0.07764f
C2150 CLK.n56 VSUBS 0.023072f
C2151 CLK.n57 VSUBS 1.01462f
C2152 CLK.t28 VSUBS 0.042487f
C2153 CLK.t31 VSUBS 0.028426f
C2154 CLK.n58 VSUBS 0.07764f
C2155 CLK.n59 VSUBS 0.023072f
C2156 CLK.n60 VSUBS 0.894705f
C2157 CLK.t11 VSUBS 0.042487f
C2158 CLK.t9 VSUBS 0.028426f
C2159 CLK.n61 VSUBS 0.07764f
C2160 CLK.n62 VSUBS 0.023072f
C2161 CLK.n63 VSUBS 1.00243f
C2162 CLK.n64 VSUBS 3.34046f
C2163 CLK.n65 VSUBS 21.8766f
C2164 out_latch_0.FINAL.t8 VSUBS 0.020864f
C2165 out_latch_0.FINAL.t10 VSUBS 0.020864f
C2166 out_latch_0.FINAL.n0 VSUBS 0.044497f
C2167 out_latch_0.FINAL.t4 VSUBS 0.013562f
C2168 out_latch_0.FINAL.t0 VSUBS 0.013562f
C2169 out_latch_0.FINAL.n1 VSUBS 0.028495f
C2170 out_latch_0.FINAL.t6 VSUBS 0.013562f
C2171 out_latch_0.FINAL.t2 VSUBS 0.013562f
C2172 out_latch_0.FINAL.n2 VSUBS 0.028495f
C2173 out_latch_0.FINAL.t7 VSUBS 0.013562f
C2174 out_latch_0.FINAL.t5 VSUBS 0.013562f
C2175 out_latch_0.FINAL.n3 VSUBS 0.040686f
C2176 out_latch_0.FINAL.n4 VSUBS 0.106188f
C2177 out_latch_0.FINAL.n5 VSUBS 0.063525f
C2178 out_latch_0.FINAL.t1 VSUBS 0.013562f
C2179 out_latch_0.FINAL.t3 VSUBS 0.013562f
C2180 out_latch_0.FINAL.n6 VSUBS 0.029068f
C2181 out_latch_0.FINAL.n7 VSUBS 0.052102f
C2182 out_latch_0.FINAL.t18 VSUBS 0.015724f
C2183 out_latch_0.FINAL.t19 VSUBS 0.022881f
C2184 out_latch_0.FINAL.n8 VSUBS 0.06649f
C2185 out_latch_0.FINAL.n9 VSUBS 0.023229f
C2186 out_latch_0.FINAL.t17 VSUBS 0.022881f
C2187 out_latch_0.FINAL.t16 VSUBS 0.015724f
C2188 out_latch_0.FINAL.n10 VSUBS 0.06649f
C2189 out_latch_0.FINAL.n11 VSUBS 0.015841f
C2190 out_latch_0.FINAL.n12 VSUBS 0.037347f
C2191 out_latch_0.FINAL.n13 VSUBS 0.401317f
C2192 out_latch_0.FINAL.n14 VSUBS 16.4227f
C2193 out_latch_0.FINAL.n15 VSUBS 0.025223f
C2194 out_latch_0.FINAL.t13 VSUBS 0.020864f
C2195 out_latch_0.FINAL.t9 VSUBS 0.020864f
C2196 out_latch_0.FINAL.n16 VSUBS 0.044497f
C2197 out_latch_0.FINAL.t14 VSUBS 0.020864f
C2198 out_latch_0.FINAL.t12 VSUBS 0.020864f
C2199 out_latch_0.FINAL.n17 VSUBS 0.05604f
C2200 out_latch_0.FINAL.n18 VSUBS 0.142927f
C2201 out_latch_0.FINAL.t11 VSUBS 0.020864f
C2202 out_latch_0.FINAL.t15 VSUBS 0.020864f
C2203 out_latch_0.FINAL.n19 VSUBS 0.044497f
C2204 out_latch_0.FINAL.n20 VSUBS 0.08157f
C2205 out_latch_0.FINAL.n21 VSUBS 0.02962f
C2206 cdac_ctrl_0.x2.X.t2 VSUBS 0.035376f
C2207 cdac_ctrl_0.x2.X.t8 VSUBS 0.035376f
C2208 cdac_ctrl_0.x2.X.n0 VSUBS 0.070779f
C2209 cdac_ctrl_0.x2.X.t21 VSUBS 0.044432f
C2210 cdac_ctrl_0.x2.X.t16 VSUBS 0.048911f
C2211 cdac_ctrl_0.x2.X.n1 VSUBS 0.140546f
C2212 cdac_ctrl_0.x2.X.t30 VSUBS 0.044432f
C2213 cdac_ctrl_0.x2.X.t25 VSUBS 0.048911f
C2214 cdac_ctrl_0.x2.X.n2 VSUBS 0.140546f
C2215 cdac_ctrl_0.x2.X.n3 VSUBS 1.34878f
C2216 cdac_ctrl_0.x2.X.t27 VSUBS 0.044432f
C2217 cdac_ctrl_0.x2.X.t33 VSUBS 0.048911f
C2218 cdac_ctrl_0.x2.X.n4 VSUBS 0.140546f
C2219 cdac_ctrl_0.x2.X.n5 VSUBS 0.930404f
C2220 cdac_ctrl_0.x2.X.t34 VSUBS 0.044432f
C2221 cdac_ctrl_0.x2.X.t32 VSUBS 0.048911f
C2222 cdac_ctrl_0.x2.X.n6 VSUBS 0.140546f
C2223 cdac_ctrl_0.x2.X.n7 VSUBS 0.930404f
C2224 cdac_ctrl_0.x2.X.t28 VSUBS 0.044432f
C2225 cdac_ctrl_0.x2.X.t18 VSUBS 0.048911f
C2226 cdac_ctrl_0.x2.X.n8 VSUBS 0.140546f
C2227 cdac_ctrl_0.x2.X.n9 VSUBS 0.930404f
C2228 cdac_ctrl_0.x2.X.t26 VSUBS 0.044432f
C2229 cdac_ctrl_0.x2.X.t29 VSUBS 0.048911f
C2230 cdac_ctrl_0.x2.X.n10 VSUBS 0.140546f
C2231 cdac_ctrl_0.x2.X.n11 VSUBS 0.930404f
C2232 cdac_ctrl_0.x2.X.t22 VSUBS 0.044432f
C2233 cdac_ctrl_0.x2.X.t24 VSUBS 0.048911f
C2234 cdac_ctrl_0.x2.X.n12 VSUBS 0.140546f
C2235 cdac_ctrl_0.x2.X.n13 VSUBS 0.930404f
C2236 cdac_ctrl_0.x2.X.t19 VSUBS 0.044432f
C2237 cdac_ctrl_0.x2.X.t20 VSUBS 0.048911f
C2238 cdac_ctrl_0.x2.X.n14 VSUBS 0.140546f
C2239 cdac_ctrl_0.x2.X.n15 VSUBS 0.930404f
C2240 cdac_ctrl_0.x2.X.t23 VSUBS 0.044432f
C2241 cdac_ctrl_0.x2.X.t35 VSUBS 0.048911f
C2242 cdac_ctrl_0.x2.X.n16 VSUBS 0.140546f
C2243 cdac_ctrl_0.x2.X.n17 VSUBS 0.930404f
C2244 cdac_ctrl_0.x2.X.t17 VSUBS 0.044432f
C2245 cdac_ctrl_0.x2.X.t31 VSUBS 0.048911f
C2246 cdac_ctrl_0.x2.X.n18 VSUBS 0.140546f
C2247 cdac_ctrl_0.x2.X.n19 VSUBS 0.774865f
C2248 cdac_ctrl_0.x2.X.n20 VSUBS 0.036632f
C2249 cdac_ctrl_0.x2.X.t13 VSUBS 0.022994f
C2250 cdac_ctrl_0.x2.X.t12 VSUBS 0.022994f
C2251 cdac_ctrl_0.x2.X.n21 VSUBS 0.048313f
C2252 cdac_ctrl_0.x2.X.t0 VSUBS 0.022994f
C2253 cdac_ctrl_0.x2.X.t14 VSUBS 0.022994f
C2254 cdac_ctrl_0.x2.X.n22 VSUBS 0.048313f
C2255 cdac_ctrl_0.x2.X.t6 VSUBS 0.022994f
C2256 cdac_ctrl_0.x2.X.t4 VSUBS 0.022994f
C2257 cdac_ctrl_0.x2.X.n23 VSUBS 0.068982f
C2258 cdac_ctrl_0.x2.X.n24 VSUBS 0.180043f
C2259 cdac_ctrl_0.x2.X.n25 VSUBS 0.107706f
C2260 cdac_ctrl_0.x2.X.t11 VSUBS 0.022994f
C2261 cdac_ctrl_0.x2.X.t9 VSUBS 0.022994f
C2262 cdac_ctrl_0.x2.X.n26 VSUBS 0.049285f
C2263 cdac_ctrl_0.x2.X.n27 VSUBS 0.088339f
C2264 cdac_ctrl_0.x2.X.t10 VSUBS 0.035376f
C2265 cdac_ctrl_0.x2.X.t3 VSUBS 0.035376f
C2266 cdac_ctrl_0.x2.X.n28 VSUBS 0.075445f
C2267 cdac_ctrl_0.x2.X.t7 VSUBS 0.035376f
C2268 cdac_ctrl_0.x2.X.t15 VSUBS 0.035376f
C2269 cdac_ctrl_0.x2.X.n29 VSUBS 0.075445f
C2270 cdac_ctrl_0.x2.X.t1 VSUBS 0.035376f
C2271 cdac_ctrl_0.x2.X.t5 VSUBS 0.035376f
C2272 cdac_ctrl_0.x2.X.n30 VSUBS 0.095016f
C2273 cdac_ctrl_0.x2.X.n31 VSUBS 0.242333f
C2274 cdac_ctrl_0.x2.X.n32 VSUBS 0.138303f
C2275 cdac_ctrl_0.x2.X.n33 VSUBS 0.052552f
C2276 VSSD.t260 VSUBS 0.13659f
C2277 VSSD.t418 VSUBS 0.155048f
C2278 VSSD.t258 VSUBS 0.155048f
C2279 VSSD.t170 VSUBS 0.155048f
C2280 VSSD.t172 VSUBS 0.155048f
C2281 VSSD.t191 VSUBS 0.155048f
C2282 VSSD.t193 VSUBS 0.155048f
C2283 VSSD.t246 VSUBS 0.155048f
C2284 VSSD.t248 VSUBS 0.155048f
C2285 VSSD.t349 VSUBS 0.155048f
C2286 VSSD.t351 VSUBS 0.261183f
C2287 VSSD.t370 VSUBS 0.137513f
C2288 VSSD.t631 VSUBS 0.312866f
C2289 VSSD.t365 VSUBS 0.323018f
C2290 VSSD.t116 VSUBS 0.176275f
C2291 VSSD.t135 VSUBS 0.241802f
C2292 VSSD.t320 VSUBS 0.219652f
C2293 VSSD.t1071 VSUBS 0.188273f
C2294 VSSD.t85 VSUBS 0.213192f
C2295 VSSD.t787 VSUBS 0.191965f
C2296 VSSD.t630 VSUBS 0.189196f
C2297 VSSD.t7 VSUBS 0.226112f
C2298 VSSD.t1026 VSUBS 0.221498f
C2299 VSSD.t531 VSUBS 0.275949f
C2300 VSSD.t32 VSUBS 0.269489f
C2301 VSSD.t26 VSUBS 0.198425f
C2302 VSSD.t81 VSUBS 0.137513f
C2303 VSSD.t521 VSUBS 0.312866f
C2304 VSSD.t625 VSUBS 0.323018f
C2305 VSSD.t4 VSUBS 0.176275f
C2306 VSSD.t890 VSUBS 0.241802f
C2307 VSSD.t151 VSUBS 0.219652f
C2308 VSSD.t1041 VSUBS 0.188273f
C2309 VSSD.t404 VSUBS 0.213192f
C2310 VSSD.t889 VSUBS 0.191965f
C2311 VSSD.t520 VSUBS 0.189196f
C2312 VSSD.t286 VSUBS 0.226112f
C2313 VSSD.t1078 VSUBS 0.221498f
C2314 VSSD.t756 VSUBS 0.275949f
C2315 VSSD.t288 VSUBS 0.269489f
C2316 VSSD.t684 VSUBS 0.198425f
C2317 VSSD.t673 VSUBS 0.137513f
C2318 VSSD.t424 VSUBS 0.312866f
C2319 VSSD.t536 VSUBS 0.323018f
C2320 VSSD.t711 VSUBS 0.176275f
C2321 VSSD.t614 VSUBS 0.241802f
C2322 VSSD.t464 VSUBS 0.219652f
C2323 VSSD.t1047 VSUBS 0.188273f
C2324 VSSD.t834 VSUBS 0.213192f
C2325 VSSD.t615 VSUBS 0.191965f
C2326 VSSD.t426 VSUBS 0.189196f
C2327 VSSD.t77 VSUBS 0.226112f
C2328 VSSD.t1024 VSUBS 0.221498f
C2329 VSSD.t560 VSUBS 0.275949f
C2330 VSSD.t502 VSUBS 0.269489f
C2331 VSSD.t75 VSUBS 0.198425f
C2332 VSSD.t654 VSUBS 0.137513f
C2333 VSSD.t59 VSUBS 0.312866f
C2334 VSSD.t30 VSUBS 0.323018f
C2335 VSSD.t58 VSUBS 0.176275f
C2336 VSSD.t335 VSUBS 0.241802f
C2337 VSSD.t142 VSUBS 0.219652f
C2338 VSSD.t1053 VSUBS 0.188273f
C2339 VSSD.t34 VSUBS 0.213192f
C2340 VSSD.t157 VSUBS 0.191965f
C2341 VSSD.t61 VSUBS 0.189196f
C2342 VSSD.t127 VSUBS 0.226112f
C2343 VSSD.t1035 VSUBS 0.221498f
C2344 VSSD.t380 VSUBS 0.275949f
C2345 VSSD.t87 VSUBS 0.269489f
C2346 VSSD.t89 VSUBS 0.198425f
C2347 VSSD.t2 VSUBS 0.137513f
C2348 VSSD.t870 VSUBS 0.312866f
C2349 VSSD.t363 VSUBS 0.323018f
C2350 VSSD.t284 VSUBS 0.176275f
C2351 VSSD.t590 VSUBS 0.241802f
C2352 VSSD.t272 VSUBS 0.219652f
C2353 VSSD.t1020 VSUBS 0.188273f
C2354 VSSD.t388 VSUBS 0.213192f
C2355 VSSD.t775 VSUBS 0.191965f
C2356 VSSD.t285 VSUBS 0.189196f
C2357 VSSD.t137 VSUBS 0.226112f
C2358 VSSD.t1006 VSUBS 0.221498f
C2359 VSSD.t273 VSUBS 0.275949f
C2360 VSSD.t139 VSUBS 0.269489f
C2361 VSSD.t168 VSUBS 0.198425f
C2362 VSSD.t447 VSUBS 0.137513f
C2363 VSSD.t28 VSUBS 0.312866f
C2364 VSSD.t899 VSUBS 0.323018f
C2365 VSSD.t112 VSUBS 0.176275f
C2366 VSSD.t591 VSUBS 0.241802f
C2367 VSSD.t133 VSUBS 0.219652f
C2368 VSSD.t1030 VSUBS 0.188273f
C2369 VSSD.t493 VSUBS 0.213192f
C2370 VSSD.t95 VSUBS 0.191965f
C2371 VSSD.t601 VSUBS 0.189196f
C2372 VSSD.t801 VSUBS 0.226112f
C2373 VSSD.t1061 VSUBS 0.221498f
C2374 VSSD.t68 VSUBS 0.275949f
C2375 VSSD.t585 VSUBS 0.269489f
C2376 VSSD.t959 VSUBS 0.198425f
C2377 VSSD.t123 VSUBS 0.137513f
C2378 VSSD.t790 VSUBS 0.312866f
C2379 VSSD.t97 VSUBS 0.323018f
C2380 VSSD.t190 VSUBS 0.176275f
C2381 VSSD.t444 VSUBS 0.241802f
C2382 VSSD.t538 VSUBS 0.219652f
C2383 VSSD.t1022 VSUBS 0.188273f
C2384 VSSD.t178 VSUBS 0.213192f
C2385 VSSD.t589 VSUBS 0.191965f
C2386 VSSD.t839 VSUBS 0.189196f
C2387 VSSD.t578 VSUBS 0.226112f
C2388 VSSD.t1058 VSUBS 0.221498f
C2389 VSSD.t465 VSUBS 0.275949f
C2390 VSSD.t41 VSUBS 0.269489f
C2391 VSSD.t79 VSUBS 0.198425f
C2392 VSSD.t229 VSUBS 0.137513f
C2393 VSSD.t436 VSUBS 0.312866f
C2394 VSSD.t570 VSUBS 0.323018f
C2395 VSSD.t150 VSUBS 0.176275f
C2396 VSSD.t935 VSUBS 0.241802f
C2397 VSSD.t926 VSUBS 0.219652f
C2398 VSSD.t1008 VSUBS 0.188273f
C2399 VSSD.t678 VSUBS 0.213192f
C2400 VSSD.t534 VSUBS 0.191965f
C2401 VSSD.t149 VSUBS 0.189196f
C2402 VSSD.t566 VSUBS 0.226112f
C2403 VSSD.t1039 VSUBS 0.221498f
C2404 VSSD.t243 VSUBS 0.275949f
C2405 VSSD.t564 VSUBS 0.269489f
C2406 VSSD.t602 VSUBS 0.198425f
C2407 VSSD.t523 VSUBS 0.137513f
C2408 VSSD.t202 VSUBS 0.312866f
C2409 VSSD.t227 VSUBS 0.323018f
C2410 VSSD.t201 VSUBS 0.176275f
C2411 VSSD.t443 VSUBS 0.241802f
C2412 VSSD.t505 VSUBS 0.219652f
C2413 VSSD.t1045 VSUBS 0.188273f
C2414 VSSD.t840 VSUBS 0.213192f
C2415 VSSD.t744 VSUBS 0.191965f
C2416 VSSD.t200 VSUBS 0.189196f
C2417 VSSD.t303 VSUBS 0.226112f
C2418 VSSD.t1012 VSUBS 0.221498f
C2419 VSSD.t584 VSUBS 0.275949f
C2420 VSSD.t733 VSUBS 0.269489f
C2421 VSSD.t917 VSUBS 0.198425f
C2422 VSSD.t256 VSUBS 0.137513f
C2423 VSSD.t24 VSUBS 0.312866f
C2424 VSSD.t897 VSUBS 0.323018f
C2425 VSSD.t23 VSUBS 0.176275f
C2426 VSSD.t69 VSUBS 0.241802f
C2427 VSSD.t452 VSUBS 0.219652f
C2428 VSSD.t1037 VSUBS 0.188273f
C2429 VSSD.t344 VSUBS 0.213192f
C2430 VSSD.t70 VSUBS 0.191965f
C2431 VSSD.t22 VSUBS 0.189196f
C2432 VSSD.t498 VSUBS 0.226112f
C2433 VSSD.t1018 VSUBS 0.221498f
C2434 VSSD.t519 VSUBS 0.275949f
C2435 VSSD.t798 VSUBS 0.269489f
C2436 VSSD.t106 VSUBS 0.206731f
C2437 VSSD.n1 VSUBS 0.249247p
C2438 VSSD.n2 VSUBS 0.221083p
C2439 VSSD.t639 VSUBS 8.68217f
C2440 VSSD.n3 VSUBS 0.156946p
C2441 VSSD.t293 VSUBS 0.024414f
C2442 VSSD.n4 VSUBS 0.028345f
C2443 VSSD.t291 VSUBS 0.028005f
C2444 VSSD.n6 VSUBS 0.03123f
C2445 VSSD.n7 VSUBS 0.03123f
C2446 VSSD.t183 VSUBS 0.024724f
C2447 VSSD.n9 VSUBS 0.03123f
C2448 VSSD.t1087 VSUBS 0.010396f
C2449 VSSD.n10 VSUBS 0.018748f
C2450 VSSD.n11 VSUBS 0.018565f
C2451 VSSD.n13 VSUBS 0.03123f
C2452 VSSD.t92 VSUBS 0.013879f
C2453 VSSD.n14 VSUBS 0.017846f
C2454 VSSD.n15 VSUBS 0.029746f
C2455 VSSD.t401 VSUBS 0.013879f
C2456 VSSD.n16 VSUBS 0.017846f
C2457 VSSD.n17 VSUBS 0.011061f
C2458 VSSD.n18 VSUBS 0.03123f
C2459 VSSD.t1089 VSUBS 0.010396f
C2460 VSSD.n19 VSUBS 0.018748f
C2461 VSSD.t575 VSUBS 0.024724f
C2462 VSSD.n20 VSUBS 0.036733f
C2463 VSSD.n21 VSUBS 0.03123f
C2464 VSSD.t383 VSUBS 0.028005f
C2465 VSSD.n23 VSUBS 0.018501f
C2466 VSSD.t385 VSUBS 0.024414f
C2467 VSSD.t846 VSUBS 0.024414f
C2468 VSSD.n24 VSUBS 0.010693f
C2469 VSSD.n25 VSUBS 0.028345f
C2470 VSSD.t848 VSUBS 0.028005f
C2471 VSSD.n27 VSUBS 0.03123f
C2472 VSSD.n28 VSUBS 0.03123f
C2473 VSSD.t1 VSUBS 0.024724f
C2474 VSSD.n30 VSUBS 0.03123f
C2475 VSSD.t1092 VSUBS 0.010396f
C2476 VSSD.n31 VSUBS 0.018748f
C2477 VSSD.n32 VSUBS 0.018565f
C2478 VSSD.n34 VSUBS 0.03123f
C2479 VSSD.t541 VSUBS 0.013879f
C2480 VSSD.n35 VSUBS 0.017846f
C2481 VSSD.n36 VSUBS 0.029746f
C2482 VSSD.t40 VSUBS 0.013879f
C2483 VSSD.n37 VSUBS 0.017846f
C2484 VSSD.n38 VSUBS 0.011061f
C2485 VSSD.n39 VSUBS 0.03123f
C2486 VSSD.t1064 VSUBS 0.010396f
C2487 VSSD.n40 VSUBS 0.018748f
C2488 VSSD.t777 VSUBS 0.024724f
C2489 VSSD.n41 VSUBS 0.036733f
C2490 VSSD.n42 VSUBS 0.03123f
C2491 VSSD.t815 VSUBS 0.028005f
C2492 VSSD.n44 VSUBS 0.018501f
C2493 VSSD.t817 VSUBS 0.024414f
C2494 VSSD.t554 VSUBS 0.024414f
C2495 VSSD.n45 VSUBS 0.010693f
C2496 VSSD.n46 VSUBS 0.028345f
C2497 VSSD.t181 VSUBS 0.028005f
C2498 VSSD.n48 VSUBS 0.03123f
C2499 VSSD.n49 VSUBS 0.03123f
C2500 VSSD.t657 VSUBS 0.024724f
C2501 VSSD.n51 VSUBS 0.03123f
C2502 VSSD.t1068 VSUBS 0.010396f
C2503 VSSD.n52 VSUBS 0.018748f
C2504 VSSD.n53 VSUBS 0.018565f
C2505 VSSD.n55 VSUBS 0.03123f
C2506 VSSD.t702 VSUBS 0.013879f
C2507 VSSD.n56 VSUBS 0.017846f
C2508 VSSD.n57 VSUBS 0.029746f
C2509 VSSD.t196 VSUBS 0.013879f
C2510 VSSD.n58 VSUBS 0.017846f
C2511 VSSD.n59 VSUBS 0.011061f
C2512 VSSD.n60 VSUBS 0.03123f
C2513 VSSD.t1044 VSUBS 0.010396f
C2514 VSSD.n61 VSUBS 0.018748f
C2515 VSSD.t526 VSUBS 0.024724f
C2516 VSSD.n62 VSUBS 0.036733f
C2517 VSSD.n63 VSUBS 0.03123f
C2518 VSSD.t990 VSUBS 0.028005f
C2519 VSSD.n65 VSUBS 0.018501f
C2520 VSSD.t992 VSUBS 0.024414f
C2521 VSSD.t1137 VSUBS 0.024414f
C2522 VSSD.n66 VSUBS 0.010693f
C2523 VSSD.n67 VSUBS 0.028345f
C2524 VSSD.t1139 VSUBS 0.028005f
C2525 VSSD.n69 VSUBS 0.03123f
C2526 VSSD.n70 VSUBS 0.03123f
C2527 VSSD.t545 VSUBS 0.024724f
C2528 VSSD.n72 VSUBS 0.03123f
C2529 VSSD.t1105 VSUBS 0.010396f
C2530 VSSD.n73 VSUBS 0.018748f
C2531 VSSD.n74 VSUBS 0.018565f
C2532 VSSD.n76 VSUBS 0.03123f
C2533 VSSD.t412 VSUBS 0.013879f
C2534 VSSD.n77 VSUBS 0.017846f
C2535 VSSD.n78 VSUBS 0.029746f
C2536 VSSD.t718 VSUBS 0.013879f
C2537 VSSD.n79 VSUBS 0.017846f
C2538 VSSD.n80 VSUBS 0.011061f
C2539 VSSD.n81 VSUBS 0.03123f
C2540 VSSD.t1108 VSUBS 0.010396f
C2541 VSSD.n82 VSUBS 0.018748f
C2542 VSSD.t255 VSUBS 0.024724f
C2543 VSSD.n83 VSUBS 0.036733f
C2544 VSSD.n84 VSUBS 0.03123f
C2545 VSSD.t789 VSUBS 0.028005f
C2546 VSSD.n86 VSUBS 0.018501f
C2547 VSSD.t974 VSUBS 0.024414f
C2548 VSSD.t220 VSUBS 0.024414f
C2549 VSSD.n87 VSUBS 0.010693f
C2550 VSSD.t218 VSUBS 0.028005f
C2551 VSSD.n88 VSUBS 0.03344f
C2552 VSSD.n90 VSUBS 0.03123f
C2553 VSSD.t1110 VSUBS 0.010396f
C2554 VSSD.n91 VSUBS 0.018748f
C2555 VSSD.n92 VSUBS 0.018565f
C2556 VSSD.n93 VSUBS 0.03123f
C2557 VSSD.n95 VSUBS 0.03123f
C2558 VSSD.t1003 VSUBS 0.013879f
C2559 VSSD.n96 VSUBS 0.017846f
C2560 VSSD.n97 VSUBS 0.029746f
C2561 VSSD.n98 VSUBS 0.011061f
C2562 VSSD.n99 VSUBS 0.03123f
C2563 VSSD.t12 VSUBS 0.024724f
C2564 VSSD.n100 VSUBS 0.036733f
C2565 VSSD.n101 VSUBS 0.03123f
C2566 VSSD.n103 VSUBS 0.03123f
C2567 VSSD.n105 VSUBS 0.03123f
C2568 VSSD.n106 VSUBS 0.01373f
C2569 VSSD.n107 VSUBS 0.030584f
C2570 VSSD.n108 VSUBS 0.01373f
C2571 VSSD.n109 VSUBS 0.036114f
C2572 VSSD.n110 VSUBS 0.214581f
C2573 VSSD.n111 VSUBS 0.971351f
C2574 VSSD.n112 VSUBS 1.71988f
C2575 VSSD.n113 VSUBS 0.821251f
C2576 VSSD.n114 VSUBS 0.03123f
C2577 VSSD.t507 VSUBS 0.022291f
C2578 VSSD.t617 VSUBS 0.022309f
C2579 VSSD.n115 VSUBS 0.011262f
C2580 VSSD.n116 VSUBS 0.03123f
C2581 VSSD.n117 VSUBS 0.013217f
C2582 VSSD.t175 VSUBS 0.022003f
C2583 VSSD.n118 VSUBS 0.028916f
C2584 VSSD.t163 VSUBS 0.021956f
C2585 VSSD.n119 VSUBS 0.029108f
C2586 VSSD.n120 VSUBS 0.03123f
C2587 VSSD.t413 VSUBS 0.575862f
C2588 VSSD.t466 VSUBS 0.902264f
C2589 VSSD.t346 VSUBS 0.678213f
C2590 VSSD.t212 VSUBS 0.767816f
C2591 VSSD.t1184 VSUBS 0.767816f
C2592 VSSD.t158 VSUBS 0.767816f
C2593 VSSD.t1182 VSUBS 0.767816f
C2594 VSSD.t210 VSUBS 0.767816f
C2595 VSSD.t160 VSUBS 1.0329f
C2596 VSSD.t1014 VSUBS 1.30254f
C2597 VSSD.n122 VSUBS 0.011835f
C2598 VSSD.t251 VSUBS 0.023899f
C2599 VSSD.n123 VSUBS 0.037275f
C2600 VSSD.n124 VSUBS 0.03123f
C2601 VSSD.n126 VSUBS 0.015053f
C2602 VSSD.t688 VSUBS 0.024724f
C2603 VSSD.n127 VSUBS 0.03123f
C2604 VSSD.n128 VSUBS 0.021146f
C2605 VSSD.n129 VSUBS 0.03123f
C2606 VSSD.n130 VSUBS 0.021146f
C2607 VSSD.n131 VSUBS 0.03123f
C2608 VSSD.t1123 VSUBS 0.010396f
C2609 VSSD.n132 VSUBS 0.018413f
C2610 VSSD.n133 VSUBS 0.021146f
C2611 VSSD.n134 VSUBS 0.03123f
C2612 VSSD.t153 VSUBS 0.027635f
C2613 VSSD.t407 VSUBS 0.023899f
C2614 VSSD.n135 VSUBS 0.037275f
C2615 VSSD.n136 VSUBS 0.022892f
C2616 VSSD.n137 VSUBS 0.03123f
C2617 VSSD.n138 VSUBS 0.021146f
C2618 VSSD.n139 VSUBS 0.03123f
C2619 VSSD.n140 VSUBS 0.012984f
C2620 VSSD.n141 VSUBS 0.03123f
C2621 VSSD.n142 VSUBS 0.021146f
C2622 VSSD.n143 VSUBS 0.03123f
C2623 VSSD.t279 VSUBS 0.010396f
C2624 VSSD.n144 VSUBS 0.018413f
C2625 VSSD.n145 VSUBS 0.021146f
C2626 VSSD.n146 VSUBS 0.03123f
C2627 VSSD.t56 VSUBS 0.027635f
C2628 VSSD.t54 VSUBS 0.023899f
C2629 VSSD.n147 VSUBS 0.017122f
C2630 VSSD.n148 VSUBS 0.03123f
C2631 VSSD.n150 VSUBS 0.015053f
C2632 VSSD.t118 VSUBS 0.024724f
C2633 VSSD.n151 VSUBS 0.03123f
C2634 VSSD.n152 VSUBS 0.021146f
C2635 VSSD.n153 VSUBS 0.03123f
C2636 VSSD.n154 VSUBS 0.021146f
C2637 VSSD.n155 VSUBS 0.03123f
C2638 VSSD.t692 VSUBS 0.010396f
C2639 VSSD.n156 VSUBS 0.018413f
C2640 VSSD.n157 VSUBS 0.021146f
C2641 VSSD.n158 VSUBS 0.03123f
C2642 VSSD.t358 VSUBS 0.027635f
C2643 VSSD.t723 VSUBS 0.023899f
C2644 VSSD.n159 VSUBS 0.043227f
C2645 VSSD.t295 VSUBS 0.022506f
C2646 VSSD.n160 VSUBS 0.047644f
C2647 VSSD.t226 VSUBS 0.023899f
C2648 VSSD.n161 VSUBS 0.037275f
C2649 VSSD.n162 VSUBS 0.03123f
C2650 VSSD.t224 VSUBS 0.027635f
C2651 VSSD.n163 VSUBS 0.021146f
C2652 VSSD.n164 VSUBS 0.03123f
C2653 VSSD.t1170 VSUBS 0.010396f
C2654 VSSD.n165 VSUBS 0.018413f
C2655 VSSD.n166 VSUBS 0.021146f
C2656 VSSD.n167 VSUBS 0.03123f
C2657 VSSD.t369 VSUBS 0.013879f
C2658 VSSD.n168 VSUBS 0.018245f
C2659 VSSD.n169 VSUBS 0.021146f
C2660 VSSD.n170 VSUBS 0.03123f
C2661 VSSD.n171 VSUBS 0.015053f
C2662 VSSD.n172 VSUBS 0.03123f
C2663 VSSD.t332 VSUBS 0.024724f
C2664 VSSD.n174 VSUBS 0.022624f
C2665 VSSD.n175 VSUBS 0.011262f
C2666 VSSD.n176 VSUBS 0.03123f
C2667 VSSD.n177 VSUBS 0.03123f
C2668 VSSD.t101 VSUBS 0.023899f
C2669 VSSD.n178 VSUBS 0.037275f
C2670 VSSD.t103 VSUBS 0.027635f
C2671 VSSD.n179 VSUBS 0.021146f
C2672 VSSD.n180 VSUBS 0.03123f
C2673 VSSD.t731 VSUBS 0.010396f
C2674 VSSD.n181 VSUBS 0.018413f
C2675 VSSD.n182 VSUBS 0.021146f
C2676 VSSD.n183 VSUBS 0.03123f
C2677 VSSD.t360 VSUBS 0.013879f
C2678 VSSD.n184 VSUBS 0.018245f
C2679 VSSD.n185 VSUBS 0.021146f
C2680 VSSD.n186 VSUBS 0.03123f
C2681 VSSD.n187 VSUBS 0.015053f
C2682 VSSD.n188 VSUBS 0.03123f
C2683 VSSD.t642 VSUBS 0.024724f
C2684 VSSD.n190 VSUBS 0.022624f
C2685 VSSD.n191 VSUBS 0.011262f
C2686 VSSD.n192 VSUBS 0.03123f
C2687 VSSD.n193 VSUBS 0.03123f
C2688 VSSD.t484 VSUBS 0.023899f
C2689 VSSD.n194 VSUBS 0.037275f
C2690 VSSD.t750 VSUBS 0.027635f
C2691 VSSD.n195 VSUBS 0.021146f
C2692 VSSD.n196 VSUBS 0.03123f
C2693 VSSD.t698 VSUBS 0.010396f
C2694 VSSD.n197 VSUBS 0.018413f
C2695 VSSD.n198 VSUBS 0.021146f
C2696 VSSD.n199 VSUBS 0.03123f
C2697 VSSD.t706 VSUBS 0.013879f
C2698 VSSD.n200 VSUBS 0.018245f
C2699 VSSD.n201 VSUBS 0.021146f
C2700 VSSD.n202 VSUBS 0.03123f
C2701 VSSD.n203 VSUBS 0.015053f
C2702 VSSD.n204 VSUBS 0.03123f
C2703 VSSD.t588 VSUBS 0.024724f
C2704 VSSD.n206 VSUBS 0.022624f
C2705 VSSD.t294 VSUBS 0.125098f
C2706 VSSD.t880 VSUBS 0.902264f
C2707 VSSD.t441 VSUBS 2.0528f
C2708 VSSD.t687 VSUBS 2.11941f
C2709 VSSD.t417 VSUBS 1.15659f
C2710 VSSD.t771 VSUBS 1.58653f
C2711 VSSD.t741 VSUBS 1.4412f
C2712 VSSD.t826 VSUBS 1.23532f
C2713 VSSD.t680 VSUBS 1.39881f
C2714 VSSD.t772 VSUBS 1.25954f
C2715 VSSD.t416 VSUBS 1.24137f
C2716 VSSD.t114 VSUBS 1.48359f
C2717 VSSD.t1122 VSUBS 1.45331f
C2718 VSSD.t296 VSUBS 1.81059f
C2719 VSSD.t152 VSUBS 1.7682f
C2720 VSSD.t406 VSUBS 1.30193f
C2721 VSSD.t824 VSUBS 0.902264f
C2722 VSSD.t322 VSUBS 2.0528f
C2723 VSSD.t1118 VSUBS 2.11941f
C2724 VSSD.t321 VSUBS 1.15659f
C2725 VSSD.t6 VSUBS 1.58653f
C2726 VSSD.t156 VSUBS 1.4412f
C2727 VSSD.t513 VSUBS 1.23532f
C2728 VSSD.t18 VSUBS 1.39881f
C2729 VSSD.t57 VSUBS 1.25954f
C2730 VSSD.t17 VSUBS 1.24137f
C2731 VSSD.t580 VSUBS 1.48359f
C2732 VSSD.t278 VSUBS 1.45331f
C2733 VSSD.t627 VSUBS 1.81059f
C2734 VSSD.t55 VSUBS 1.7682f
C2735 VSSD.t53 VSUBS 1.30193f
C2736 VSSD.t805 VSUBS 0.902264f
C2737 VSSD.t235 VSUBS 2.0528f
C2738 VSSD.t117 VSUBS 2.11941f
C2739 VSSD.t923 VSUBS 1.15659f
C2740 VSSD.t338 VSUBS 1.58653f
C2741 VSSD.t981 VSUBS 1.4412f
C2742 VSSD.t15 VSUBS 1.23532f
C2743 VSSD.t861 VSUBS 1.39881f
C2744 VSSD.t337 VSUBS 1.25954f
C2745 VSSD.t237 VSUBS 1.24137f
C2746 VSSD.t355 VSUBS 1.48359f
C2747 VSSD.t691 VSUBS 1.45331f
C2748 VSSD.t555 VSUBS 1.81059f
C2749 VSSD.t357 VSUBS 1.7682f
C2750 VSSD.t722 VSUBS 4.45446f
C2751 VSSD.n207 VSUBS 0.101664f
C2752 VSSD.n208 VSUBS 0.046796f
C2753 VSSD.t225 VSUBS 0.197283f
C2754 VSSD.t223 VSUBS 0.26794f
C2755 VSSD.t390 VSUBS 0.274362f
C2756 VSSD.t1169 VSUBS 0.220221f
C2757 VSSD.t221 VSUBS 0.224811f
C2758 VSSD.t948 VSUBS 0.188107f
C2759 VSSD.t592 VSUBS 0.190858f
C2760 VSSD.t368 VSUBS 0.211965f
C2761 VSSD.t515 VSUBS 0.187191f
C2762 VSSD.t126 VSUBS 0.21839f
C2763 VSSD.t1135 VSUBS 0.240412f
C2764 VSSD.t1005 VSUBS 0.17526f
C2765 VSSD.t331 VSUBS 0.321158f
C2766 VSSD.t946 VSUBS 0.311066f
C2767 VSSD.t307 VSUBS 0.136721f
C2768 VSSD.t100 VSUBS 0.197283f
C2769 VSSD.t102 VSUBS 0.26794f
C2770 VSSD.t99 VSUBS 0.274362f
C2771 VSSD.t730 VSUBS 0.220221f
C2772 VSSD.t1133 VSUBS 0.224811f
C2773 VSSD.t317 VSUBS 0.188107f
C2774 VSSD.t446 VSUBS 0.190858f
C2775 VSSD.t359 VSUBS 0.211965f
C2776 VSSD.t689 VSUBS 0.187191f
C2777 VSSD.t528 VSUBS 0.21839f
C2778 VSSD.t445 VSUBS 0.240412f
C2779 VSSD.t318 VSUBS 0.17526f
C2780 VSSD.t641 VSUBS 0.321158f
C2781 VSSD.t66 VSUBS 0.311066f
C2782 VSSD.t882 VSUBS 0.136721f
C2783 VSSD.t483 VSUBS 0.197283f
C2784 VSSD.t749 VSUBS 0.26794f
C2785 VSSD.t770 VSUBS 0.274362f
C2786 VSSD.t697 VSUBS 0.220221f
C2787 VSSD.t747 VSUBS 0.224811f
C2788 VSSD.t1128 VSUBS 0.188107f
C2789 VSSD.t501 VSUBS 0.190858f
C2790 VSSD.t705 VSUBS 0.211965f
C2791 VSSD.t276 VSUBS 0.187191f
C2792 VSSD.t700 VSUBS 0.21839f
C2793 VSSD.t500 VSUBS 0.240412f
C2794 VSSD.t675 VSUBS 0.17526f
C2795 VSSD.t587 VSUBS 0.321158f
C2796 VSSD.t676 VSUBS 0.270691f
C2797 VSSD.t468 VSUBS 0.136721f
C2798 VSSD.t830 VSUBS 0.311066f
C2799 VSSD.t1186 VSUBS 0.321158f
C2800 VSSD.t829 VSUBS 0.17526f
C2801 VSSD.t238 VSUBS 0.240412f
C2802 VSSD.t361 VSUBS 0.21839f
C2803 VSSD.t621 VSUBS 0.187191f
C2804 VSSD.t843 VSUBS 0.211965f
C2805 VSSD.t239 VSUBS 0.190858f
C2806 VSSD.t832 VSUBS 0.188107f
C2807 VSSD.t1130 VSUBS 0.224811f
C2808 VSSD.t1171 VSUBS 0.220221f
C2809 VSSD.t1147 VSUBS 0.274362f
C2810 VSSD.t893 VSUBS 0.26794f
C2811 VSSD.t891 VSUBS 0.197283f
C2812 VSSD.t309 VSUBS 0.136721f
C2813 VSSD.t773 VSUBS 0.311066f
C2814 VSSD.t582 VSUBS 0.321158f
C2815 VSSD.t643 VSUBS 0.17526f
C2816 VSSD.t20 VSUBS 0.240412f
C2817 VSSD.t573 VSUBS 0.21839f
C2818 VSSD.t268 VSUBS 0.187191f
C2819 VSSD.t298 VSUBS 0.211965f
C2820 VSSD.t21 VSUBS 0.190858f
C2821 VSSD.t1194 VSUBS 0.188107f
C2822 VSSD.t341 VSUBS 0.224811f
C2823 VSSD.t1175 VSUBS 0.220221f
C2824 VSSD.t504 VSUBS 0.274362f
C2825 VSSD.t462 VSUBS 0.26794f
C2826 VSSD.t460 VSUBS 0.197283f
C2827 VSSD.t558 VSUBS 0.136721f
C2828 VSSD.t427 VSUBS 0.311066f
C2829 VSSD.t785 VSUBS 0.321158f
C2830 VSSD.t535 VSUBS 0.17526f
C2831 VSSD.t956 VSUBS 0.240412f
C2832 VSSD.t319 VSUBS 0.21839f
C2833 VSSD.t1120 VSUBS 0.187191f
C2834 VSSD.t315 VSUBS 0.211965f
C2835 VSSD.t399 VSUBS 0.190858f
C2836 VSSD.t429 VSUBS 0.188107f
C2837 VSSD.t951 VSUBS 0.224811f
C2838 VSSD.t724 VSUBS 0.220221f
C2839 VSSD.t457 VSUBS 0.274362f
C2840 VSSD.t781 VSUBS 0.26794f
C2841 VSSD.t779 VSUBS 0.197283f
C2842 VSSD.t803 VSUBS 0.100017f
C2843 VSSD.n209 VSUBS -0.849272f
C2844 VSSD.n210 VSUBS 0.011262f
C2845 VSSD.n211 VSUBS 0.03123f
C2846 VSSD.n212 VSUBS 0.03123f
C2847 VSSD.t780 VSUBS 0.023899f
C2848 VSSD.n213 VSUBS 0.037275f
C2849 VSSD.t782 VSUBS 0.027635f
C2850 VSSD.n214 VSUBS 0.021146f
C2851 VSSD.n215 VSUBS 0.03123f
C2852 VSSD.t725 VSUBS 0.010396f
C2853 VSSD.n216 VSUBS 0.018413f
C2854 VSSD.n217 VSUBS 0.021146f
C2855 VSSD.n218 VSUBS 0.03123f
C2856 VSSD.t316 VSUBS 0.013879f
C2857 VSSD.n219 VSUBS 0.018245f
C2858 VSSD.n220 VSUBS 0.021146f
C2859 VSSD.n221 VSUBS 0.03123f
C2860 VSSD.n222 VSUBS 0.015053f
C2861 VSSD.n223 VSUBS 0.03123f
C2862 VSSD.t786 VSUBS 0.024724f
C2863 VSSD.n225 VSUBS 0.022624f
C2864 VSSD.n226 VSUBS 0.011262f
C2865 VSSD.n227 VSUBS 0.03123f
C2866 VSSD.n228 VSUBS 0.03123f
C2867 VSSD.t461 VSUBS 0.023899f
C2868 VSSD.n229 VSUBS 0.037275f
C2869 VSSD.t463 VSUBS 0.027635f
C2870 VSSD.n230 VSUBS 0.021146f
C2871 VSSD.n231 VSUBS 0.03123f
C2872 VSSD.t1176 VSUBS 0.010396f
C2873 VSSD.n232 VSUBS 0.018413f
C2874 VSSD.n233 VSUBS 0.021146f
C2875 VSSD.n234 VSUBS 0.03123f
C2876 VSSD.t299 VSUBS 0.013879f
C2877 VSSD.n235 VSUBS 0.018245f
C2878 VSSD.n236 VSUBS 0.021146f
C2879 VSSD.n237 VSUBS 0.03123f
C2880 VSSD.n238 VSUBS 0.015053f
C2881 VSSD.n239 VSUBS 0.03123f
C2882 VSSD.t583 VSUBS 0.024724f
C2883 VSSD.n241 VSUBS 0.022624f
C2884 VSSD.n242 VSUBS 0.011262f
C2885 VSSD.n243 VSUBS 0.03123f
C2886 VSSD.n244 VSUBS 0.03123f
C2887 VSSD.t892 VSUBS 0.023899f
C2888 VSSD.n245 VSUBS 0.037275f
C2889 VSSD.t894 VSUBS 0.027635f
C2890 VSSD.n246 VSUBS 0.021146f
C2891 VSSD.n247 VSUBS 0.03123f
C2892 VSSD.t1172 VSUBS 0.010396f
C2893 VSSD.n248 VSUBS 0.018413f
C2894 VSSD.n249 VSUBS 0.021146f
C2895 VSSD.n250 VSUBS 0.03123f
C2896 VSSD.t844 VSUBS 0.013879f
C2897 VSSD.n251 VSUBS 0.018245f
C2898 VSSD.n252 VSUBS 0.021146f
C2899 VSSD.n253 VSUBS 0.03123f
C2900 VSSD.n254 VSUBS 0.015053f
C2901 VSSD.n255 VSUBS 0.03123f
C2902 VSSD.t1187 VSUBS 0.024724f
C2903 VSSD.n257 VSUBS 0.022624f
C2904 VSSD.n258 VSUBS 0.03123f
C2905 VSSD.n259 VSUBS 0.025373f
C2906 VSSD.n260 VSUBS 0.028587f
C2907 VSSD.n261 VSUBS 0.016086f
C2908 VSSD.n262 VSUBS 0.022892f
C2909 VSSD.n263 VSUBS 0.029102f
C2910 VSSD.n264 VSUBS 0.03123f
C2911 VSSD.n265 VSUBS 0.03123f
C2912 VSSD.n266 VSUBS 0.03123f
C2913 VSSD.n267 VSUBS 0.021146f
C2914 VSSD.n268 VSUBS 0.021146f
C2915 VSSD.n269 VSUBS 0.021146f
C2916 VSSD.n270 VSUBS 0.03123f
C2917 VSSD.n271 VSUBS 0.03123f
C2918 VSSD.n272 VSUBS 0.03123f
C2919 VSSD.n273 VSUBS 0.012984f
C2920 VSSD.n274 VSUBS 0.038003f
C2921 VSSD.n275 VSUBS 0.011146f
C2922 VSSD.n276 VSUBS 0.021146f
C2923 VSSD.n277 VSUBS 0.03123f
C2924 VSSD.n278 VSUBS 0.03123f
C2925 VSSD.n279 VSUBS 0.03123f
C2926 VSSD.n280 VSUBS 0.021146f
C2927 VSSD.n281 VSUBS 0.013561f
C2928 VSSD.n282 VSUBS 0.021657f
C2929 VSSD.n283 VSUBS 0.018158f
C2930 VSSD.n284 VSUBS 0.03123f
C2931 VSSD.n285 VSUBS 0.03123f
C2932 VSSD.n286 VSUBS 0.03123f
C2933 VSSD.n287 VSUBS 0.021146f
C2934 VSSD.n288 VSUBS 0.011033f
C2935 VSSD.n289 VSUBS 0.032298f
C2936 VSSD.n290 VSUBS 0.019996f
C2937 VSSD.n291 VSUBS 0.03123f
C2938 VSSD.n292 VSUBS 0.023423f
C2939 VSSD.n293 VSUBS 0.018501f
C2940 VSSD.n294 VSUBS 0.017122f
C2941 VSSD.n295 VSUBS 0.022892f
C2942 VSSD.n296 VSUBS 0.016086f
C2943 VSSD.n297 VSUBS 0.022892f
C2944 VSSD.n298 VSUBS 0.029102f
C2945 VSSD.n299 VSUBS 0.03123f
C2946 VSSD.n300 VSUBS 0.03123f
C2947 VSSD.n301 VSUBS 0.03123f
C2948 VSSD.n302 VSUBS 0.021146f
C2949 VSSD.n303 VSUBS 0.021146f
C2950 VSSD.n304 VSUBS 0.021146f
C2951 VSSD.n305 VSUBS 0.03123f
C2952 VSSD.n306 VSUBS 0.03123f
C2953 VSSD.n307 VSUBS 0.03123f
C2954 VSSD.n308 VSUBS 0.012984f
C2955 VSSD.n309 VSUBS 0.038003f
C2956 VSSD.n310 VSUBS 0.011146f
C2957 VSSD.n311 VSUBS 0.021146f
C2958 VSSD.n312 VSUBS 0.03123f
C2959 VSSD.n313 VSUBS 0.03123f
C2960 VSSD.n314 VSUBS 0.03123f
C2961 VSSD.n315 VSUBS 0.021146f
C2962 VSSD.n316 VSUBS 0.013561f
C2963 VSSD.n317 VSUBS 0.021657f
C2964 VSSD.n318 VSUBS 0.018158f
C2965 VSSD.n319 VSUBS 0.03123f
C2966 VSSD.n320 VSUBS 0.03123f
C2967 VSSD.n321 VSUBS 0.03123f
C2968 VSSD.n322 VSUBS 0.021146f
C2969 VSSD.n323 VSUBS 0.011033f
C2970 VSSD.n324 VSUBS 0.032298f
C2971 VSSD.n325 VSUBS 0.019996f
C2972 VSSD.n326 VSUBS 0.03123f
C2973 VSSD.n327 VSUBS 0.023423f
C2974 VSSD.n328 VSUBS 0.018501f
C2975 VSSD.n329 VSUBS 0.017122f
C2976 VSSD.n330 VSUBS 0.022892f
C2977 VSSD.n331 VSUBS 0.016086f
C2978 VSSD.n332 VSUBS 0.022892f
C2979 VSSD.n333 VSUBS 0.029102f
C2980 VSSD.n334 VSUBS 0.03123f
C2981 VSSD.n335 VSUBS 0.03123f
C2982 VSSD.n336 VSUBS 0.03123f
C2983 VSSD.n337 VSUBS 0.021146f
C2984 VSSD.n338 VSUBS 0.021146f
C2985 VSSD.n339 VSUBS 0.021146f
C2986 VSSD.n340 VSUBS 0.03123f
C2987 VSSD.n341 VSUBS 0.03123f
C2988 VSSD.n342 VSUBS 0.03123f
C2989 VSSD.n343 VSUBS 0.012984f
C2990 VSSD.n344 VSUBS 0.038003f
C2991 VSSD.n345 VSUBS 0.011146f
C2992 VSSD.n346 VSUBS 0.021146f
C2993 VSSD.n347 VSUBS 0.03123f
C2994 VSSD.n348 VSUBS 0.03123f
C2995 VSSD.n349 VSUBS 0.03123f
C2996 VSSD.n350 VSUBS 0.021146f
C2997 VSSD.n351 VSUBS 0.013561f
C2998 VSSD.n352 VSUBS 0.021657f
C2999 VSSD.n353 VSUBS 0.018158f
C3000 VSSD.n354 VSUBS 0.03123f
C3001 VSSD.n355 VSUBS 0.03123f
C3002 VSSD.n356 VSUBS 0.03123f
C3003 VSSD.n357 VSUBS 0.021146f
C3004 VSSD.n358 VSUBS 0.011033f
C3005 VSSD.n359 VSUBS 0.032298f
C3006 VSSD.n360 VSUBS 0.019996f
C3007 VSSD.n361 VSUBS 0.03123f
C3008 VSSD.n362 VSUBS 0.023423f
C3009 VSSD.n363 VSUBS 0.018501f
C3010 VSSD.n364 VSUBS 0.017122f
C3011 VSSD.n365 VSUBS -0.476391f
C3012 VSSD.n366 VSUBS 0.016086f
C3013 VSSD.n367 VSUBS 0.022892f
C3014 VSSD.n368 VSUBS 0.029102f
C3015 VSSD.n369 VSUBS 0.03123f
C3016 VSSD.n370 VSUBS 0.03123f
C3017 VSSD.n371 VSUBS 0.03123f
C3018 VSSD.n372 VSUBS 0.021146f
C3019 VSSD.n373 VSUBS 0.021146f
C3020 VSSD.n374 VSUBS 0.021146f
C3021 VSSD.n375 VSUBS 0.03123f
C3022 VSSD.n376 VSUBS 0.03123f
C3023 VSSD.n377 VSUBS 0.03123f
C3024 VSSD.n378 VSUBS 0.012984f
C3025 VSSD.n379 VSUBS 0.038003f
C3026 VSSD.n380 VSUBS 0.011146f
C3027 VSSD.n381 VSUBS 0.021146f
C3028 VSSD.n382 VSUBS 0.03123f
C3029 VSSD.n383 VSUBS 0.03123f
C3030 VSSD.n384 VSUBS 0.03123f
C3031 VSSD.n385 VSUBS 0.021146f
C3032 VSSD.n386 VSUBS 0.013561f
C3033 VSSD.n387 VSUBS 0.021657f
C3034 VSSD.n388 VSUBS 0.018158f
C3035 VSSD.n389 VSUBS 0.03123f
C3036 VSSD.n390 VSUBS 0.03123f
C3037 VSSD.n391 VSUBS 0.03123f
C3038 VSSD.n392 VSUBS 0.021146f
C3039 VSSD.n393 VSUBS 0.011033f
C3040 VSSD.n394 VSUBS 0.032298f
C3041 VSSD.n395 VSUBS 0.019996f
C3042 VSSD.n396 VSUBS 0.03123f
C3043 VSSD.n397 VSUBS 0.023423f
C3044 VSSD.n398 VSUBS 0.018501f
C3045 VSSD.n399 VSUBS 0.017122f
C3046 VSSD.n400 VSUBS 0.022892f
C3047 VSSD.n401 VSUBS 0.016086f
C3048 VSSD.n402 VSUBS 0.022892f
C3049 VSSD.n403 VSUBS 0.029102f
C3050 VSSD.n404 VSUBS 0.03123f
C3051 VSSD.n405 VSUBS 0.03123f
C3052 VSSD.n406 VSUBS 0.03123f
C3053 VSSD.n407 VSUBS 0.021146f
C3054 VSSD.n408 VSUBS 0.021146f
C3055 VSSD.n409 VSUBS 0.021146f
C3056 VSSD.n410 VSUBS 0.03123f
C3057 VSSD.n411 VSUBS 0.03123f
C3058 VSSD.n412 VSUBS 0.03123f
C3059 VSSD.n413 VSUBS 0.012984f
C3060 VSSD.n414 VSUBS 0.038003f
C3061 VSSD.n415 VSUBS 0.011146f
C3062 VSSD.n416 VSUBS 0.021146f
C3063 VSSD.n417 VSUBS 0.03123f
C3064 VSSD.n418 VSUBS 0.03123f
C3065 VSSD.n419 VSUBS 0.03123f
C3066 VSSD.n420 VSUBS 0.021146f
C3067 VSSD.n421 VSUBS 0.013561f
C3068 VSSD.n422 VSUBS 0.021657f
C3069 VSSD.n423 VSUBS 0.018158f
C3070 VSSD.n424 VSUBS 0.03123f
C3071 VSSD.n425 VSUBS 0.03123f
C3072 VSSD.n426 VSUBS 0.03123f
C3073 VSSD.n427 VSUBS 0.021146f
C3074 VSSD.n428 VSUBS 0.011033f
C3075 VSSD.n429 VSUBS 0.032298f
C3076 VSSD.n430 VSUBS 0.019996f
C3077 VSSD.n431 VSUBS 0.03123f
C3078 VSSD.n432 VSUBS 0.023423f
C3079 VSSD.n433 VSUBS 0.018501f
C3080 VSSD.n434 VSUBS 0.017122f
C3081 VSSD.n435 VSUBS 0.022892f
C3082 VSSD.n436 VSUBS 0.016086f
C3083 VSSD.n437 VSUBS 0.022892f
C3084 VSSD.n438 VSUBS 0.029102f
C3085 VSSD.n439 VSUBS 0.03123f
C3086 VSSD.n440 VSUBS 0.03123f
C3087 VSSD.n441 VSUBS 0.03123f
C3088 VSSD.n442 VSUBS 0.021146f
C3089 VSSD.n443 VSUBS 0.021146f
C3090 VSSD.n444 VSUBS 0.021146f
C3091 VSSD.n445 VSUBS 0.03123f
C3092 VSSD.n446 VSUBS 0.03123f
C3093 VSSD.n447 VSUBS 0.03123f
C3094 VSSD.n448 VSUBS 0.012984f
C3095 VSSD.n449 VSUBS 0.038003f
C3096 VSSD.n450 VSUBS 0.011146f
C3097 VSSD.n451 VSUBS 0.021146f
C3098 VSSD.n452 VSUBS 0.03123f
C3099 VSSD.n453 VSUBS 0.03123f
C3100 VSSD.n454 VSUBS 0.03123f
C3101 VSSD.n455 VSUBS 0.021146f
C3102 VSSD.n456 VSUBS 0.013561f
C3103 VSSD.n457 VSUBS 0.021657f
C3104 VSSD.n458 VSUBS 0.018158f
C3105 VSSD.n459 VSUBS 0.03123f
C3106 VSSD.n460 VSUBS 0.03123f
C3107 VSSD.n461 VSUBS 0.03123f
C3108 VSSD.n462 VSUBS 0.021146f
C3109 VSSD.n463 VSUBS 0.011033f
C3110 VSSD.n464 VSUBS 0.032298f
C3111 VSSD.n465 VSUBS 0.019996f
C3112 VSSD.n466 VSUBS 0.03123f
C3113 VSSD.n467 VSUBS 0.023423f
C3114 VSSD.n468 VSUBS 0.011262f
C3115 VSSD.n469 VSUBS 0.015283f
C3116 VSSD.n470 VSUBS 0.024879f
C3117 VSSD.n471 VSUBS 0.243513f
C3118 VSSD.t1015 VSUBS 0.022506f
C3119 VSSD.n472 VSUBS 0.047644f
C3120 VSSD.t161 VSUBS 0.021939f
C3121 VSSD.n473 VSUBS 0.032378f
C3122 VSSD.n474 VSUBS 0.03123f
C3123 VSSD.n475 VSUBS 0.013217f
C3124 VSSD.n476 VSUBS 0.013217f
C3125 VSSD.n477 VSUBS 0.020824f
C3126 VSSD.n478 VSUBS 0.03123f
C3127 VSSD.n479 VSUBS 0.013217f
C3128 VSSD.n480 VSUBS 0.020824f
C3129 VSSD.n481 VSUBS 0.018501f
C3130 VSSD.n482 VSUBS 0.011375f
C3131 VSSD.n483 VSUBS 0.03123f
C3132 VSSD.n484 VSUBS 0.03123f
C3133 VSSD.n485 VSUBS 0.019303f
C3134 VSSD.n486 VSUBS 0.020824f
C3135 VSSD.n487 VSUBS 0.011605f
C3136 VSSD.n488 VSUBS 0.019767f
C3137 VSSD.n489 VSUBS 0.03123f
C3138 VSSD.n490 VSUBS 0.023423f
C3139 VSSD.n491 VSUBS 0.011952f
C3140 VSSD.n492 VSUBS 0.015283f
C3141 VSSD.n493 VSUBS 0.024879f
C3142 VSSD.n494 VSUBS 1.53123f
C3143 VSSD.n495 VSUBS 1.82097f
C3144 VSSD.n496 VSUBS 0.11804f
C3145 VSSD.n497 VSUBS 0.03123f
C3146 VSSD.n498 VSUBS 0.019996f
C3147 VSSD.n499 VSUBS 0.032298f
C3148 VSSD.n500 VSUBS 0.011033f
C3149 VSSD.n501 VSUBS 0.021146f
C3150 VSSD.n502 VSUBS 0.03123f
C3151 VSSD.n503 VSUBS 0.03123f
C3152 VSSD.n504 VSUBS 0.03123f
C3153 VSSD.n505 VSUBS 0.018158f
C3154 VSSD.n506 VSUBS 0.021657f
C3155 VSSD.n507 VSUBS 0.013561f
C3156 VSSD.n508 VSUBS 0.021146f
C3157 VSSD.n509 VSUBS 0.03123f
C3158 VSSD.n510 VSUBS 0.03123f
C3159 VSSD.n511 VSUBS 0.03123f
C3160 VSSD.n512 VSUBS 0.021146f
C3161 VSSD.n513 VSUBS 0.011146f
C3162 VSSD.t862 VSUBS 0.013879f
C3163 VSSD.n514 VSUBS 0.018245f
C3164 VSSD.n515 VSUBS 0.038003f
C3165 VSSD.n516 VSUBS 0.012984f
C3166 VSSD.n517 VSUBS 0.03123f
C3167 VSSD.n518 VSUBS 0.03123f
C3168 VSSD.n519 VSUBS 0.03123f
C3169 VSSD.n520 VSUBS 0.021146f
C3170 VSSD.n521 VSUBS 0.021146f
C3171 VSSD.n522 VSUBS 0.021146f
C3172 VSSD.n523 VSUBS 0.03123f
C3173 VSSD.n524 VSUBS 0.03123f
C3174 VSSD.n525 VSUBS 0.03123f
C3175 VSSD.n526 VSUBS 0.029102f
C3176 VSSD.n527 VSUBS 0.022892f
C3177 VSSD.n528 VSUBS 0.016086f
C3178 VSSD.n529 VSUBS 0.022892f
C3179 VSSD.n530 VSUBS 0.022624f
C3180 VSSD.n531 VSUBS 0.03123f
C3181 VSSD.n532 VSUBS 0.018501f
C3182 VSSD.n533 VSUBS 0.023423f
C3183 VSSD.n534 VSUBS 0.011262f
C3184 VSSD.n535 VSUBS 0.037275f
C3185 VSSD.n536 VSUBS 0.019996f
C3186 VSSD.n537 VSUBS 0.032298f
C3187 VSSD.n538 VSUBS 0.011033f
C3188 VSSD.n539 VSUBS 0.03123f
C3189 VSSD.n540 VSUBS 0.03123f
C3190 VSSD.n541 VSUBS 0.03123f
C3191 VSSD.n542 VSUBS 0.021146f
C3192 VSSD.n543 VSUBS 0.018158f
C3193 VSSD.n544 VSUBS 0.021657f
C3194 VSSD.n545 VSUBS 0.013561f
C3195 VSSD.n546 VSUBS 0.03123f
C3196 VSSD.n547 VSUBS 0.03123f
C3197 VSSD.n548 VSUBS 0.03123f
C3198 VSSD.n549 VSUBS 0.021146f
C3199 VSSD.n550 VSUBS 0.021146f
C3200 VSSD.t19 VSUBS 0.013879f
C3201 VSSD.n551 VSUBS 0.018245f
C3202 VSSD.n552 VSUBS 0.038003f
C3203 VSSD.n553 VSUBS 0.011146f
C3204 VSSD.n554 VSUBS 0.03123f
C3205 VSSD.n555 VSUBS 0.03123f
C3206 VSSD.n556 VSUBS 0.03123f
C3207 VSSD.n557 VSUBS 0.021146f
C3208 VSSD.n558 VSUBS 0.021146f
C3209 VSSD.n559 VSUBS 0.021146f
C3210 VSSD.n560 VSUBS 0.03123f
C3211 VSSD.n561 VSUBS 0.03123f
C3212 VSSD.n562 VSUBS 0.03123f
C3213 VSSD.n563 VSUBS 0.015053f
C3214 VSSD.t1119 VSUBS 0.024724f
C3215 VSSD.n564 VSUBS 0.029102f
C3216 VSSD.n565 VSUBS 0.022892f
C3217 VSSD.n566 VSUBS 0.016086f
C3218 VSSD.n567 VSUBS 0.03123f
C3219 VSSD.n569 VSUBS 0.022624f
C3220 VSSD.n570 VSUBS 0.03123f
C3221 VSSD.n571 VSUBS 0.018501f
C3222 VSSD.n572 VSUBS 0.017122f
C3223 VSSD.n573 VSUBS 0.011262f
C3224 VSSD.n574 VSUBS 0.023423f
C3225 VSSD.n575 VSUBS 0.03123f
C3226 VSSD.n576 VSUBS 0.019996f
C3227 VSSD.n577 VSUBS 0.032298f
C3228 VSSD.n578 VSUBS 0.011033f
C3229 VSSD.n579 VSUBS 0.021146f
C3230 VSSD.n580 VSUBS 0.03123f
C3231 VSSD.n581 VSUBS 0.03123f
C3232 VSSD.n582 VSUBS 0.03123f
C3233 VSSD.n583 VSUBS 0.018158f
C3234 VSSD.n584 VSUBS 0.021657f
C3235 VSSD.n585 VSUBS 0.013561f
C3236 VSSD.n586 VSUBS 0.021146f
C3237 VSSD.n587 VSUBS 0.03123f
C3238 VSSD.n588 VSUBS 0.03123f
C3239 VSSD.n589 VSUBS 0.03123f
C3240 VSSD.n590 VSUBS 0.021146f
C3241 VSSD.n591 VSUBS 0.011146f
C3242 VSSD.t681 VSUBS 0.013879f
C3243 VSSD.n592 VSUBS 0.018245f
C3244 VSSD.n593 VSUBS 0.038003f
C3245 VSSD.n594 VSUBS 0.012984f
C3246 VSSD.n595 VSUBS 0.03123f
C3247 VSSD.n596 VSUBS 0.03123f
C3248 VSSD.n597 VSUBS 0.03123f
C3249 VSSD.n598 VSUBS 0.021146f
C3250 VSSD.n599 VSUBS 0.021146f
C3251 VSSD.n600 VSUBS 0.021146f
C3252 VSSD.n601 VSUBS 0.03123f
C3253 VSSD.n602 VSUBS 0.03123f
C3254 VSSD.n603 VSUBS 0.03123f
C3255 VSSD.n604 VSUBS 0.029102f
C3256 VSSD.n605 VSUBS 0.022892f
C3257 VSSD.n606 VSUBS 0.016086f
C3258 VSSD.n607 VSUBS 0.022892f
C3259 VSSD.n608 VSUBS 0.022624f
C3260 VSSD.n609 VSUBS 0.03123f
C3261 VSSD.n610 VSUBS 0.018501f
C3262 VSSD.n611 VSUBS 0.03123f
C3263 VSSD.t809 VSUBS 0.027635f
C3264 VSSD.n612 VSUBS 0.021146f
C3265 VSSD.n613 VSUBS 0.03123f
C3266 VSSD.t696 VSUBS 0.010396f
C3267 VSSD.n614 VSUBS 0.018413f
C3268 VSSD.n615 VSUBS 0.021146f
C3269 VSSD.n616 VSUBS 0.03123f
C3270 VSSD.t929 VSUBS 0.013879f
C3271 VSSD.n617 VSUBS 0.018245f
C3272 VSSD.n618 VSUBS 0.021146f
C3273 VSSD.n619 VSUBS 0.03123f
C3274 VSSD.n620 VSUBS 0.015053f
C3275 VSSD.n621 VSUBS 0.03123f
C3276 VSSD.t968 VSUBS 0.024724f
C3277 VSSD.n623 VSUBS 0.022624f
C3278 VSSD.n624 VSUBS 0.011262f
C3279 VSSD.n625 VSUBS 0.03123f
C3280 VSSD.n626 VSUBS 0.03123f
C3281 VSSD.t49 VSUBS 0.023899f
C3282 VSSD.n627 VSUBS 0.037275f
C3283 VSSD.t51 VSUBS 0.027635f
C3284 VSSD.n628 VSUBS 0.021146f
C3285 VSSD.n629 VSUBS 0.03123f
C3286 VSSD.t283 VSUBS 0.010396f
C3287 VSSD.n630 VSUBS 0.018413f
C3288 VSSD.n631 VSUBS 0.021146f
C3289 VSSD.n632 VSUBS 0.03123f
C3290 VSSD.t909 VSUBS 0.013879f
C3291 VSSD.n633 VSUBS 0.018245f
C3292 VSSD.n634 VSUBS 0.021146f
C3293 VSSD.n635 VSUBS 0.03123f
C3294 VSSD.n636 VSUBS 0.015053f
C3295 VSSD.n637 VSUBS 0.03123f
C3296 VSSD.t619 VSUBS 0.024724f
C3297 VSSD.n639 VSUBS 0.022624f
C3298 VSSD.n640 VSUBS 0.011262f
C3299 VSSD.n641 VSUBS 0.03123f
C3300 VSSD.n642 VSUBS 0.03123f
C3301 VSSD.t1163 VSUBS 0.023899f
C3302 VSSD.n643 VSUBS 0.037275f
C3303 VSSD.t185 VSUBS 0.027635f
C3304 VSSD.n644 VSUBS 0.021146f
C3305 VSSD.n645 VSUBS 0.03123f
C3306 VSSD.t945 VSUBS 0.010396f
C3307 VSSD.n646 VSUBS 0.018413f
C3308 VSSD.n647 VSUBS 0.021146f
C3309 VSSD.n648 VSUBS 0.03123f
C3310 VSSD.t459 VSUBS 0.013879f
C3311 VSSD.n649 VSUBS 0.018245f
C3312 VSSD.n650 VSUBS 0.021146f
C3313 VSSD.n651 VSUBS 0.03123f
C3314 VSSD.n652 VSUBS 0.015053f
C3315 VSSD.n653 VSUBS 0.03123f
C3316 VSSD.t613 VSUBS 0.024724f
C3317 VSSD.n655 VSUBS 0.022624f
C3318 VSSD.n656 VSUBS 0.03123f
C3319 VSSD.n657 VSUBS 0.025373f
C3320 VSSD.n658 VSUBS 0.028587f
C3321 VSSD.n659 VSUBS 0.016086f
C3322 VSSD.n660 VSUBS 0.022892f
C3323 VSSD.n661 VSUBS 0.029102f
C3324 VSSD.n662 VSUBS 0.03123f
C3325 VSSD.n663 VSUBS 0.03123f
C3326 VSSD.n664 VSUBS 0.03123f
C3327 VSSD.n665 VSUBS 0.021146f
C3328 VSSD.n666 VSUBS 0.021146f
C3329 VSSD.n667 VSUBS 0.021146f
C3330 VSSD.n668 VSUBS 0.03123f
C3331 VSSD.n669 VSUBS 0.03123f
C3332 VSSD.n670 VSUBS 0.03123f
C3333 VSSD.n671 VSUBS 0.012984f
C3334 VSSD.n672 VSUBS 0.038003f
C3335 VSSD.n673 VSUBS 0.011146f
C3336 VSSD.n674 VSUBS 0.021146f
C3337 VSSD.n675 VSUBS 0.03123f
C3338 VSSD.n676 VSUBS 0.03123f
C3339 VSSD.n677 VSUBS 0.03123f
C3340 VSSD.n678 VSUBS 0.021146f
C3341 VSSD.n679 VSUBS 0.013561f
C3342 VSSD.n680 VSUBS 0.021657f
C3343 VSSD.n681 VSUBS 0.018158f
C3344 VSSD.n682 VSUBS 0.03123f
C3345 VSSD.n683 VSUBS 0.03123f
C3346 VSSD.n684 VSUBS 0.03123f
C3347 VSSD.n685 VSUBS 0.021146f
C3348 VSSD.n686 VSUBS 0.011033f
C3349 VSSD.n687 VSUBS 0.032298f
C3350 VSSD.n688 VSUBS 0.019996f
C3351 VSSD.n689 VSUBS 0.03123f
C3352 VSSD.n690 VSUBS 0.023423f
C3353 VSSD.n691 VSUBS 0.018501f
C3354 VSSD.n692 VSUBS 0.017122f
C3355 VSSD.n693 VSUBS 0.022892f
C3356 VSSD.n694 VSUBS 0.016086f
C3357 VSSD.n695 VSUBS 0.022892f
C3358 VSSD.n696 VSUBS 0.029102f
C3359 VSSD.n697 VSUBS 0.03123f
C3360 VSSD.n698 VSUBS 0.03123f
C3361 VSSD.n699 VSUBS 0.03123f
C3362 VSSD.n700 VSUBS 0.021146f
C3363 VSSD.n701 VSUBS 0.021146f
C3364 VSSD.n702 VSUBS 0.021146f
C3365 VSSD.n703 VSUBS 0.03123f
C3366 VSSD.n704 VSUBS 0.03123f
C3367 VSSD.n705 VSUBS 0.03123f
C3368 VSSD.n706 VSUBS 0.012984f
C3369 VSSD.n707 VSUBS 0.038003f
C3370 VSSD.n708 VSUBS 0.011146f
C3371 VSSD.n709 VSUBS 0.021146f
C3372 VSSD.n710 VSUBS 0.03123f
C3373 VSSD.n711 VSUBS 0.03123f
C3374 VSSD.n712 VSUBS 0.03123f
C3375 VSSD.n713 VSUBS 0.021146f
C3376 VSSD.n714 VSUBS 0.013561f
C3377 VSSD.n715 VSUBS 0.021657f
C3378 VSSD.n716 VSUBS 0.018158f
C3379 VSSD.n717 VSUBS 0.03123f
C3380 VSSD.n718 VSUBS 0.03123f
C3381 VSSD.n719 VSUBS 0.03123f
C3382 VSSD.n720 VSUBS 0.021146f
C3383 VSSD.n721 VSUBS 0.011033f
C3384 VSSD.n722 VSUBS 0.032298f
C3385 VSSD.n723 VSUBS 0.019996f
C3386 VSSD.n724 VSUBS 0.03123f
C3387 VSSD.n725 VSUBS 0.023423f
C3388 VSSD.n726 VSUBS 0.018501f
C3389 VSSD.n727 VSUBS 0.017122f
C3390 VSSD.n728 VSUBS 0.022892f
C3391 VSSD.n729 VSUBS 0.016086f
C3392 VSSD.n730 VSUBS 0.022892f
C3393 VSSD.n731 VSUBS 0.029102f
C3394 VSSD.n732 VSUBS 0.03123f
C3395 VSSD.n733 VSUBS 0.03123f
C3396 VSSD.n734 VSUBS 0.03123f
C3397 VSSD.n735 VSUBS 0.021146f
C3398 VSSD.n736 VSUBS 0.021146f
C3399 VSSD.n737 VSUBS 0.021146f
C3400 VSSD.n738 VSUBS 0.03123f
C3401 VSSD.n739 VSUBS 0.03123f
C3402 VSSD.n740 VSUBS 0.03123f
C3403 VSSD.n741 VSUBS 0.012984f
C3404 VSSD.n742 VSUBS 0.038003f
C3405 VSSD.n743 VSUBS 0.011146f
C3406 VSSD.n744 VSUBS 0.021146f
C3407 VSSD.n745 VSUBS 0.03123f
C3408 VSSD.n746 VSUBS 0.03123f
C3409 VSSD.n747 VSUBS 0.03123f
C3410 VSSD.n748 VSUBS 0.021146f
C3411 VSSD.n749 VSUBS 0.013561f
C3412 VSSD.n750 VSUBS 0.021657f
C3413 VSSD.n751 VSUBS 0.018158f
C3414 VSSD.n752 VSUBS 0.03123f
C3415 VSSD.n753 VSUBS 0.03123f
C3416 VSSD.n754 VSUBS 0.03123f
C3417 VSSD.n755 VSUBS 0.021146f
C3418 VSSD.n756 VSUBS 0.011033f
C3419 VSSD.n757 VSUBS 0.032298f
C3420 VSSD.n758 VSUBS 0.019996f
C3421 VSSD.n759 VSUBS 0.03123f
C3422 VSSD.n760 VSUBS 0.023423f
C3423 VSSD.n762 VSUBS -0.685653f
C3424 VSSD.n763 VSUBS 0.09704f
C3425 VSSD.t250 VSUBS 1.12632f
C3426 VSSD.t808 VSUBS 1.7682f
C3427 VSSD.t529 VSUBS 1.81059f
C3428 VSSD.t695 VSUBS 1.45331f
C3429 VSSD.t810 VSUBS 1.48359f
C3430 VSSD.t671 VSUBS 1.24137f
C3431 VSSD.t362 VSUBS 1.25954f
C3432 VSSD.t928 VSUBS 1.39881f
C3433 VSSD.t942 VSUBS 1.23532f
C3434 VSSD.t367 VSUBS 1.4412f
C3435 VSSD.t300 VSUBS 1.58653f
C3436 VSSD.t395 VSUBS 1.15659f
C3437 VSSD.t967 VSUBS 0.738764f
C3438 VSSD.n764 VSUBS 1.1908f
C3439 VSSD.t396 VSUBS 0.286292f
C3440 VSSD.t474 VSUBS 0.136721f
C3441 VSSD.t48 VSUBS 0.197283f
C3442 VSSD.t50 VSUBS 0.26794f
C3443 VSSD.t1132 VSUBS 0.274362f
C3444 VSSD.t282 VSUBS 0.220221f
C3445 VSSD.t46 VSUBS 0.224811f
C3446 VSSD.t669 VSUBS 0.188107f
C3447 VSSD.t708 VSUBS 0.190858f
C3448 VSSD.t908 VSUBS 0.211965f
C3449 VSSD.t186 VSUBS 0.187191f
C3450 VSSD.t672 VSUBS 0.21839f
C3451 VSSD.t707 VSUBS 0.240412f
C3452 VSSD.t670 VSUBS 0.17526f
C3453 VSSD.t618 VSUBS 0.305736f
C3454 VSSD.n765 VSUBS 1.72333f
C3455 VSSD.t506 VSUBS 0.690119f
C3456 VSSD.t616 VSUBS 0.955198f
C3457 VSSD.t119 VSUBS 0.726682f
C3458 VSSD.t121 VSUBS 0.767816f
C3459 VSSD.t792 VSUBS 0.767816f
C3460 VSSD.t174 VSUBS 0.991761f
C3461 VSSD.t162 VSUBS 0.639847f
C3462 VSSD.n766 VSUBS 0.272159f
C3463 VSSD.n767 VSUBS -0.10118f
C3464 VSSD.n768 VSUBS 0.010686f
C3465 VSSD.n769 VSUBS 0.03123f
C3466 VSSD.n770 VSUBS 0.018501f
C3467 VSSD.n771 VSUBS 0.01402f
C3468 VSSD.n772 VSUBS 0.011492f
C3469 VSSD.n773 VSUBS 0.023423f
C3470 VSSD.n774 VSUBS 0.03123f
C3471 VSSD.n775 VSUBS 0.020226f
C3472 VSSD.n776 VSUBS 0.031401f
C3473 VSSD.t120 VSUBS 0.021952f
C3474 VSSD.n777 VSUBS 0.029763f
C3475 VSSD.n778 VSUBS 0.020456f
C3476 VSSD.n779 VSUBS 0.03123f
C3477 VSSD.n780 VSUBS 0.018501f
C3478 VSSD.n781 VSUBS 0.023423f
C3479 VSSD.n782 VSUBS 0.011033f
C3480 VSSD.n783 VSUBS 0.036523f
C3481 VSSD.n784 VSUBS 0.020456f
C3482 VSSD.n785 VSUBS 0.04738f
C3483 VSSD.n786 VSUBS 0.018861f
C3484 VSSD.n787 VSUBS 2.34906f
C3485 VSSD.n788 VSUBS 2.02298f
C3486 VSSD.n789 VSUBS 1.52304f
C3487 VSSD.n790 VSUBS 1.96735f
C3488 VSSD.n791 VSUBS 0.03123f
C3489 VSSD.n792 VSUBS 0.01373f
C3490 VSSD.n793 VSUBS 0.01373f
C3491 VSSD.n794 VSUBS 0.01373f
C3492 VSSD.n795 VSUBS 0.03123f
C3493 VSSD.n796 VSUBS 0.01373f
C3494 VSSD.n797 VSUBS 0.01373f
C3495 VSSD.n798 VSUBS 0.01373f
C3496 VSSD.n799 VSUBS 0.05167f
C3497 VSSD.n800 VSUBS 0.03123f
C3498 VSSD.n801 VSUBS 0.01373f
C3499 VSSD.n802 VSUBS 0.01373f
C3500 VSSD.n803 VSUBS 0.01373f
C3501 VSSD.n804 VSUBS 0.01373f
C3502 VSSD.n805 VSUBS 0.0572f
C3503 VSSD.n806 VSUBS 0.03123f
C3504 VSSD.t721 VSUBS 0.02316f
C3505 VSSD.t352 VSUBS 0.02316f
C3506 VSSD.n808 VSUBS 0.03123f
C3507 VSSD.t366 VSUBS 0.024724f
C3508 VSSD.n811 VSUBS 0.03123f
C3509 VSSD.t568 VSUBS 0.024724f
C3510 VSSD.n812 VSUBS 0.011061f
C3511 VSSD.n813 VSUBS 0.03123f
C3512 VSSD.n815 VSUBS 0.03123f
C3513 VSSD.n816 VSUBS 0.011061f
C3514 VSSD.n817 VSUBS 0.03123f
C3515 VSSD.t1027 VSUBS 0.010396f
C3516 VSSD.n818 VSUBS 0.018748f
C3517 VSSD.t1098 VSUBS 0.010396f
C3518 VSSD.n819 VSUBS 0.018748f
C3519 VSSD.n821 VSUBS 0.03123f
C3520 VSSD.t964 VSUBS 0.028005f
C3521 VSSD.t33 VSUBS 0.028005f
C3522 VSSD.t154 VSUBS 0.024414f
C3523 VSSD.n822 VSUBS 0.023423f
C3524 VSSD.t27 VSUBS 0.024414f
C3525 VSSD.n825 VSUBS 0.048607f
C3526 VSSD.n826 VSUBS 0.03123f
C3527 VSSD.t896 VSUBS 0.024724f
C3528 VSSD.t626 VSUBS 0.024724f
C3529 VSSD.n827 VSUBS 0.011061f
C3530 VSSD.n828 VSUBS 0.03123f
C3531 VSSD.n830 VSUBS 0.03123f
C3532 VSSD.n831 VSUBS 0.011061f
C3533 VSSD.n832 VSUBS 0.03123f
C3534 VSSD.t1100 VSUBS 0.010396f
C3535 VSSD.n833 VSUBS 0.018748f
C3536 VSSD.t1079 VSUBS 0.010396f
C3537 VSSD.n834 VSUBS 0.018748f
C3538 VSSD.n836 VSUBS 0.03123f
C3539 VSSD.t348 VSUBS 0.028005f
C3540 VSSD.t289 VSUBS 0.028005f
C3541 VSSD.t685 VSUBS 0.024414f
C3542 VSSD.n837 VSUBS 0.023423f
C3543 VSSD.t873 VSUBS 0.024414f
C3544 VSSD.n840 VSUBS 0.048607f
C3545 VSSD.n841 VSUBS 0.03123f
C3546 VSSD.t537 VSUBS 0.024724f
C3547 VSSD.t812 VSUBS 0.024724f
C3548 VSSD.n842 VSUBS 0.011061f
C3549 VSSD.n843 VSUBS 0.03123f
C3550 VSSD.n845 VSUBS 0.03123f
C3551 VSSD.n846 VSUBS 0.011061f
C3552 VSSD.n847 VSUBS 0.03123f
C3553 VSSD.t1066 VSUBS 0.010396f
C3554 VSSD.n848 VSUBS 0.018748f
C3555 VSSD.t1025 VSUBS 0.010396f
C3556 VSSD.n849 VSUBS 0.018748f
C3557 VSSD.n851 VSUBS 0.03123f
C3558 VSSD.t503 VSUBS 0.028005f
C3559 VSSD.t686 VSUBS 0.028005f
C3560 VSSD.t1113 VSUBS 0.024414f
C3561 VSSD.n852 VSUBS 0.023423f
C3562 VSSD.t76 VSUBS 0.024414f
C3563 VSSD.n855 VSUBS 0.048607f
C3564 VSSD.n856 VSUBS 0.03123f
C3565 VSSD.t31 VSUBS 0.024724f
C3566 VSSD.t813 VSUBS 0.024724f
C3567 VSSD.n857 VSUBS 0.011061f
C3568 VSSD.n858 VSUBS 0.03123f
C3569 VSSD.n860 VSUBS 0.03123f
C3570 VSSD.n861 VSUBS 0.011061f
C3571 VSSD.n862 VSUBS 0.03123f
C3572 VSSD.t1073 VSUBS 0.010396f
C3573 VSSD.n863 VSUBS 0.018748f
C3574 VSSD.t1036 VSUBS 0.010396f
C3575 VSSD.n864 VSUBS 0.018748f
C3576 VSSD.n866 VSUBS 0.03123f
C3577 VSSD.t88 VSUBS 0.028005f
C3578 VSSD.t129 VSUBS 0.028005f
C3579 VSSD.t90 VSUBS 0.024414f
C3580 VSSD.n867 VSUBS 0.023423f
C3581 VSSD.t130 VSUBS 0.024414f
C3582 VSSD.n870 VSUBS 0.048607f
C3583 VSSD.n871 VSUBS 0.03123f
C3584 VSSD.t364 VSUBS 0.024724f
C3585 VSSD.t885 VSUBS 0.024724f
C3586 VSSD.n872 VSUBS 0.011061f
C3587 VSSD.n873 VSUBS 0.03123f
C3588 VSSD.n875 VSUBS 0.03123f
C3589 VSSD.n876 VSUBS 0.011061f
C3590 VSSD.n877 VSUBS 0.03123f
C3591 VSSD.t1055 VSUBS 0.010396f
C3592 VSSD.n878 VSUBS 0.018748f
C3593 VSSD.t1007 VSUBS 0.010396f
C3594 VSSD.n879 VSUBS 0.018748f
C3595 VSSD.n881 VSUBS 0.03123f
C3596 VSSD.t736 VSUBS 0.028005f
C3597 VSSD.t140 VSUBS 0.028005f
C3598 VSSD.t198 VSUBS 0.024414f
C3599 VSSD.n882 VSUBS 0.023423f
C3600 VSSD.t169 VSUBS 0.024414f
C3601 VSSD.n885 VSUBS 0.048607f
C3602 VSSD.n886 VSUBS 0.03123f
C3603 VSSD.t900 VSUBS 0.024724f
C3604 VSSD.t937 VSUBS 0.024724f
C3605 VSSD.n887 VSUBS 0.011061f
C3606 VSSD.n888 VSUBS 0.03123f
C3607 VSSD.n890 VSUBS 0.03123f
C3608 VSSD.n891 VSUBS 0.011061f
C3609 VSSD.n892 VSUBS 0.03123f
C3610 VSSD.t1090 VSUBS 0.010396f
C3611 VSSD.n893 VSUBS 0.018748f
C3612 VSSD.t1062 VSUBS 0.010396f
C3613 VSSD.n894 VSUBS 0.018748f
C3614 VSSD.n896 VSUBS 0.03123f
C3615 VSSD.t586 VSUBS 0.028005f
C3616 VSSD.t958 VSUBS 0.028005f
C3617 VSSD.t1179 VSUBS 0.024414f
C3618 VSSD.n897 VSUBS 0.023423f
C3619 VSSD.t960 VSUBS 0.024414f
C3620 VSSD.n900 VSUBS 0.048607f
C3621 VSSD.n901 VSUBS 0.03123f
C3622 VSSD.t98 VSUBS 0.024724f
C3623 VSSD.t569 VSUBS 0.024724f
C3624 VSSD.n902 VSUBS 0.011061f
C3625 VSSD.n903 VSUBS 0.03123f
C3626 VSSD.n905 VSUBS 0.03123f
C3627 VSSD.n906 VSUBS 0.011061f
C3628 VSSD.n907 VSUBS 0.03123f
C3629 VSSD.t1085 VSUBS 0.010396f
C3630 VSSD.n908 VSUBS 0.018748f
C3631 VSSD.t1059 VSUBS 0.010396f
C3632 VSSD.n909 VSUBS 0.018748f
C3633 VSSD.n911 VSUBS 0.03123f
C3634 VSSD.t42 VSUBS 0.028005f
C3635 VSSD.t620 VSUBS 0.028005f
C3636 VSSD.t1148 VSUBS 0.024414f
C3637 VSSD.n912 VSUBS 0.023423f
C3638 VSSD.t80 VSUBS 0.024414f
C3639 VSSD.n915 VSUBS 0.048607f
C3640 VSSD.n916 VSUBS 0.03123f
C3641 VSSD.t1192 VSUBS 0.024724f
C3642 VSSD.t571 VSUBS 0.024724f
C3643 VSSD.n917 VSUBS 0.011061f
C3644 VSSD.n918 VSUBS 0.03123f
C3645 VSSD.n920 VSUBS 0.03123f
C3646 VSSD.n921 VSUBS 0.011061f
C3647 VSSD.n922 VSUBS 0.03123f
C3648 VSSD.t1040 VSUBS 0.010396f
C3649 VSSD.n923 VSUBS 0.018748f
C3650 VSSD.t1103 VSUBS 0.010396f
C3651 VSSD.n924 VSUBS 0.018748f
C3652 VSSD.n926 VSUBS 0.03123f
C3653 VSSD.t565 VSUBS 0.028005f
C3654 VSSD.t755 VSUBS 0.028005f
C3655 VSSD.t603 VSUBS 0.024414f
C3656 VSSD.n927 VSUBS 0.023423f
C3657 VSSD.t754 VSUBS 0.024414f
C3658 VSSD.n930 VSUBS 0.048607f
C3659 VSSD.n931 VSUBS 0.03123f
C3660 VSSD.t228 VSUBS 0.024724f
C3661 VSSD.t884 VSUBS 0.024724f
C3662 VSSD.n932 VSUBS 0.011061f
C3663 VSSD.n933 VSUBS 0.03123f
C3664 VSSD.n935 VSUBS 0.03123f
C3665 VSSD.n936 VSUBS 0.011061f
C3666 VSSD.n937 VSUBS 0.03123f
C3667 VSSD.t1013 VSUBS 0.010396f
C3668 VSSD.n938 VSUBS 0.018748f
C3669 VSSD.t1034 VSUBS 0.010396f
C3670 VSSD.n939 VSUBS 0.018748f
C3671 VSSD.n941 VSUBS 0.03123f
C3672 VSSD.t734 VSUBS 0.028005f
C3673 VSSD.t1150 VSUBS 0.028005f
C3674 VSSD.t918 VSUBS 0.024414f
C3675 VSSD.n942 VSUBS 0.023423f
C3676 VSSD.t1151 VSUBS 0.024414f
C3677 VSSD.n945 VSUBS 0.048607f
C3678 VSSD.n946 VSUBS 0.03123f
C3679 VSSD.t898 VSUBS 0.024724f
C3680 VSSD.t936 VSUBS 0.024724f
C3681 VSSD.n947 VSUBS 0.011061f
C3682 VSSD.n948 VSUBS 0.03123f
C3683 VSSD.n950 VSUBS 0.03123f
C3684 VSSD.n951 VSUBS 0.011061f
C3685 VSSD.n952 VSUBS 0.03123f
C3686 VSSD.t1065 VSUBS 0.010396f
C3687 VSSD.n953 VSUBS 0.018748f
C3688 VSSD.t1019 VSUBS 0.010396f
C3689 VSSD.n954 VSUBS 0.018748f
C3690 VSSD.t1140 VSUBS 0.024414f
C3691 VSSD.t107 VSUBS 0.024414f
C3692 VSSD.n956 VSUBS 0.06129f
C3693 VSSD.t1141 VSUBS 0.028005f
C3694 VSSD.t799 VSUBS 0.028005f
C3695 VSSD.n957 VSUBS 0.058811f
C3696 VSSD.n958 VSUBS 0.023247f
C3697 VSSD.n959 VSUBS 0.104916f
C3698 VSSD.n960 VSUBS 0.03123f
C3699 VSSD.n961 VSUBS 0.011061f
C3700 VSSD.n963 VSUBS 0.029315f
C3701 VSSD.n965 VSUBS 0.03123f
C3702 VSSD.n966 VSUBS 0.03123f
C3703 VSSD.n967 VSUBS 0.03123f
C3704 VSSD.n968 VSUBS 0.011061f
C3705 VSSD.n969 VSUBS 0.011061f
C3706 VSSD.t962 VSUBS 0.013879f
C3707 VSSD.n970 VSUBS 0.017846f
C3708 VSSD.t345 VSUBS 0.013879f
C3709 VSSD.n971 VSUBS 0.017846f
C3710 VSSD.n972 VSUBS 0.049994f
C3711 VSSD.n974 VSUBS 0.03123f
C3712 VSSD.n975 VSUBS 0.03123f
C3713 VSSD.n976 VSUBS 0.03123f
C3714 VSSD.n977 VSUBS 0.011061f
C3715 VSSD.n978 VSUBS 0.011061f
C3716 VSSD.n979 VSUBS 0.011061f
C3717 VSSD.n980 VSUBS 0.03123f
C3718 VSSD.n981 VSUBS 0.03123f
C3719 VSSD.n982 VSUBS 0.03123f
C3720 VSSD.n984 VSUBS 0.061563f
C3721 VSSD.n986 VSUBS 0.03123f
C3722 VSSD.n987 VSUBS 0.03123f
C3723 VSSD.n988 VSUBS 0.018501f
C3724 VSSD.n990 VSUBS 0.06644f
C3725 VSSD.n992 VSUBS 0.057443f
C3726 VSSD.n993 VSUBS 0.03123f
C3727 VSSD.n994 VSUBS 0.03123f
C3728 VSSD.n995 VSUBS 0.03123f
C3729 VSSD.n996 VSUBS 0.011061f
C3730 VSSD.n998 VSUBS 0.029315f
C3731 VSSD.n1000 VSUBS 0.03123f
C3732 VSSD.n1001 VSUBS 0.03123f
C3733 VSSD.n1002 VSUBS 0.03123f
C3734 VSSD.n1003 VSUBS 0.011061f
C3735 VSSD.n1004 VSUBS 0.011061f
C3736 VSSD.t841 VSUBS 0.013879f
C3737 VSSD.n1005 VSUBS 0.017846f
C3738 VSSD.t941 VSUBS 0.013879f
C3739 VSSD.n1006 VSUBS 0.017846f
C3740 VSSD.n1007 VSUBS 0.049994f
C3741 VSSD.n1009 VSUBS 0.03123f
C3742 VSSD.n1010 VSUBS 0.03123f
C3743 VSSD.n1011 VSUBS 0.03123f
C3744 VSSD.n1012 VSUBS 0.011061f
C3745 VSSD.n1013 VSUBS 0.011061f
C3746 VSSD.n1014 VSUBS 0.011061f
C3747 VSSD.n1015 VSUBS 0.03123f
C3748 VSSD.n1016 VSUBS 0.03123f
C3749 VSSD.n1017 VSUBS 0.03123f
C3750 VSSD.n1019 VSUBS 0.061563f
C3751 VSSD.n1021 VSUBS 0.03123f
C3752 VSSD.n1022 VSUBS 0.03123f
C3753 VSSD.n1023 VSUBS 0.018501f
C3754 VSSD.n1025 VSUBS 0.06644f
C3755 VSSD.n1027 VSUBS 0.057443f
C3756 VSSD.n1028 VSUBS 0.03123f
C3757 VSSD.n1029 VSUBS 0.03123f
C3758 VSSD.n1030 VSUBS 0.03123f
C3759 VSSD.n1031 VSUBS 0.011061f
C3760 VSSD.n1033 VSUBS 0.029315f
C3761 VSSD.n1035 VSUBS 0.03123f
C3762 VSSD.n1036 VSUBS 0.03123f
C3763 VSSD.n1037 VSUBS 0.03123f
C3764 VSSD.n1038 VSUBS 0.011061f
C3765 VSSD.n1039 VSUBS 0.011061f
C3766 VSSD.t957 VSUBS 0.013879f
C3767 VSSD.n1040 VSUBS 0.017846f
C3768 VSSD.t679 VSUBS 0.013879f
C3769 VSSD.n1041 VSUBS 0.017846f
C3770 VSSD.n1042 VSUBS 0.049994f
C3771 VSSD.n1044 VSUBS 0.03123f
C3772 VSSD.n1045 VSUBS 0.03123f
C3773 VSSD.n1046 VSUBS 0.03123f
C3774 VSSD.n1047 VSUBS 0.011061f
C3775 VSSD.n1048 VSUBS 0.011061f
C3776 VSSD.n1049 VSUBS 0.011061f
C3777 VSSD.n1050 VSUBS 0.03123f
C3778 VSSD.n1051 VSUBS 0.03123f
C3779 VSSD.n1052 VSUBS 0.03123f
C3780 VSSD.n1054 VSUBS 0.061563f
C3781 VSSD.n1056 VSUBS 0.03123f
C3782 VSSD.n1057 VSUBS 0.03123f
C3783 VSSD.n1058 VSUBS 0.018501f
C3784 VSSD.n1060 VSUBS 0.06644f
C3785 VSSD.n1062 VSUBS 0.057443f
C3786 VSSD.n1063 VSUBS 0.03123f
C3787 VSSD.n1064 VSUBS 0.03123f
C3788 VSSD.n1065 VSUBS 0.03123f
C3789 VSSD.n1066 VSUBS 0.011061f
C3790 VSSD.n1068 VSUBS 0.029315f
C3791 VSSD.n1070 VSUBS 0.03123f
C3792 VSSD.n1071 VSUBS 0.03123f
C3793 VSSD.n1072 VSUBS 0.03123f
C3794 VSSD.n1073 VSUBS 0.011061f
C3795 VSSD.n1074 VSUBS 0.011061f
C3796 VSSD.t607 VSUBS 0.013879f
C3797 VSSD.n1075 VSUBS 0.017846f
C3798 VSSD.t179 VSUBS 0.013879f
C3799 VSSD.n1076 VSUBS 0.017846f
C3800 VSSD.n1077 VSUBS 0.049994f
C3801 VSSD.n1079 VSUBS 0.03123f
C3802 VSSD.n1080 VSUBS 0.03123f
C3803 VSSD.n1081 VSUBS 0.03123f
C3804 VSSD.n1082 VSUBS 0.011061f
C3805 VSSD.n1083 VSUBS 0.011061f
C3806 VSSD.n1084 VSUBS 0.011061f
C3807 VSSD.n1085 VSUBS 0.03123f
C3808 VSSD.n1086 VSUBS 0.03123f
C3809 VSSD.n1087 VSUBS 0.03123f
C3810 VSSD.n1089 VSUBS 0.061563f
C3811 VSSD.n1091 VSUBS 0.03123f
C3812 VSSD.n1092 VSUBS 0.03123f
C3813 VSSD.n1093 VSUBS 0.018501f
C3814 VSSD.n1095 VSUBS 0.06644f
C3815 VSSD.n1097 VSUBS 0.057443f
C3816 VSSD.n1098 VSUBS 0.03123f
C3817 VSSD.n1099 VSUBS 0.03123f
C3818 VSSD.n1100 VSUBS 0.03123f
C3819 VSSD.n1101 VSUBS 0.011061f
C3820 VSSD.n1103 VSUBS 0.029315f
C3821 VSSD.n1105 VSUBS 0.03123f
C3822 VSSD.n1106 VSUBS 0.03123f
C3823 VSSD.n1107 VSUBS 0.03123f
C3824 VSSD.n1108 VSUBS 0.011061f
C3825 VSSD.n1109 VSUBS 0.011061f
C3826 VSSD.t828 VSUBS 0.013879f
C3827 VSSD.n1110 VSUBS 0.017846f
C3828 VSSD.t494 VSUBS 0.013879f
C3829 VSSD.n1111 VSUBS 0.017846f
C3830 VSSD.n1112 VSUBS 0.049994f
C3831 VSSD.n1114 VSUBS 0.03123f
C3832 VSSD.n1115 VSUBS 0.03123f
C3833 VSSD.n1116 VSUBS 0.03123f
C3834 VSSD.n1117 VSUBS 0.011061f
C3835 VSSD.n1118 VSUBS 0.011061f
C3836 VSSD.n1119 VSUBS 0.011061f
C3837 VSSD.n1120 VSUBS 0.03123f
C3838 VSSD.n1121 VSUBS 0.03123f
C3839 VSSD.n1122 VSUBS 0.03123f
C3840 VSSD.n1124 VSUBS 0.061563f
C3841 VSSD.n1126 VSUBS 0.03123f
C3842 VSSD.n1127 VSUBS 0.03123f
C3843 VSSD.n1128 VSUBS 0.018501f
C3844 VSSD.n1130 VSUBS 0.06644f
C3845 VSSD.n1132 VSUBS 0.057443f
C3846 VSSD.n1133 VSUBS 0.03123f
C3847 VSSD.n1134 VSUBS 0.03123f
C3848 VSSD.n1135 VSUBS 0.03123f
C3849 VSSD.n1136 VSUBS 0.011061f
C3850 VSSD.n1138 VSUBS 0.029315f
C3851 VSSD.n1140 VSUBS 0.03123f
C3852 VSSD.n1141 VSUBS 0.03123f
C3853 VSSD.n1142 VSUBS 0.03123f
C3854 VSSD.n1143 VSUBS 0.011061f
C3855 VSSD.n1144 VSUBS 0.011061f
C3856 VSSD.t389 VSUBS 0.013879f
C3857 VSSD.n1145 VSUBS 0.017846f
C3858 VSSD.t489 VSUBS 0.013879f
C3859 VSSD.n1146 VSUBS 0.017846f
C3860 VSSD.n1147 VSUBS 0.049994f
C3861 VSSD.n1149 VSUBS 0.03123f
C3862 VSSD.n1150 VSUBS 0.03123f
C3863 VSSD.n1151 VSUBS 0.03123f
C3864 VSSD.n1152 VSUBS 0.011061f
C3865 VSSD.n1153 VSUBS 0.011061f
C3866 VSSD.n1154 VSUBS 0.011061f
C3867 VSSD.n1155 VSUBS 0.03123f
C3868 VSSD.n1156 VSUBS 0.03123f
C3869 VSSD.n1157 VSUBS 0.03123f
C3870 VSSD.n1159 VSUBS 0.061563f
C3871 VSSD.n1161 VSUBS 0.03123f
C3872 VSSD.n1162 VSUBS 0.03123f
C3873 VSSD.n1163 VSUBS 0.018501f
C3874 VSSD.n1165 VSUBS 0.06644f
C3875 VSSD.n1167 VSUBS 0.057443f
C3876 VSSD.n1168 VSUBS 0.03123f
C3877 VSSD.n1169 VSUBS 0.03123f
C3878 VSSD.n1170 VSUBS 0.03123f
C3879 VSSD.n1171 VSUBS 0.011061f
C3880 VSSD.n1173 VSUBS 0.029315f
C3881 VSSD.n1175 VSUBS 0.03123f
C3882 VSSD.n1176 VSUBS 0.03123f
C3883 VSSD.n1177 VSUBS 0.03123f
C3884 VSSD.n1178 VSUBS 0.011061f
C3885 VSSD.n1179 VSUBS 0.011061f
C3886 VSSD.t63 VSUBS 0.013879f
C3887 VSSD.n1180 VSUBS 0.017846f
C3888 VSSD.t35 VSUBS 0.013879f
C3889 VSSD.n1181 VSUBS 0.017846f
C3890 VSSD.n1182 VSUBS 0.049994f
C3891 VSSD.n1184 VSUBS 0.03123f
C3892 VSSD.n1185 VSUBS 0.03123f
C3893 VSSD.n1186 VSUBS 0.03123f
C3894 VSSD.n1187 VSUBS 0.011061f
C3895 VSSD.n1188 VSUBS 0.011061f
C3896 VSSD.n1189 VSUBS 0.011061f
C3897 VSSD.n1190 VSUBS 0.03123f
C3898 VSSD.n1191 VSUBS 0.03123f
C3899 VSSD.n1192 VSUBS 0.03123f
C3900 VSSD.n1194 VSUBS 0.061563f
C3901 VSSD.n1196 VSUBS 0.03123f
C3902 VSSD.n1197 VSUBS 0.03123f
C3903 VSSD.n1198 VSUBS 0.018501f
C3904 VSSD.n1200 VSUBS 0.06644f
C3905 VSSD.n1202 VSUBS 0.057443f
C3906 VSSD.n1203 VSUBS 0.03123f
C3907 VSSD.n1204 VSUBS 0.03123f
C3908 VSSD.n1205 VSUBS 0.03123f
C3909 VSSD.n1206 VSUBS 0.011061f
C3910 VSSD.n1208 VSUBS 0.029315f
C3911 VSSD.n1210 VSUBS 0.03123f
C3912 VSSD.n1211 VSUBS 0.03123f
C3913 VSSD.n1212 VSUBS 0.03123f
C3914 VSSD.n1213 VSUBS 0.011061f
C3915 VSSD.n1214 VSUBS 0.011061f
C3916 VSSD.t836 VSUBS 0.013879f
C3917 VSSD.n1215 VSUBS 0.017846f
C3918 VSSD.t835 VSUBS 0.013879f
C3919 VSSD.n1216 VSUBS 0.017846f
C3920 VSSD.n1217 VSUBS 0.049994f
C3921 VSSD.n1219 VSUBS 0.03123f
C3922 VSSD.n1220 VSUBS 0.03123f
C3923 VSSD.n1221 VSUBS 0.03123f
C3924 VSSD.n1222 VSUBS 0.011061f
C3925 VSSD.n1223 VSUBS 0.011061f
C3926 VSSD.n1224 VSUBS 0.011061f
C3927 VSSD.n1225 VSUBS 0.03123f
C3928 VSSD.n1226 VSUBS 0.03123f
C3929 VSSD.n1227 VSUBS 0.03123f
C3930 VSSD.n1229 VSUBS 0.061563f
C3931 VSSD.n1231 VSUBS 0.03123f
C3932 VSSD.n1232 VSUBS 0.03123f
C3933 VSSD.n1233 VSUBS 0.018501f
C3934 VSSD.n1235 VSUBS 0.06644f
C3935 VSSD.n1237 VSUBS 0.057443f
C3936 VSSD.n1238 VSUBS 0.03123f
C3937 VSSD.n1239 VSUBS 0.03123f
C3938 VSSD.n1240 VSUBS 0.03123f
C3939 VSSD.n1241 VSUBS 0.011061f
C3940 VSSD.n1243 VSUBS 0.029315f
C3941 VSSD.n1245 VSUBS 0.03123f
C3942 VSSD.n1246 VSUBS 0.03123f
C3943 VSSD.n1247 VSUBS 0.03123f
C3944 VSSD.n1248 VSUBS 0.011061f
C3945 VSSD.n1249 VSUBS 0.011061f
C3946 VSSD.t405 VSUBS 0.013879f
C3947 VSSD.n1250 VSUBS 0.017846f
C3948 VSSD.t984 VSUBS 0.013879f
C3949 VSSD.n1251 VSUBS 0.017846f
C3950 VSSD.n1252 VSUBS 0.049994f
C3951 VSSD.n1254 VSUBS 0.03123f
C3952 VSSD.n1255 VSUBS 0.03123f
C3953 VSSD.n1256 VSUBS 0.03123f
C3954 VSSD.n1257 VSUBS 0.011061f
C3955 VSSD.n1258 VSUBS 0.011061f
C3956 VSSD.n1259 VSUBS 0.011061f
C3957 VSSD.n1260 VSUBS 0.03123f
C3958 VSSD.n1261 VSUBS 0.03123f
C3959 VSSD.n1262 VSUBS 0.03123f
C3960 VSSD.n1264 VSUBS 0.061563f
C3961 VSSD.n1266 VSUBS 0.03123f
C3962 VSSD.n1267 VSUBS 0.03123f
C3963 VSSD.n1268 VSUBS 0.018501f
C3964 VSSD.n1270 VSUBS 0.06644f
C3965 VSSD.n1272 VSUBS 0.057443f
C3966 VSSD.n1273 VSUBS 0.03123f
C3967 VSSD.n1274 VSUBS 0.03123f
C3968 VSSD.n1275 VSUBS 0.03123f
C3969 VSSD.n1276 VSUBS 0.011061f
C3970 VSSD.n1278 VSUBS 0.029315f
C3971 VSSD.n1280 VSUBS 0.03123f
C3972 VSSD.n1281 VSUBS 0.03123f
C3973 VSSD.n1282 VSUBS 0.03123f
C3974 VSSD.n1283 VSUBS 0.011061f
C3975 VSSD.n1284 VSUBS 0.011061f
C3976 VSSD.t336 VSUBS 0.013879f
C3977 VSSD.n1285 VSUBS 0.017846f
C3978 VSSD.t86 VSUBS 0.013879f
C3979 VSSD.n1286 VSUBS 0.017846f
C3980 VSSD.n1287 VSUBS 0.049994f
C3981 VSSD.n1289 VSUBS 0.03123f
C3982 VSSD.n1290 VSUBS 0.03123f
C3983 VSSD.n1291 VSUBS 0.03123f
C3984 VSSD.n1292 VSUBS 0.011061f
C3985 VSSD.n1293 VSUBS 0.011061f
C3986 VSSD.n1294 VSUBS 0.011061f
C3987 VSSD.n1295 VSUBS 0.03123f
C3988 VSSD.n1296 VSUBS 0.03123f
C3989 VSSD.n1297 VSUBS 0.03123f
C3990 VSSD.n1299 VSUBS 0.061563f
C3991 VSSD.n1301 VSUBS 0.048607f
C3992 VSSD.n1302 VSUBS 0.03123f
C3993 VSSD.n1303 VSUBS 0.018501f
C3994 VSSD.n1304 VSUBS 0.023423f
C3995 VSSD.n1306 VSUBS 0.091197f
C3996 VSSD.n1308 VSUBS 0.03123f
C3997 VSSD.n1309 VSUBS 0.03123f
C3998 VSSD.n1310 VSUBS 0.03123f
C3999 VSSD.n1312 VSUBS 0.05167f
C4000 VSSD.n1315 VSUBS 0.03123f
C4001 VSSD.n1316 VSUBS 0.03123f
C4002 VSSD.n1318 VSUBS 0.0572f
C4003 VSSD.n1320 VSUBS 0.0572f
C4004 VSSD.n1321 VSUBS 0.03123f
C4005 VSSD.n1322 VSUBS 0.016464f
C4006 VSSD.n1323 VSUBS 0.2361f
C4007 VSSD.n1324 VSUBS 2.54819f
C4008 VSSD.n1325 VSUBS 2.55828f
C4009 VSSD.n1326 VSUBS 0.03123f
C4010 VSSD.t636 VSUBS 0.028005f
C4011 VSSD.n1328 VSUBS 0.03123f
C4012 VSSD.n1329 VSUBS 0.011061f
C4013 VSSD.n1330 VSUBS 0.03123f
C4014 VSSD.t611 VSUBS 0.013879f
C4015 VSSD.n1331 VSUBS 0.017846f
C4016 VSSD.n1332 VSUBS 0.029746f
C4017 VSSD.n1333 VSUBS 0.03123f
C4018 VSSD.n1334 VSUBS 0.011061f
C4019 VSSD.n1335 VSUBS 0.03123f
C4020 VSSD.t976 VSUBS 0.024724f
C4021 VSSD.t714 VSUBS 0.024414f
C4022 VSSD.n1337 VSUBS 0.040253f
C4023 VSSD.n1338 VSUBS 0.03123f
C4024 VSSD.n1339 VSUBS 0.011061f
C4025 VSSD.n1340 VSUBS 0.03123f
C4026 VSSD.n1341 VSUBS 0.011061f
C4027 VSSD.n1342 VSUBS 0.03123f
C4028 VSSD.n1343 VSUBS 0.011061f
C4029 VSSD.n1344 VSUBS 0.03123f
C4030 VSSD.n1346 VSUBS 0.03123f
C4031 VSSD.n1349 VSUBS 0.03123f
C4032 VSSD.t664 VSUBS 0.028005f
C4033 VSSD.n1351 VSUBS 0.03123f
C4034 VSSD.n1352 VSUBS 0.011061f
C4035 VSSD.n1353 VSUBS 0.03123f
C4036 VSSD.t606 VSUBS 0.013879f
C4037 VSSD.n1354 VSUBS 0.017846f
C4038 VSSD.n1355 VSUBS 0.029746f
C4039 VSSD.n1356 VSUBS 0.03123f
C4040 VSSD.n1357 VSUBS 0.011061f
C4041 VSSD.n1358 VSUBS 0.03123f
C4042 VSSD.t105 VSUBS 0.024724f
C4043 VSSD.t903 VSUBS 0.024414f
C4044 VSSD.n1360 VSUBS 0.040253f
C4045 VSSD.n1361 VSUBS 0.03123f
C4046 VSSD.n1362 VSUBS 0.011061f
C4047 VSSD.n1363 VSUBS 0.03123f
C4048 VSSD.n1364 VSUBS 0.011061f
C4049 VSSD.n1365 VSUBS 0.03123f
C4050 VSSD.n1366 VSUBS 0.011061f
C4051 VSSD.n1367 VSUBS 0.03123f
C4052 VSSD.n1369 VSUBS 0.03123f
C4053 VSSD.n1372 VSUBS 0.03123f
C4054 VSSD.t144 VSUBS 0.028005f
C4055 VSSD.n1374 VSUBS 0.03123f
C4056 VSSD.n1375 VSUBS 0.011061f
C4057 VSSD.n1376 VSUBS 0.03123f
C4058 VSSD.t241 VSUBS 0.013879f
C4059 VSSD.n1377 VSUBS 0.017846f
C4060 VSSD.n1378 VSUBS 0.029746f
C4061 VSSD.n1379 VSUBS 0.03123f
C4062 VSSD.n1380 VSUBS 0.011061f
C4063 VSSD.n1381 VSUBS 0.03123f
C4064 VSSD.t983 VSUBS 0.024724f
C4065 VSSD.n1383 VSUBS 0.011001f
C4066 VSSD.n1384 VSUBS 0.03123f
C4067 VSSD.t635 VSUBS 1.82705f
C4068 VSSD.t628 VSUBS 1.87085f
C4069 VSSD.t274 VSUBS 1.50168f
C4070 VSSD.t637 VSUBS 1.53297f
C4071 VSSD.t993 VSUBS 1.28269f
C4072 VSSD.t745 VSUBS 1.30146f
C4073 VSSD.t610 VSUBS 1.44537f
C4074 VSSD.t728 VSUBS 1.27643f
C4075 VSSD.t783 VSUBS 1.48917f
C4076 VSSD.t746 VSUBS 1.63934f
C4077 VSSD.t994 VSUBS 1.19509f
C4078 VSSD.t975 VSUBS 2.18996f
C4079 VSSD.t933 VSUBS 2.12113f
C4080 VSSD.t204 VSUBS 0.719557f
C4081 VSSD.t713 VSUBS 1.558f
C4082 VSSD.t252 VSUBS 1.82705f
C4083 VSSD.t940 VSUBS 1.87085f
C4084 VSSD.t1126 VSUBS 1.50168f
C4085 VSSD.t715 VSUBS 1.53297f
C4086 VSSD.t919 VSUBS 1.28269f
C4087 VSSD.t1178 VSUBS 1.30146f
C4088 VSSD.t1144 VSUBS 1.44537f
C4089 VSSD.t726 VSUBS 1.27643f
C4090 VSSD.t52 VSUBS 1.48917f
C4091 VSSD.t842 VSUBS 1.63934f
C4092 VSSD.t922 VSUBS 1.19509f
C4093 VSSD.t1152 VSUBS 2.18996f
C4094 VSSD.t920 VSUBS 2.12113f
C4095 VSSD.t1155 VSUBS 0.719557f
C4096 VSSD.t661 VSUBS 1.558f
C4097 VSSD.t663 VSUBS 1.82705f
C4098 VSSD.t593 VSUBS 1.87085f
C4099 VSSD.t998 VSUBS 1.50168f
C4100 VSSD.t131 VSUBS 1.53297f
C4101 VSSD.t394 VSUBS 1.28269f
C4102 VSSD.t784 VSUBS 1.30146f
C4103 VSSD.t605 VSUBS 1.44537f
C4104 VSSD.t511 VSUBS 1.27643f
C4105 VSSD.t703 VSUBS 1.48917f
C4106 VSSD.t704 VSUBS 1.63934f
C4107 VSSD.t1142 VSUBS 1.19509f
C4108 VSSD.t104 VSUBS 2.18996f
C4109 VSSD.t453 VSUBS 2.12113f
C4110 VSSD.t71 VSUBS 0.719557f
C4111 VSSD.t902 VSUBS 1.558f
C4112 VSSD.t906 VSUBS 1.82705f
C4113 VSSD.t214 VSUBS 1.87085f
C4114 VSSD.t13 VSUBS 1.50168f
C4115 VSSD.t904 VSUBS 1.53297f
C4116 VSSD.t609 VSUBS 1.28269f
C4117 VSSD.t939 VSUBS 1.30146f
C4118 VSSD.t485 VSUBS 1.44537f
C4119 VSSD.t266 VSUBS 1.27643f
C4120 VSSD.t767 VSUBS 1.48917f
C4121 VSSD.t938 VSUBS 1.63934f
C4122 VSSD.t608 VSUBS 1.19509f
C4123 VSSD.t652 VSUBS 2.18996f
C4124 VSSD.t765 VSUBS 2.12113f
C4125 VSSD.t208 VSUBS 0.719557f
C4126 VSSD.t145 VSUBS 1.558f
C4127 VSSD.t143 VSUBS 1.82705f
C4128 VSSD.t155 VSUBS 1.87085f
C4129 VSSD.t623 VSUBS 1.50168f
C4130 VSSD.t147 VSUBS 1.53297f
C4131 VSSD.t423 VSUBS 1.28269f
C4132 VSSD.t141 VSUBS 1.30146f
C4133 VSSD.t240 VSUBS 1.44537f
C4134 VSSD.t270 VSUBS 1.27643f
C4135 VSSD.t43 VSUBS 1.48917f
C4136 VSSD.t699 VSUBS 1.63934f
C4137 VSSD.t422 VSUBS 1.19509f
C4138 VSSD.t982 VSUBS 2.18996f
C4139 VSSD.t420 VSUBS 2.12113f
C4140 VSSD.t73 VSUBS 0.719557f
C4141 VSSD.t455 VSUBS 1.92716f
C4142 VSSD.t1028 VSUBS 1.20135f
C4143 VSSD.t759 VSUBS 0.94481f
C4144 VSSD.t1157 VSUBS 0.839305f
C4145 VSSD.t64 VSUBS 1.90956f
C4146 VSSD.t886 VSUBS 1.97152f
C4147 VSSD.t955 VSUBS 1.07589f
C4148 VSSD.t563 VSUBS 1.47582f
C4149 VSSD.t888 VSUBS 1.34063f
C4150 VSSD.t164 VSUBS 1.14912f
C4151 VSSD.t709 VSUBS 1.3012f
C4152 VSSD.t977 VSUBS 1.17165f
C4153 VSSD.t954 VSUBS 1.15475f
C4154 VSSD.t868 VSUBS 1.38006f
C4155 VSSD.t166 VSUBS 1.3519f
C4156 VSSD.t764 VSUBS 1.68424f
C4157 VSSD.t313 VSUBS 1.64481f
C4158 VSSD.t311 VSUBS 1.21108f
C4159 VSSD.t1188 VSUBS 0.839305f
C4160 VSSD.t438 VSUBS 1.90956f
C4161 VSSD.t44 VSUBS 1.97152f
C4162 VSSD.t440 VSUBS 1.07589f
C4163 VSSD.t451 VSUBS 1.47582f
C4164 VSSD.t197 VSUBS 1.34063f
C4165 VSSD.t693 VSUBS 1.14912f
C4166 VSSD.t176 VSUBS 1.3012f
C4167 VSSD.t450 VSUBS 1.17165f
C4168 VSSD.t1112 VSUBS 1.15475f
C4169 VSSD.t596 VSUBS 1.38006f
C4170 VSSD.t280 VSUBS 1.3519f
C4171 VSSD.t988 VSUBS 1.68424f
C4172 VSSD.t598 VSUBS 1.64481f
C4173 VSSD.t594 VSUBS 1.21108f
C4174 VSSD.t1114 VSUBS 0.839305f
C4175 VSSD.t931 VSUBS 1.90956f
C4176 VSSD.t633 VSUBS 1.97152f
C4177 VSSD.t374 VSUBS 1.07589f
C4178 VSSD.t737 VSUBS 1.47582f
C4179 VSSD.t93 VSUBS 1.34063f
C4180 VSSD.t9 VSUBS 1.14912f
C4181 VSSD.t301 VSUBS 1.3012f
C4182 VSSD.t738 VSUBS 1.17165f
C4183 VSSD.t94 VSUBS 1.15475f
C4184 VSSD.t430 VSUBS 1.38006f
C4185 VSSD.t1167 VSUBS 1.3519f
C4186 VSSD.t837 VSUBS 1.68424f
C4187 VSSD.t434 VSUBS 1.64481f
C4188 VSSD.t432 VSUBS 1.21108f
C4189 VSSD.t1116 VSUBS 0.839305f
C4190 VSSD.t491 VSUBS 1.90956f
C4191 VSSD.t979 VSUBS 1.97152f
C4192 VSSD.t604 VSUBS 1.07589f
C4193 VSSD.t1166 VSUBS 1.47582f
C4194 VSSD.t330 VSUBS 1.34063f
C4195 VSSD.t1173 VSUBS 1.14912f
C4196 VSSD.t487 VSUBS 1.3012f
C4197 VSSD.t576 VSUBS 1.17165f
C4198 VSSD.t490 VSUBS 1.15475f
C4199 VSSD.t532 VSUBS 1.38006f
C4200 VSSD.t517 VSUBS 1.3519f
C4201 VSSD.t343 VSUBS 1.68424f
C4202 VSSD.t264 VSUBS 1.64481f
C4203 VSSD.t262 VSUBS 1.21108f
C4204 VSSD.t206 VSUBS 0.839305f
C4205 VSSD.t409 VSUBS 1.90956f
C4206 VSSD.t768 VSUBS 1.97152f
C4207 VSSD.t719 VSUBS 1.07589f
C4208 VSSD.t577 VSUBS 1.47582f
C4209 VSSD.t108 VSUBS 1.34063f
C4210 VSSD.t188 VSUBS 1.14912f
C4211 VSSD.t476 VSUBS 1.3012f
C4212 VSSD.t763 VSUBS 1.17165f
C4213 VSSD.t408 VSUBS 1.15475f
C4214 VSSD.t479 VSUBS 1.38006f
C4215 VSSD.t1000 VSUBS 1.3519f
C4216 VSSD.t242 VSUBS 1.68424f
C4217 VSSD.t481 VSUBS 1.64481f
C4218 VSSD.t751 VSUBS 1.81943f
C4219 VSSD.t874 VSUBS 1.95462f
C4220 VSSD.t1080 VSUBS 1.08152f
C4221 VSSD.t760 VSUBS 0.85057f
C4222 VSSD.n1386 VSUBS 0.023423f
C4223 VSSD.n1387 VSUBS 0.027816f
C4224 VSSD.n1388 VSUBS 0.023607f
C4225 VSSD.n1390 VSUBS 0.03123f
C4226 VSSD.n1392 VSUBS 0.03123f
C4227 VSSD.t1001 VSUBS 0.010396f
C4228 VSSD.n1393 VSUBS 0.018748f
C4229 VSSD.n1394 VSUBS 0.018565f
C4230 VSSD.n1395 VSUBS 0.011061f
C4231 VSSD.n1396 VSUBS 0.03123f
C4232 VSSD.n1397 VSUBS 0.011061f
C4233 VSSD.n1398 VSUBS 0.03123f
C4234 VSSD.t769 VSUBS 0.024724f
C4235 VSSD.n1399 VSUBS 0.038296f
C4236 VSSD.n1400 VSUBS 0.03123f
C4237 VSSD.t263 VSUBS 0.024414f
C4238 VSSD.n1401 VSUBS 0.040253f
C4239 VSSD.n1402 VSUBS 0.03123f
C4240 VSSD.n1403 VSUBS 0.011061f
C4241 VSSD.n1404 VSUBS 0.03123f
C4242 VSSD.n1405 VSUBS 0.011061f
C4243 VSSD.n1406 VSUBS 0.03123f
C4244 VSSD.n1407 VSUBS 0.011061f
C4245 VSSD.n1408 VSUBS 0.03123f
C4246 VSSD.n1410 VSUBS 0.03123f
C4247 VSSD.n1412 VSUBS 0.03123f
C4248 VSSD.n1414 VSUBS 0.03123f
C4249 VSSD.n1415 VSUBS 0.011061f
C4250 VSSD.n1416 VSUBS 0.03123f
C4251 VSSD.t302 VSUBS 0.013879f
C4252 VSSD.n1417 VSUBS 0.017846f
C4253 VSSD.n1418 VSUBS 0.029746f
C4254 VSSD.n1419 VSUBS 0.03123f
C4255 VSSD.n1420 VSUBS 0.011061f
C4256 VSSD.n1421 VSUBS 0.03123f
C4257 VSSD.n1423 VSUBS 0.018501f
C4258 VSSD.n1425 VSUBS 0.03123f
C4259 VSSD.n1427 VSUBS 0.03123f
C4260 VSSD.t281 VSUBS 0.010396f
C4261 VSSD.n1428 VSUBS 0.018748f
C4262 VSSD.n1429 VSUBS 0.018565f
C4263 VSSD.n1430 VSUBS 0.011061f
C4264 VSSD.n1431 VSUBS 0.03123f
C4265 VSSD.n1432 VSUBS 0.011061f
C4266 VSSD.n1433 VSUBS 0.03123f
C4267 VSSD.t45 VSUBS 0.024724f
C4268 VSSD.n1434 VSUBS 0.038296f
C4269 VSSD.n1435 VSUBS 0.03123f
C4270 VSSD.t312 VSUBS 0.024414f
C4271 VSSD.n1436 VSUBS 0.040253f
C4272 VSSD.n1437 VSUBS 0.03123f
C4273 VSSD.n1438 VSUBS 0.011061f
C4274 VSSD.n1439 VSUBS 0.03123f
C4275 VSSD.n1440 VSUBS 0.011061f
C4276 VSSD.n1441 VSUBS 0.03123f
C4277 VSSD.n1442 VSUBS 0.011061f
C4278 VSSD.n1443 VSUBS 0.03123f
C4279 VSSD.n1445 VSUBS 0.037186f
C4280 VSSD.n1446 VSUBS 0.030066f
C4281 VSSD.n1448 VSUBS 0.034526f
C4282 VSSD.t887 VSUBS 0.024724f
C4283 VSSD.n1450 VSUBS 0.038296f
C4284 VSSD.n1451 VSUBS 0.03123f
C4285 VSSD.n1452 VSUBS 0.03123f
C4286 VSSD.n1453 VSUBS 0.03123f
C4287 VSSD.n1454 VSUBS 0.011061f
C4288 VSSD.n1455 VSUBS 0.011061f
C4289 VSSD.n1456 VSUBS 0.011061f
C4290 VSSD.n1457 VSUBS 0.03123f
C4291 VSSD.n1458 VSUBS 0.03123f
C4292 VSSD.n1459 VSUBS 0.03123f
C4293 VSSD.t710 VSUBS 0.013879f
C4294 VSSD.n1461 VSUBS 0.017846f
C4295 VSSD.n1462 VSUBS 0.029746f
C4296 VSSD.n1464 VSUBS 0.011061f
C4297 VSSD.n1465 VSUBS 0.03123f
C4298 VSSD.n1466 VSUBS 0.03123f
C4299 VSSD.n1467 VSUBS 0.03123f
C4300 VSSD.n1468 VSUBS 0.011061f
C4301 VSSD.t167 VSUBS 0.010396f
C4302 VSSD.n1470 VSUBS 0.018748f
C4303 VSSD.n1471 VSUBS 0.018565f
C4304 VSSD.n1473 VSUBS 0.03123f
C4305 VSSD.n1474 VSUBS 0.03123f
C4306 VSSD.n1475 VSUBS 0.03123f
C4307 VSSD.t314 VSUBS 0.028005f
C4308 VSSD.n1477 VSUBS 0.036086f
C4309 VSSD.n1479 VSUBS 0.03123f
C4310 VSSD.n1480 VSUBS 0.023423f
C4311 VSSD.n1481 VSUBS 0.018501f
C4312 VSSD.n1484 VSUBS 0.031818f
C4313 VSSD.n1486 VSUBS 0.03123f
C4314 VSSD.n1487 VSUBS 0.03123f
C4315 VSSD.n1488 VSUBS 0.03123f
C4316 VSSD.n1490 VSUBS 0.011061f
C4317 VSSD.n1491 VSUBS 0.011061f
C4318 VSSD.n1492 VSUBS 0.03123f
C4319 VSSD.n1493 VSUBS 0.03123f
C4320 VSSD.n1494 VSUBS 0.03123f
C4321 VSSD.n1495 VSUBS 0.011061f
C4322 VSSD.t177 VSUBS 0.013879f
C4323 VSSD.n1497 VSUBS 0.017846f
C4324 VSSD.n1498 VSUBS 0.029746f
C4325 VSSD.n1500 VSUBS 0.03123f
C4326 VSSD.n1501 VSUBS 0.03123f
C4327 VSSD.n1502 VSUBS 0.03123f
C4328 VSSD.n1503 VSUBS 0.011061f
C4329 VSSD.n1504 VSUBS 0.011061f
C4330 VSSD.n1506 VSUBS 0.03123f
C4331 VSSD.n1507 VSUBS 0.03123f
C4332 VSSD.n1508 VSUBS 0.03123f
C4333 VSSD.n1509 VSUBS 0.011061f
C4334 VSSD.t599 VSUBS 0.028005f
C4335 VSSD.n1511 VSUBS 0.036086f
C4336 VSSD.n1512 VSUBS 0.03123f
C4337 VSSD.n1513 VSUBS 0.03123f
C4338 VSSD.n1514 VSUBS 0.023423f
C4339 VSSD.t595 VSUBS 0.024414f
C4340 VSSD.n1515 VSUBS 0.040253f
C4341 VSSD.n1518 VSUBS 0.031818f
C4342 VSSD.n1519 VSUBS 0.03123f
C4343 VSSD.n1520 VSUBS 0.03123f
C4344 VSSD.n1521 VSUBS 0.03123f
C4345 VSSD.t634 VSUBS 0.024724f
C4346 VSSD.n1522 VSUBS 0.038296f
C4347 VSSD.n1524 VSUBS 0.011061f
C4348 VSSD.n1525 VSUBS 0.03123f
C4349 VSSD.n1526 VSUBS 0.03123f
C4350 VSSD.n1527 VSUBS 0.03123f
C4351 VSSD.n1528 VSUBS 0.011061f
C4352 VSSD.n1529 VSUBS 0.011061f
C4353 VSSD.n1531 VSUBS 0.03123f
C4354 VSSD.n1532 VSUBS 0.03123f
C4355 VSSD.n1534 VSUBS 0.011061f
C4356 VSSD.n1535 VSUBS 0.011061f
C4357 VSSD.n1536 VSUBS 0.03123f
C4358 VSSD.n1537 VSUBS 0.03123f
C4359 VSSD.n1538 VSUBS 0.03123f
C4360 VSSD.t1168 VSUBS 0.010396f
C4361 VSSD.n1540 VSUBS 0.018748f
C4362 VSSD.n1541 VSUBS 0.018565f
C4363 VSSD.n1543 VSUBS 0.011061f
C4364 VSSD.n1544 VSUBS 0.03123f
C4365 VSSD.n1545 VSUBS 0.03123f
C4366 VSSD.n1546 VSUBS 0.03123f
C4367 VSSD.t435 VSUBS 0.028005f
C4368 VSSD.n1547 VSUBS 0.036086f
C4369 VSSD.t433 VSUBS 0.024414f
C4370 VSSD.n1549 VSUBS 0.040253f
C4371 VSSD.n1550 VSUBS 0.023423f
C4372 VSSD.n1551 VSUBS 0.018501f
C4373 VSSD.n1552 VSUBS 0.03123f
C4374 VSSD.n1554 VSUBS 0.031818f
C4375 VSSD.t980 VSUBS 0.024724f
C4376 VSSD.n1556 VSUBS 0.038296f
C4377 VSSD.n1557 VSUBS 0.03123f
C4378 VSSD.n1558 VSUBS 0.03123f
C4379 VSSD.n1559 VSUBS 0.03123f
C4380 VSSD.n1560 VSUBS 0.011061f
C4381 VSSD.n1561 VSUBS 0.011061f
C4382 VSSD.n1562 VSUBS 0.011061f
C4383 VSSD.n1563 VSUBS 0.03123f
C4384 VSSD.n1564 VSUBS 0.03123f
C4385 VSSD.n1565 VSUBS 0.03123f
C4386 VSSD.t488 VSUBS 0.013879f
C4387 VSSD.n1567 VSUBS 0.017846f
C4388 VSSD.n1568 VSUBS 0.029746f
C4389 VSSD.n1570 VSUBS 0.011061f
C4390 VSSD.n1571 VSUBS 0.03123f
C4391 VSSD.n1572 VSUBS 0.03123f
C4392 VSSD.n1573 VSUBS 0.03123f
C4393 VSSD.n1574 VSUBS 0.011061f
C4394 VSSD.t518 VSUBS 0.010396f
C4395 VSSD.n1576 VSUBS 0.018748f
C4396 VSSD.n1577 VSUBS 0.018565f
C4397 VSSD.n1579 VSUBS 0.03123f
C4398 VSSD.n1580 VSUBS 0.03123f
C4399 VSSD.n1581 VSUBS 0.03123f
C4400 VSSD.t265 VSUBS 0.028005f
C4401 VSSD.n1583 VSUBS 0.036086f
C4402 VSSD.n1585 VSUBS 0.03123f
C4403 VSSD.n1586 VSUBS 0.023423f
C4404 VSSD.n1587 VSUBS 0.018501f
C4405 VSSD.n1590 VSUBS 0.031818f
C4406 VSSD.n1592 VSUBS 0.03123f
C4407 VSSD.n1593 VSUBS 0.03123f
C4408 VSSD.n1594 VSUBS 0.03123f
C4409 VSSD.n1596 VSUBS 0.011061f
C4410 VSSD.n1597 VSUBS 0.011061f
C4411 VSSD.n1598 VSUBS 0.03123f
C4412 VSSD.n1599 VSUBS 0.03123f
C4413 VSSD.n1600 VSUBS 0.03123f
C4414 VSSD.n1601 VSUBS 0.011061f
C4415 VSSD.t477 VSUBS 0.013879f
C4416 VSSD.n1603 VSUBS 0.017846f
C4417 VSSD.n1604 VSUBS 0.029746f
C4418 VSSD.n1606 VSUBS 0.03123f
C4419 VSSD.n1607 VSUBS 0.03123f
C4420 VSSD.n1608 VSUBS 0.03123f
C4421 VSSD.n1609 VSUBS 0.011061f
C4422 VSSD.n1610 VSUBS 0.011061f
C4423 VSSD.n1612 VSUBS 0.03123f
C4424 VSSD.n1613 VSUBS 0.03123f
C4425 VSSD.n1614 VSUBS 0.03123f
C4426 VSSD.n1615 VSUBS 0.011061f
C4427 VSSD.t482 VSUBS 0.028005f
C4428 VSSD.n1617 VSUBS 0.036086f
C4429 VSSD.n1618 VSUBS 0.03123f
C4430 VSSD.n1619 VSUBS 0.03123f
C4431 VSSD.n1620 VSUBS 0.023253f
C4432 VSSD.t752 VSUBS 0.024414f
C4433 VSSD.n1621 VSUBS 0.040193f
C4434 VSSD.n1624 VSUBS 0.03123f
C4435 VSSD.n1625 VSUBS 0.03123f
C4436 VSSD.n1626 VSUBS 0.028345f
C4437 VSSD.n1627 VSUBS 0.013402f
C4438 VSSD.n1628 VSUBS 0.778863f
C4439 VSSD.n1629 VSUBS 23.913f
C4440 VSSD.n1630 VSUBS 0.131045p
C4441 VSSD.n1631 VSUBS 56.717396f
C4442 VSSD.n1632 VSUBS 0.667373f
C4443 VSSD.n1633 VSUBS 0.028345f
C4444 VSSD.n1634 VSUBS 0.013402f
C4445 VSSD.n1636 VSUBS 0.027816f
C4446 VSSD.n1637 VSUBS 0.023607f
C4447 VSSD.n1639 VSUBS 0.03123f
C4448 VSSD.n1640 VSUBS 0.023423f
C4449 VSSD.n1641 VSUBS 0.010523f
C4450 VSSD.n1644 VSUBS 0.031818f
C4451 VSSD.n1645 VSUBS 0.028345f
C4452 VSSD.n1646 VSUBS 0.03123f
C4453 VSSD.n1647 VSUBS 0.03123f
C4454 VSSD.n1648 VSUBS 0.038296f
C4455 VSSD.n1650 VSUBS 0.011061f
C4456 VSSD.n1651 VSUBS 0.03123f
C4457 VSSD.n1652 VSUBS 0.03123f
C4458 VSSD.n1653 VSUBS 0.03123f
C4459 VSSD.n1654 VSUBS 0.011061f
C4460 VSSD.n1655 VSUBS 0.011061f
C4461 VSSD.n1657 VSUBS 0.03123f
C4462 VSSD.n1658 VSUBS 0.03123f
C4463 VSSD.n1660 VSUBS 0.011061f
C4464 VSSD.n1661 VSUBS 0.011061f
C4465 VSSD.n1662 VSUBS 0.03123f
C4466 VSSD.n1663 VSUBS 0.03123f
C4467 VSSD.n1664 VSUBS 0.03123f
C4468 VSSD.t624 VSUBS 0.010396f
C4469 VSSD.n1666 VSUBS 0.018748f
C4470 VSSD.n1667 VSUBS 0.018565f
C4471 VSSD.n1669 VSUBS 0.011061f
C4472 VSSD.n1670 VSUBS 0.03123f
C4473 VSSD.n1671 VSUBS 0.03123f
C4474 VSSD.n1672 VSUBS 0.03123f
C4475 VSSD.n1673 VSUBS 0.036086f
C4476 VSSD.t146 VSUBS 0.024414f
C4477 VSSD.n1675 VSUBS 0.040253f
C4478 VSSD.n1676 VSUBS 0.023423f
C4479 VSSD.n1677 VSUBS 0.010693f
C4480 VSSD.n1678 VSUBS 0.028345f
C4481 VSSD.n1679 VSUBS 0.031818f
C4482 VSSD.t653 VSUBS 0.024724f
C4483 VSSD.n1681 VSUBS 0.038296f
C4484 VSSD.n1682 VSUBS 0.03123f
C4485 VSSD.n1683 VSUBS 0.03123f
C4486 VSSD.n1684 VSUBS 0.03123f
C4487 VSSD.n1685 VSUBS 0.011061f
C4488 VSSD.n1686 VSUBS 0.011061f
C4489 VSSD.n1687 VSUBS 0.011061f
C4490 VSSD.n1688 VSUBS 0.03123f
C4491 VSSD.n1689 VSUBS 0.03123f
C4492 VSSD.n1690 VSUBS 0.03123f
C4493 VSSD.t486 VSUBS 0.013879f
C4494 VSSD.n1692 VSUBS 0.017846f
C4495 VSSD.n1693 VSUBS 0.029746f
C4496 VSSD.n1695 VSUBS 0.011061f
C4497 VSSD.n1696 VSUBS 0.03123f
C4498 VSSD.n1697 VSUBS 0.03123f
C4499 VSSD.n1698 VSUBS 0.03123f
C4500 VSSD.n1699 VSUBS 0.011061f
C4501 VSSD.t14 VSUBS 0.010396f
C4502 VSSD.n1701 VSUBS 0.018748f
C4503 VSSD.n1702 VSUBS 0.018565f
C4504 VSSD.n1704 VSUBS 0.03123f
C4505 VSSD.n1705 VSUBS 0.03123f
C4506 VSSD.n1706 VSUBS 0.03123f
C4507 VSSD.t907 VSUBS 0.028005f
C4508 VSSD.n1708 VSUBS 0.036086f
C4509 VSSD.n1710 VSUBS 0.03123f
C4510 VSSD.n1711 VSUBS 0.023423f
C4511 VSSD.n1712 VSUBS 0.010693f
C4512 VSSD.n1715 VSUBS 0.031818f
C4513 VSSD.n1716 VSUBS 0.028345f
C4514 VSSD.n1717 VSUBS 0.03123f
C4515 VSSD.n1718 VSUBS 0.03123f
C4516 VSSD.n1719 VSUBS 0.038296f
C4517 VSSD.n1721 VSUBS 0.011061f
C4518 VSSD.n1722 VSUBS 0.03123f
C4519 VSSD.n1723 VSUBS 0.03123f
C4520 VSSD.n1724 VSUBS 0.03123f
C4521 VSSD.n1725 VSUBS 0.011061f
C4522 VSSD.n1726 VSUBS 0.011061f
C4523 VSSD.n1728 VSUBS 0.03123f
C4524 VSSD.n1729 VSUBS 0.03123f
C4525 VSSD.n1731 VSUBS 0.011061f
C4526 VSSD.n1732 VSUBS 0.011061f
C4527 VSSD.n1733 VSUBS 0.03123f
C4528 VSSD.n1734 VSUBS 0.03123f
C4529 VSSD.n1735 VSUBS 0.03123f
C4530 VSSD.t999 VSUBS 0.010396f
C4531 VSSD.n1737 VSUBS 0.018748f
C4532 VSSD.n1738 VSUBS 0.018565f
C4533 VSSD.n1740 VSUBS 0.011061f
C4534 VSSD.n1741 VSUBS 0.03123f
C4535 VSSD.n1742 VSUBS 0.03123f
C4536 VSSD.n1743 VSUBS 0.03123f
C4537 VSSD.n1744 VSUBS 0.036086f
C4538 VSSD.t662 VSUBS 0.024414f
C4539 VSSD.n1746 VSUBS 0.040253f
C4540 VSSD.n1747 VSUBS 0.023423f
C4541 VSSD.n1748 VSUBS 0.010693f
C4542 VSSD.n1749 VSUBS 0.028345f
C4543 VSSD.n1750 VSUBS 0.031818f
C4544 VSSD.t1153 VSUBS 0.024724f
C4545 VSSD.n1752 VSUBS 0.038296f
C4546 VSSD.n1753 VSUBS 0.03123f
C4547 VSSD.n1754 VSUBS 0.03123f
C4548 VSSD.n1755 VSUBS 0.03123f
C4549 VSSD.n1756 VSUBS 0.011061f
C4550 VSSD.n1757 VSUBS 0.011061f
C4551 VSSD.n1758 VSUBS 0.011061f
C4552 VSSD.n1759 VSUBS 0.03123f
C4553 VSSD.n1760 VSUBS 0.03123f
C4554 VSSD.n1761 VSUBS 0.03123f
C4555 VSSD.t1145 VSUBS 0.013879f
C4556 VSSD.n1763 VSUBS 0.017846f
C4557 VSSD.n1764 VSUBS 0.029746f
C4558 VSSD.n1766 VSUBS 0.011061f
C4559 VSSD.n1767 VSUBS 0.03123f
C4560 VSSD.n1768 VSUBS 0.03123f
C4561 VSSD.n1769 VSUBS 0.03123f
C4562 VSSD.n1770 VSUBS 0.011061f
C4563 VSSD.t1127 VSUBS 0.010396f
C4564 VSSD.n1772 VSUBS 0.018748f
C4565 VSSD.n1773 VSUBS 0.018565f
C4566 VSSD.n1775 VSUBS 0.03123f
C4567 VSSD.n1776 VSUBS 0.03123f
C4568 VSSD.n1777 VSUBS 0.03123f
C4569 VSSD.t253 VSUBS 0.028005f
C4570 VSSD.n1779 VSUBS 0.036086f
C4571 VSSD.n1781 VSUBS 0.03123f
C4572 VSSD.n1782 VSUBS 0.023423f
C4573 VSSD.n1783 VSUBS 0.010693f
C4574 VSSD.n1786 VSUBS 0.031818f
C4575 VSSD.n1787 VSUBS 0.028345f
C4576 VSSD.n1788 VSUBS 0.03123f
C4577 VSSD.n1789 VSUBS 0.03123f
C4578 VSSD.n1790 VSUBS 0.038296f
C4579 VSSD.n1792 VSUBS 0.011061f
C4580 VSSD.n1793 VSUBS 0.03123f
C4581 VSSD.n1794 VSUBS 0.03123f
C4582 VSSD.n1795 VSUBS 0.03123f
C4583 VSSD.n1796 VSUBS 0.011061f
C4584 VSSD.n1797 VSUBS 0.011061f
C4585 VSSD.n1799 VSUBS 0.03123f
C4586 VSSD.n1800 VSUBS 0.03123f
C4587 VSSD.n1802 VSUBS 0.011061f
C4588 VSSD.n1803 VSUBS 0.011061f
C4589 VSSD.n1804 VSUBS 0.03123f
C4590 VSSD.n1805 VSUBS 0.03123f
C4591 VSSD.n1806 VSUBS 0.03123f
C4592 VSSD.t275 VSUBS 0.010396f
C4593 VSSD.n1808 VSUBS 0.018748f
C4594 VSSD.n1809 VSUBS 0.018565f
C4595 VSSD.n1811 VSUBS 0.011061f
C4596 VSSD.n1812 VSUBS 0.03123f
C4597 VSSD.n1813 VSUBS 0.03123f
C4598 VSSD.n1814 VSUBS 0.03123f
C4599 VSSD.n1815 VSUBS 0.036086f
C4600 VSSD.t640 VSUBS 0.024414f
C4601 VSSD.n1817 VSUBS 0.032619f
C4602 VSSD.n1818 VSUBS 0.023423f
C4603 VSSD.n1819 VSUBS 2.61656f
C4604 VSSD.n1820 VSUBS 1.76436f
C4605 VSSD.n1821 VSUBS 0.215918f
C4606 VSSD.n1822 VSUBS 1.71988f
C4607 VSSD.n1823 VSUBS 0.812406f
C4608 VSSD.n1824 VSUBS 0.214921f
C4609 VSSD.n1825 VSUBS 2.62148f
C4610 VSSD.n1826 VSUBS 0.812406f
C4611 VSSD.n1827 VSUBS 1.13383f
C4612 VSSD.n1828 VSUBS 2.51964f
C4613 VSSD.n1829 VSUBS 0.036513f
C4614 VSSD.t856 VSUBS 0.02316f
C4615 VSSD.n1830 VSUBS 0.055953f
C4616 VSSD.n1832 VSUBS 0.037564f
C4617 VSSD.n1833 VSUBS 0.03123f
C4618 VSSD.n1834 VSUBS 0.03123f
C4619 VSSD.n1836 VSUBS 0.01373f
C4620 VSSD.n1837 VSUBS 0.030584f
C4621 VSSD.n1840 VSUBS 0.03123f
C4622 VSSD.n1841 VSUBS 0.03123f
C4623 VSSD.n1842 VSUBS 0.03123f
C4624 VSSD.n1843 VSUBS 0.01373f
C4625 VSSD.n1844 VSUBS 0.036114f
C4626 VSSD.n1846 VSUBS 0.01373f
C4627 VSSD.n1847 VSUBS 0.036114f
C4628 VSSD.n1848 VSUBS 0.028175f
C4629 VSSD.n1849 VSUBS 0.010693f
C4630 VSSD.n1850 VSUBS 0.018501f
C4631 VSSD.t911 VSUBS 0.024414f
C4632 VSSD.n1851 VSUBS 0.038089f
C4633 VSSD.n1853 VSUBS 0.02785f
C4634 VSSD.t915 VSUBS 0.028005f
C4635 VSSD.n1854 VSUBS 0.03344f
C4636 VSSD.n1855 VSUBS 0.03123f
C4637 VSSD.n1856 VSUBS 0.03123f
C4638 VSSD.n1857 VSUBS 0.03123f
C4639 VSSD.t1084 VSUBS 0.010396f
C4640 VSSD.n1860 VSUBS 0.018748f
C4641 VSSD.n1861 VSUBS 0.018565f
C4642 VSSD.n1863 VSUBS 0.03123f
C4643 VSSD.n1864 VSUBS 0.03123f
C4644 VSSD.n1865 VSUBS 0.03123f
C4645 VSSD.n1866 VSUBS 0.011061f
C4646 VSSD.t403 VSUBS 0.013879f
C4647 VSSD.n1868 VSUBS 0.017846f
C4648 VSSD.n1869 VSUBS 0.029746f
C4649 VSSD.n1871 VSUBS 0.03123f
C4650 VSSD.n1872 VSUBS 0.03123f
C4651 VSSD.n1873 VSUBS 0.03123f
C4652 VSSD.n1874 VSUBS 0.011061f
C4653 VSSD.n1875 VSUBS 0.011061f
C4654 VSSD.n1877 VSUBS 0.03123f
C4655 VSSD.n1878 VSUBS 0.03123f
C4656 VSSD.t84 VSUBS 0.024724f
C4657 VSSD.n1881 VSUBS 0.036733f
C4658 VSSD.n1882 VSUBS 0.03123f
C4659 VSSD.n1883 VSUBS 0.03123f
C4660 VSSD.n1884 VSUBS 0.028345f
C4661 VSSD.n1885 VSUBS 0.02785f
C4662 VSSD.n1886 VSUBS 0.037007f
C4663 VSSD.n1887 VSUBS 0.037007f
C4664 VSSD.n1888 VSUBS 0.02785f
C4665 VSSD.n1889 VSUBS 0.03344f
C4666 VSSD.n1890 VSUBS 0.03123f
C4667 VSSD.n1891 VSUBS 0.03123f
C4668 VSSD.n1892 VSUBS 0.03123f
C4669 VSSD.n1895 VSUBS 0.018565f
C4670 VSSD.n1897 VSUBS 0.03123f
C4671 VSSD.n1898 VSUBS 0.03123f
C4672 VSSD.n1899 VSUBS 0.03123f
C4673 VSSD.n1900 VSUBS 0.011061f
C4674 VSSD.n1902 VSUBS 0.029746f
C4675 VSSD.n1904 VSUBS 0.03123f
C4676 VSSD.n1905 VSUBS 0.03123f
C4677 VSSD.n1906 VSUBS 0.03123f
C4678 VSSD.n1907 VSUBS 0.011061f
C4679 VSSD.n1908 VSUBS 0.011061f
C4680 VSSD.n1910 VSUBS 0.03123f
C4681 VSSD.n1911 VSUBS 0.03123f
C4682 VSSD.n1912 VSUBS 0.03123f
C4683 VSSD.n1914 VSUBS 0.036733f
C4684 VSSD.n1915 VSUBS 0.03344f
C4685 VSSD.n1916 VSUBS 0.02785f
C4686 VSSD.n1917 VSUBS 0.037007f
C4687 VSSD.n1918 VSUBS 0.037007f
C4688 VSSD.n1919 VSUBS 0.02785f
C4689 VSSD.n1920 VSUBS 0.03344f
C4690 VSSD.n1921 VSUBS 0.03123f
C4691 VSSD.n1922 VSUBS 0.03123f
C4692 VSSD.n1923 VSUBS 0.03123f
C4693 VSSD.n1926 VSUBS 0.018565f
C4694 VSSD.n1928 VSUBS 0.03123f
C4695 VSSD.n1929 VSUBS 0.03123f
C4696 VSSD.n1930 VSUBS 0.03123f
C4697 VSSD.n1931 VSUBS 0.011061f
C4698 VSSD.n1933 VSUBS 0.029746f
C4699 VSSD.n1935 VSUBS 0.03123f
C4700 VSSD.n1936 VSUBS 0.03123f
C4701 VSSD.n1937 VSUBS 0.03123f
C4702 VSSD.n1938 VSUBS 0.011061f
C4703 VSSD.n1939 VSUBS 0.011061f
C4704 VSSD.n1941 VSUBS 0.03123f
C4705 VSSD.n1942 VSUBS 0.03123f
C4706 VSSD.n1943 VSUBS 0.03123f
C4707 VSSD.n1945 VSUBS 0.036733f
C4708 VSSD.n1946 VSUBS 0.03344f
C4709 VSSD.n1947 VSUBS 0.02785f
C4710 VSSD.n1948 VSUBS 0.037007f
C4711 VSSD.n1949 VSUBS 0.037007f
C4712 VSSD.n1950 VSUBS 0.02785f
C4713 VSSD.n1951 VSUBS 0.03344f
C4714 VSSD.n1952 VSUBS 0.03123f
C4715 VSSD.n1953 VSUBS 0.03123f
C4716 VSSD.n1954 VSUBS 0.03123f
C4717 VSSD.n1957 VSUBS 0.018565f
C4718 VSSD.n1959 VSUBS 0.03123f
C4719 VSSD.n1960 VSUBS 0.03123f
C4720 VSSD.n1961 VSUBS 0.03123f
C4721 VSSD.n1962 VSUBS 0.011061f
C4722 VSSD.n1964 VSUBS 0.029746f
C4723 VSSD.n1966 VSUBS 0.03123f
C4724 VSSD.n1967 VSUBS 0.03123f
C4725 VSSD.n1968 VSUBS 0.03123f
C4726 VSSD.n1969 VSUBS 0.011061f
C4727 VSSD.n1970 VSUBS 0.011061f
C4728 VSSD.n1972 VSUBS 0.03123f
C4729 VSSD.n1973 VSUBS 0.03123f
C4730 VSSD.n1974 VSUBS 0.03123f
C4731 VSSD.n1976 VSUBS 0.036733f
C4732 VSSD.n1977 VSUBS 0.03344f
C4733 VSSD.n1978 VSUBS 0.02785f
C4734 VSSD.n1979 VSUBS 0.037007f
C4735 VSSD.n1980 VSUBS 0.037007f
C4736 VSSD.n1981 VSUBS 0.02785f
C4737 VSSD.n1982 VSUBS 0.03344f
C4738 VSSD.n1983 VSUBS 0.03123f
C4739 VSSD.n1984 VSUBS 0.03123f
C4740 VSSD.n1985 VSUBS 0.03123f
C4741 VSSD.n1988 VSUBS 0.018565f
C4742 VSSD.n1990 VSUBS 0.03123f
C4743 VSSD.n1991 VSUBS 0.03123f
C4744 VSSD.n1992 VSUBS 0.03123f
C4745 VSSD.n1993 VSUBS 0.011061f
C4746 VSSD.n1995 VSUBS 0.029746f
C4747 VSSD.n1997 VSUBS 0.03123f
C4748 VSSD.n1998 VSUBS 0.03123f
C4749 VSSD.n1999 VSUBS 0.03123f
C4750 VSSD.n2000 VSUBS 0.011061f
C4751 VSSD.n2001 VSUBS 0.011061f
C4752 VSSD.n2003 VSUBS 0.03123f
C4753 VSSD.n2004 VSUBS 0.03123f
C4754 VSSD.n2005 VSUBS 0.03123f
C4755 VSSD.n2007 VSUBS 0.036733f
C4756 VSSD.n2008 VSUBS 0.03344f
C4757 VSSD.n2009 VSUBS 0.02785f
C4758 VSSD.n2010 VSUBS 0.030515f
C4759 VSSD.n2011 VSUBS 0.050341f
C4760 VSSD.n2012 VSUBS 0.641674f
C4761 VSSD.t650 VSUBS 0.035993f
C4762 VSSD.t292 VSUBS 0.077524f
C4763 VSSD.t391 VSUBS 0.077524f
C4764 VSSD.t290 VSUBS 0.199348f
C4765 VSSD.t1160 VSUBS 0.227958f
C4766 VSSD.t182 VSUBS 0.083985f
C4767 VSSD.t1086 VSUBS 0.087676f
C4768 VSSD.t393 VSUBS 0.128284f
C4769 VSSD.t668 VSUBS 0.097828f
C4770 VSSD.t665 VSUBS 0.097828f
C4771 VSSD.t969 VSUBS 0.143974f
C4772 VSSD.t297 VSUBS 0.100597f
C4773 VSSD.t950 VSUBS 0.066449f
C4774 VSSD.t1051 VSUBS 0.091368f
C4775 VSSD.t400 VSUBS 0.121824f
C4776 VSSD.t91 VSUBS 0.121824f
C4777 VSSD.t1093 VSUBS 0.091368f
C4778 VSSD.t667 VSUBS 0.066449f
C4779 VSSD.t1143 VSUBS 0.100597f
C4780 VSSD.t1004 VSUBS 0.143974f
C4781 VSSD.t386 VSUBS 0.097828f
C4782 VSSD.t949 VSUBS 0.097828f
C4783 VSSD.t508 VSUBS 0.128284f
C4784 VSSD.t1088 VSUBS 0.087676f
C4785 VSSD.t574 VSUBS 0.083985f
C4786 VSSD.t1161 VSUBS 0.227958f
C4787 VSSD.t382 VSUBS 0.199348f
C4788 VSSD.t509 VSUBS 0.077524f
C4789 VSSD.t384 VSUBS 0.077524f
C4790 VSSD.t876 VSUBS 0.067372f
C4791 VSSD.t646 VSUBS 0.035993f
C4792 VSSD.t845 VSUBS 0.077524f
C4793 VSSD.t561 VSUBS 0.077524f
C4794 VSSD.t847 VSUBS 0.199348f
C4795 VSSD.t833 VSUBS 0.227958f
C4796 VSSD.t0 VSUBS 0.083985f
C4797 VSSD.t1091 VSUBS 0.087676f
C4798 VSSD.t1180 VSUBS 0.128284f
C4799 VSSD.t740 VSUBS 0.097828f
C4800 VSSD.t849 VSUBS 0.097828f
C4801 VSSD.t328 VSUBS 0.143974f
C4802 VSSD.t530 VSUBS 0.100597f
C4803 VSSD.t539 VSUBS 0.066449f
C4804 VSSD.t1016 VSUBS 0.091368f
C4805 VSSD.t39 VSUBS 0.121824f
C4806 VSSD.t540 VSUBS 0.121824f
C4807 VSSD.t1069 VSUBS 0.091368f
C4808 VSSD.t863 VSUBS 0.066449f
C4809 VSSD.t1154 VSUBS 0.100597f
C4810 VSSD.t1181 VSUBS 0.143974f
C4811 VSSD.t818 VSUBS 0.097828f
C4812 VSSD.t62 VSUBS 0.097828f
C4813 VSSD.t329 VSUBS 0.128284f
C4814 VSSD.t1063 VSUBS 0.087676f
C4815 VSSD.t776 VSUBS 0.083985f
C4816 VSSD.t96 VSUBS 0.227958f
C4817 VSSD.t814 VSUBS 0.199348f
C4818 VSSD.t682 VSUBS 0.077524f
C4819 VSSD.t816 VSUBS 0.077524f
C4820 VSSD.t472 VSUBS 0.067372f
C4821 VSSD.t822 VSUBS 0.035993f
C4822 VSSD.t553 VSUBS 0.077524f
C4823 VSSD.t232 VSUBS 0.077524f
C4824 VSSD.t180 VSUBS 0.199348f
C4825 VSSD.t872 VSUBS 0.227958f
C4826 VSSD.t656 VSUBS 0.083985f
C4827 VSSD.t1067 VSUBS 0.087676f
C4828 VSSD.t234 VSUBS 0.128284f
C4829 VSSD.t778 VSUBS 0.097828f
C4830 VSSD.t551 VSUBS 0.097828f
C4831 VSSD.t478 VSUBS 0.143974f
C4832 VSSD.t864 VSUBS 0.100597f
C4833 VSSD.t758 VSUBS 0.066449f
C4834 VSSD.t1032 VSUBS 0.091368f
C4835 VSSD.t195 VSUBS 0.121824f
C4836 VSSD.t701 VSUBS 0.121824f
C4837 VSSD.t1076 VSUBS 0.091368f
C4838 VSSD.t995 VSUBS 0.066449f
C4839 VSSD.t244 VSUBS 0.100597f
C4840 VSSD.t972 VSUBS 0.143974f
C4841 VSSD.t965 VSUBS 0.097828f
C4842 VSSD.t757 VSUBS 0.097828f
C4843 VSSD.t109 VSUBS 0.128284f
C4844 VSSD.t1043 VSUBS 0.087676f
C4845 VSSD.t525 VSUBS 0.083985f
C4846 VSSD.t996 VSUBS 0.227958f
C4847 VSSD.t989 VSUBS 0.199348f
C4848 VSSD.t110 VSUBS 0.077524f
C4849 VSSD.t991 VSUBS 0.077524f
C4850 VSSD.t648 VSUBS 0.067372f
C4851 VSSD.t305 VSUBS 0.035993f
C4852 VSSD.t1136 VSUBS 0.077524f
C4853 VSSD.t795 VSUBS 0.077524f
C4854 VSSD.t1138 VSUBS 0.199348f
C4855 VSSD.t901 VSUBS 0.227958f
C4856 VSSD.t544 VSUBS 0.083985f
C4857 VSSD.t1104 VSUBS 0.087676f
C4858 VSSD.t797 VSUBS 0.128284f
C4859 VSSD.t660 VSUBS 0.097828f
C4860 VSSD.t333 VSUBS 0.097828f
C4861 VSSD.t38 VSUBS 0.143974f
C4862 VSSD.t761 VSUBS 0.100597f
C4863 VSSD.t557 VSUBS 0.066449f
C4864 VSSD.t1101 VSUBS 0.091368f
C4865 VSSD.t717 VSUBS 0.121824f
C4866 VSSD.t411 VSUBS 0.121824f
C4867 VSSD.t1049 VSUBS 0.091368f
C4868 VSSD.t659 VSUBS 0.066449f
C4869 VSSD.t134 VSUBS 0.100597f
C4870 VSSD.t794 VSUBS 0.143974f
C4871 VSSD.t970 VSUBS 0.097828f
C4872 VSSD.t556 VSUBS 0.097828f
C4873 VSSD.t629 VSUBS 0.128284f
C4874 VSSD.t1107 VSUBS 0.087676f
C4875 VSSD.t254 VSUBS 0.083985f
C4876 VSSD.t199 VSUBS 0.227958f
C4877 VSSD.t788 VSUBS 0.199348f
C4878 VSSD.t36 VSUBS 0.077524f
C4879 VSSD.t973 VSUBS 0.077524f
C4880 VSSD.t644 VSUBS 0.067372f
C4881 VSSD.t470 VSUBS 0.035993f
C4882 VSSD.t219 VSUBS 0.077524f
C4883 VSSD.t495 VSUBS 0.077524f
C4884 VSSD.t217 VSUBS 0.199348f
C4885 VSSD.t953 VSUBS 0.227958f
C4886 VSSD.t83 VSUBS 0.083985f
C4887 VSSD.t1109 VSUBS 0.087676f
C4888 VSSD.t497 VSUBS 0.128284f
C4889 VSSD.t867 VSUBS 0.097828f
C4890 VSSD.t215 VSUBS 0.097828f
C4891 VSSD.t325 VSUBS 0.143974f
C4892 VSSD.t712 VSUBS 0.100597f
C4893 VSSD.t866 VSUBS 0.066449f
C4894 VSSD.t1056 VSUBS 0.091368f
C4895 VSSD.t402 VSUBS 0.121824f
C4896 VSSD.t1002 VSUBS 0.121824f
C4897 VSSD.t1010 VSUBS 0.091368f
C4898 VSSD.t927 VSUBS 0.066449f
C4899 VSSD.t807 VSUBS 0.100597f
C4900 VSSD.t924 VSUBS 0.143974f
C4901 VSSD.t912 VSUBS 0.097828f
C4902 VSSD.t865 VSUBS 0.097828f
C4903 VSSD.t324 VSUBS 0.128284f
C4904 VSSD.t1083 VSUBS 0.087676f
C4905 VSSD.t11 VSUBS 0.083985f
C4906 VSSD.t415 VSUBS 0.227958f
C4907 VSSD.t914 VSUBS 0.199348f
C4908 VSSD.t326 VSUBS 0.077524f
C4909 VSSD.t910 VSUBS 0.077524f
C4910 VSSD.t878 VSUBS 0.067372f
C4911 VSSD.n2013 VSUBS 0.866992f
C4912 VSSD.t1162 VSUBS 0.226378f
C4913 VSSD.t375 VSUBS 0.633857f
C4914 VSSD.t184 VSUBS 0.633857f
C4915 VSSD.t372 VSUBS 0.799867f
C4916 VSSD.t377 VSUBS 1.26771f
C4917 VSSD.t546 VSUBS 0.769684f
C4918 VSSD.t381 VSUBS 0.633857f
C4919 VSSD.t851 VSUBS 0.686678f
C4920 VSSD.t944 VSUBS 0.633857f
C4921 VSSD.t548 VSUBS 1.07907f
C4922 VSSD.t857 VSUBS 0.679133f
C4923 VSSD.t1164 VSUBS 0.633857f
C4924 VSSD.t853 VSUBS 0.724408f
C4925 VSSD.t930 VSUBS 0.633857f
C4926 VSSD.t1190 VSUBS 0.822505f
C4927 VSSD.t379 VSUBS 0.633857f
C4928 VSSD.t859 VSUBS 0.747046f
C4929 VSSD.t458 VSUBS 0.633857f
C4930 VSSD.t855 VSUBS 0.996061f
C4931 VSSD.t1124 VSUBS 1.34317f
C4932 VSSD.t550 VSUBS 0.769684f
C4933 VSSD.n2014 VSUBS 7.95717f
C4934 VSSD.t916 VSUBS 4.87295f
C4935 VSSD.t398 VSUBS 4.01178f
C4936 VSSD.t612 VSUBS 7.35143f
C4937 VSSD.t985 VSUBS 7.12039f
C4938 VSSD.t820 VSUBS 3.12961f
C4939 VSSD.n2015 VSUBS 0.47246p
C4940 VSSD.n2016 VSUBS 0.242461p
C4941 VSSD.n2017 VSUBS 0.099854f
C4942 VSSD.n2018 VSUBS -0.034903f
C4943 CLKS.n0 VSUBS 0.010823f
C4944 CLKS.t122 VSUBS 0.033285f
C4945 CLKS.t82 VSUBS 0.020962f
C4946 CLKS.n1 VSUBS 0.064926f
C4947 CLKS.n2 VSUBS 0.01402f
C4948 CLKS.n3 VSUBS 0.020787f
C4949 CLKS.n4 VSUBS 0.032671f
C4950 CLKS.t138 VSUBS 0.038238f
C4951 CLKS.t71 VSUBS 0.016321f
C4952 CLKS.n5 VSUBS 0.067818f
C4953 CLKS.n6 VSUBS 0.076076f
C4954 CLKS.n7 VSUBS 0.093952f
C4955 CLKS.n8 VSUBS 0.238627f
C4956 CLKS.n9 VSUBS 0.045213f
C4957 CLKS.n10 VSUBS 0.010222f
C4958 CLKS.n11 VSUBS 0.010759f
C4959 CLKS.t128 VSUBS 0.020962f
C4960 CLKS.t131 VSUBS 0.033285f
C4961 CLKS.n12 VSUBS 0.064926f
C4962 CLKS.n13 VSUBS 0.01402f
C4963 CLKS.n14 VSUBS 0.030148f
C4964 CLKS.n15 VSUBS 0.010627f
C4965 CLKS.t111 VSUBS 0.016321f
C4966 CLKS.t52 VSUBS 0.038238f
C4967 CLKS.n16 VSUBS 0.067818f
C4968 CLKS.n17 VSUBS 0.076076f
C4969 CLKS.n18 VSUBS 0.093952f
C4970 CLKS.n19 VSUBS 0.238627f
C4971 CLKS.n20 VSUBS 0.032806f
C4972 CLKS.n21 VSUBS 0.41793f
C4973 CLKS.n22 VSUBS 0.010823f
C4974 CLKS.t110 VSUBS 0.033285f
C4975 CLKS.t75 VSUBS 0.020962f
C4976 CLKS.n23 VSUBS 0.064926f
C4977 CLKS.n24 VSUBS 0.01402f
C4978 CLKS.n25 VSUBS 0.020787f
C4979 CLKS.n26 VSUBS 0.032671f
C4980 CLKS.t40 VSUBS 0.038238f
C4981 CLKS.t65 VSUBS 0.016321f
C4982 CLKS.n27 VSUBS 0.067818f
C4983 CLKS.n28 VSUBS 0.076076f
C4984 CLKS.n29 VSUBS 0.093952f
C4985 CLKS.n30 VSUBS 0.238627f
C4986 CLKS.n31 VSUBS 0.045213f
C4987 CLKS.n32 VSUBS 0.010222f
C4988 CLKS.n33 VSUBS 0.010759f
C4989 CLKS.t115 VSUBS 0.020962f
C4990 CLKS.t58 VSUBS 0.033285f
C4991 CLKS.n34 VSUBS 0.064926f
C4992 CLKS.n35 VSUBS 0.01402f
C4993 CLKS.n36 VSUBS 0.030148f
C4994 CLKS.n37 VSUBS 0.010627f
C4995 CLKS.t104 VSUBS 0.016321f
C4996 CLKS.t62 VSUBS 0.038238f
C4997 CLKS.n38 VSUBS 0.067818f
C4998 CLKS.n39 VSUBS 0.076076f
C4999 CLKS.n40 VSUBS 0.093952f
C5000 CLKS.n41 VSUBS 0.238627f
C5001 CLKS.n42 VSUBS 0.032806f
C5002 CLKS.n43 VSUBS 0.237802f
C5003 CLKS.n44 VSUBS 1.91503f
C5004 CLKS.n45 VSUBS 0.010823f
C5005 CLKS.t29 VSUBS 0.033285f
C5006 CLKS.t109 VSUBS 0.020962f
C5007 CLKS.n46 VSUBS 0.064926f
C5008 CLKS.n47 VSUBS 0.01402f
C5009 CLKS.n48 VSUBS 0.020787f
C5010 CLKS.n49 VSUBS 0.032671f
C5011 CLKS.t57 VSUBS 0.038238f
C5012 CLKS.t85 VSUBS 0.016321f
C5013 CLKS.n50 VSUBS 0.067818f
C5014 CLKS.n51 VSUBS 0.076076f
C5015 CLKS.n52 VSUBS 0.093952f
C5016 CLKS.n53 VSUBS 0.238627f
C5017 CLKS.n54 VSUBS 0.045226f
C5018 CLKS.n55 VSUBS 0.010222f
C5019 CLKS.n56 VSUBS 0.010759f
C5020 CLKS.t31 VSUBS 0.020962f
C5021 CLKS.t94 VSUBS 0.033285f
C5022 CLKS.n57 VSUBS 0.064926f
C5023 CLKS.n58 VSUBS 0.01402f
C5024 CLKS.n59 VSUBS 0.030148f
C5025 CLKS.n60 VSUBS 0.010627f
C5026 CLKS.t134 VSUBS 0.016321f
C5027 CLKS.t39 VSUBS 0.038238f
C5028 CLKS.n61 VSUBS 0.067818f
C5029 CLKS.n62 VSUBS 0.076076f
C5030 CLKS.n63 VSUBS 0.093952f
C5031 CLKS.n64 VSUBS 0.238627f
C5032 CLKS.n65 VSUBS 0.03286f
C5033 CLKS.n66 VSUBS 0.235973f
C5034 CLKS.n67 VSUBS 1.37057f
C5035 CLKS.n68 VSUBS 0.010823f
C5036 CLKS.t86 VSUBS 0.033285f
C5037 CLKS.t55 VSUBS 0.020962f
C5038 CLKS.n69 VSUBS 0.064926f
C5039 CLKS.n70 VSUBS 0.01402f
C5040 CLKS.n71 VSUBS 0.020787f
C5041 CLKS.n72 VSUBS 0.032671f
C5042 CLKS.t88 VSUBS 0.038238f
C5043 CLKS.t126 VSUBS 0.016321f
C5044 CLKS.n73 VSUBS 0.067818f
C5045 CLKS.n74 VSUBS 0.076076f
C5046 CLKS.n75 VSUBS 0.093952f
C5047 CLKS.n76 VSUBS 0.238627f
C5048 CLKS.n77 VSUBS 0.045226f
C5049 CLKS.n78 VSUBS 0.010222f
C5050 CLKS.n79 VSUBS 0.010759f
C5051 CLKS.t89 VSUBS 0.020962f
C5052 CLKS.t93 VSUBS 0.033285f
C5053 CLKS.n80 VSUBS 0.064926f
C5054 CLKS.n81 VSUBS 0.01402f
C5055 CLKS.n82 VSUBS 0.030148f
C5056 CLKS.n83 VSUBS 0.010627f
C5057 CLKS.t43 VSUBS 0.016321f
C5058 CLKS.t74 VSUBS 0.038238f
C5059 CLKS.n84 VSUBS 0.067818f
C5060 CLKS.n85 VSUBS 0.076076f
C5061 CLKS.n86 VSUBS 0.093952f
C5062 CLKS.n87 VSUBS 0.238627f
C5063 CLKS.n88 VSUBS 0.03286f
C5064 CLKS.n89 VSUBS 0.235973f
C5065 CLKS.n90 VSUBS 1.37061f
C5066 CLKS.n91 VSUBS 0.010823f
C5067 CLKS.t81 VSUBS 0.033285f
C5068 CLKS.t49 VSUBS 0.020962f
C5069 CLKS.n92 VSUBS 0.064926f
C5070 CLKS.n93 VSUBS 0.01402f
C5071 CLKS.n94 VSUBS 0.020787f
C5072 CLKS.n95 VSUBS 0.032671f
C5073 CLKS.t132 VSUBS 0.038238f
C5074 CLKS.t114 VSUBS 0.016321f
C5075 CLKS.n96 VSUBS 0.067818f
C5076 CLKS.n97 VSUBS 0.076076f
C5077 CLKS.n98 VSUBS 0.093952f
C5078 CLKS.n99 VSUBS 0.238627f
C5079 CLKS.n100 VSUBS 0.045226f
C5080 CLKS.n101 VSUBS 0.010222f
C5081 CLKS.n102 VSUBS 0.010759f
C5082 CLKS.t84 VSUBS 0.020962f
C5083 CLKS.t33 VSUBS 0.033285f
C5084 CLKS.n103 VSUBS 0.064926f
C5085 CLKS.n104 VSUBS 0.01402f
C5086 CLKS.n105 VSUBS 0.030148f
C5087 CLKS.n106 VSUBS 0.010627f
C5088 CLKS.t36 VSUBS 0.016321f
C5089 CLKS.t117 VSUBS 0.038238f
C5090 CLKS.n107 VSUBS 0.067818f
C5091 CLKS.n108 VSUBS 0.076076f
C5092 CLKS.n109 VSUBS 0.093952f
C5093 CLKS.n110 VSUBS 0.238627f
C5094 CLKS.n111 VSUBS 0.03286f
C5095 CLKS.n112 VSUBS 0.235973f
C5096 CLKS.n113 VSUBS 1.37061f
C5097 CLKS.n114 VSUBS 0.010823f
C5098 CLKS.t137 VSUBS 0.033285f
C5099 CLKS.t95 VSUBS 0.020962f
C5100 CLKS.n115 VSUBS 0.064926f
C5101 CLKS.n116 VSUBS 0.01402f
C5102 CLKS.n117 VSUBS 0.020787f
C5103 CLKS.n118 VSUBS 0.032671f
C5104 CLKS.t136 VSUBS 0.038238f
C5105 CLKS.t127 VSUBS 0.016321f
C5106 CLKS.n119 VSUBS 0.067818f
C5107 CLKS.n120 VSUBS 0.076076f
C5108 CLKS.n121 VSUBS 0.093952f
C5109 CLKS.n122 VSUBS 0.238627f
C5110 CLKS.n123 VSUBS 0.045226f
C5111 CLKS.n124 VSUBS 0.010222f
C5112 CLKS.n125 VSUBS 0.010759f
C5113 CLKS.t141 VSUBS 0.020962f
C5114 CLKS.t123 VSUBS 0.033285f
C5115 CLKS.n126 VSUBS 0.064926f
C5116 CLKS.n127 VSUBS 0.01402f
C5117 CLKS.n128 VSUBS 0.030148f
C5118 CLKS.n129 VSUBS 0.010627f
C5119 CLKS.t44 VSUBS 0.016321f
C5120 CLKS.t22 VSUBS 0.038238f
C5121 CLKS.n130 VSUBS 0.067818f
C5122 CLKS.n131 VSUBS 0.076076f
C5123 CLKS.n132 VSUBS 0.093952f
C5124 CLKS.n133 VSUBS 0.238627f
C5125 CLKS.n134 VSUBS 0.03286f
C5126 CLKS.n135 VSUBS 0.235973f
C5127 CLKS.n136 VSUBS 1.37061f
C5128 CLKS.n137 VSUBS 0.010823f
C5129 CLKS.t108 VSUBS 0.033285f
C5130 CLKS.t72 VSUBS 0.020962f
C5131 CLKS.n138 VSUBS 0.064926f
C5132 CLKS.n139 VSUBS 0.01402f
C5133 CLKS.n140 VSUBS 0.020787f
C5134 CLKS.n141 VSUBS 0.032671f
C5135 CLKS.t78 VSUBS 0.038238f
C5136 CLKS.t96 VSUBS 0.016321f
C5137 CLKS.n142 VSUBS 0.067818f
C5138 CLKS.n143 VSUBS 0.076076f
C5139 CLKS.n144 VSUBS 0.093952f
C5140 CLKS.n145 VSUBS 0.238627f
C5141 CLKS.n146 VSUBS 0.045226f
C5142 CLKS.n147 VSUBS 0.010222f
C5143 CLKS.n148 VSUBS 0.010759f
C5144 CLKS.t112 VSUBS 0.020962f
C5145 CLKS.t76 VSUBS 0.033285f
C5146 CLKS.n149 VSUBS 0.064926f
C5147 CLKS.n150 VSUBS 0.01402f
C5148 CLKS.n151 VSUBS 0.030148f
C5149 CLKS.n152 VSUBS 0.010627f
C5150 CLKS.t16 VSUBS 0.016321f
C5151 CLKS.t18 VSUBS 0.038238f
C5152 CLKS.n153 VSUBS 0.067818f
C5153 CLKS.n154 VSUBS 0.076076f
C5154 CLKS.n155 VSUBS 0.093952f
C5155 CLKS.n156 VSUBS 0.238627f
C5156 CLKS.n157 VSUBS 0.03286f
C5157 CLKS.n158 VSUBS 0.235973f
C5158 CLKS.n159 VSUBS 1.37061f
C5159 CLKS.n160 VSUBS 0.010823f
C5160 CLKS.t119 VSUBS 0.033285f
C5161 CLKS.t80 VSUBS 0.020962f
C5162 CLKS.n161 VSUBS 0.064926f
C5163 CLKS.n162 VSUBS 0.01402f
C5164 CLKS.n163 VSUBS 0.020787f
C5165 CLKS.n164 VSUBS 0.032671f
C5166 CLKS.t46 VSUBS 0.038238f
C5167 CLKS.t103 VSUBS 0.016321f
C5168 CLKS.n165 VSUBS 0.067818f
C5169 CLKS.n166 VSUBS 0.076076f
C5170 CLKS.n167 VSUBS 0.093952f
C5171 CLKS.n168 VSUBS 0.238627f
C5172 CLKS.n169 VSUBS 0.045226f
C5173 CLKS.n170 VSUBS 0.010222f
C5174 CLKS.n171 VSUBS 0.010759f
C5175 CLKS.t124 VSUBS 0.020962f
C5176 CLKS.t26 VSUBS 0.033285f
C5177 CLKS.n172 VSUBS 0.064926f
C5178 CLKS.n173 VSUBS 0.01402f
C5179 CLKS.n174 VSUBS 0.030148f
C5180 CLKS.n175 VSUBS 0.010627f
C5181 CLKS.t25 VSUBS 0.016321f
C5182 CLKS.t97 VSUBS 0.038238f
C5183 CLKS.n176 VSUBS 0.067818f
C5184 CLKS.n177 VSUBS 0.076076f
C5185 CLKS.n178 VSUBS 0.093952f
C5186 CLKS.n179 VSUBS 0.238627f
C5187 CLKS.n180 VSUBS 0.03286f
C5188 CLKS.n181 VSUBS 0.235973f
C5189 CLKS.n182 VSUBS 1.37061f
C5190 CLKS.n183 VSUBS 0.010823f
C5191 CLKS.t64 VSUBS 0.033285f
C5192 CLKS.t35 VSUBS 0.020962f
C5193 CLKS.n184 VSUBS 0.064926f
C5194 CLKS.n185 VSUBS 0.01402f
C5195 CLKS.n186 VSUBS 0.020787f
C5196 CLKS.n187 VSUBS 0.032671f
C5197 CLKS.t51 VSUBS 0.038238f
C5198 CLKS.t69 VSUBS 0.016321f
C5199 CLKS.n188 VSUBS 0.067818f
C5200 CLKS.n189 VSUBS 0.076076f
C5201 CLKS.n190 VSUBS 0.093952f
C5202 CLKS.n191 VSUBS 0.238627f
C5203 CLKS.n192 VSUBS 0.045226f
C5204 CLKS.n193 VSUBS 0.010222f
C5205 CLKS.n194 VSUBS 0.010759f
C5206 CLKS.t67 VSUBS 0.020962f
C5207 CLKS.t90 VSUBS 0.033285f
C5208 CLKS.n195 VSUBS 0.064926f
C5209 CLKS.n196 VSUBS 0.01402f
C5210 CLKS.n197 VSUBS 0.030148f
C5211 CLKS.n198 VSUBS 0.010627f
C5212 CLKS.t107 VSUBS 0.016321f
C5213 CLKS.t47 VSUBS 0.038238f
C5214 CLKS.n199 VSUBS 0.067818f
C5215 CLKS.n200 VSUBS 0.076076f
C5216 CLKS.n201 VSUBS 0.093952f
C5217 CLKS.n202 VSUBS 0.238627f
C5218 CLKS.n203 VSUBS 0.03286f
C5219 CLKS.n204 VSUBS 0.235973f
C5220 CLKS.n205 VSUBS 1.37061f
C5221 CLKS.n206 VSUBS 0.010823f
C5222 CLKS.t37 VSUBS 0.033285f
C5223 CLKS.t121 VSUBS 0.020962f
C5224 CLKS.n207 VSUBS 0.064926f
C5225 CLKS.n208 VSUBS 0.01402f
C5226 CLKS.n209 VSUBS 0.020787f
C5227 CLKS.n210 VSUBS 0.032671f
C5228 CLKS.t19 VSUBS 0.038238f
C5229 CLKS.t41 VSUBS 0.016321f
C5230 CLKS.n211 VSUBS 0.067818f
C5231 CLKS.n212 VSUBS 0.076076f
C5232 CLKS.n213 VSUBS 0.093952f
C5233 CLKS.n214 VSUBS 0.238627f
C5234 CLKS.n215 VSUBS 0.045226f
C5235 CLKS.n216 VSUBS 0.010222f
C5236 CLKS.n217 VSUBS 0.010759f
C5237 CLKS.t38 VSUBS 0.020962f
C5238 CLKS.t56 VSUBS 0.033285f
C5239 CLKS.n218 VSUBS 0.064926f
C5240 CLKS.n219 VSUBS 0.01402f
C5241 CLKS.n220 VSUBS 0.030148f
C5242 CLKS.n221 VSUBS 0.010627f
C5243 CLKS.t73 VSUBS 0.016321f
C5244 CLKS.t135 VSUBS 0.038238f
C5245 CLKS.n222 VSUBS 0.067818f
C5246 CLKS.n223 VSUBS 0.076076f
C5247 CLKS.n224 VSUBS 0.093952f
C5248 CLKS.n225 VSUBS 0.238627f
C5249 CLKS.n226 VSUBS 0.03286f
C5250 CLKS.n227 VSUBS 0.235973f
C5251 CLKS.n228 VSUBS 1.70531f
C5252 CLKS.t63 VSUBS 0.039413f
C5253 CLKS.t130 VSUBS 0.024614f
C5254 CLKS.n229 VSUBS 0.073973f
C5255 CLKS.n230 VSUBS 0.021723f
C5256 CLKS.t14 VSUBS 0.023792f
C5257 CLKS.t9 VSUBS 0.023792f
C5258 CLKS.n231 VSUBS 0.052889f
C5259 CLKS.n232 VSUBS 0.147908f
C5260 CLKS.t1 VSUBS 0.015465f
C5261 CLKS.t4 VSUBS 0.015465f
C5262 CLKS.n233 VSUBS 0.035221f
C5263 CLKS.t13 VSUBS 0.015465f
C5264 CLKS.t0 VSUBS 0.015465f
C5265 CLKS.n234 VSUBS 0.035221f
C5266 CLKS.t15 VSUBS 0.015465f
C5267 CLKS.t6 VSUBS 0.015465f
C5268 CLKS.n235 VSUBS 0.035221f
C5269 CLKS.t8 VSUBS 0.015465f
C5270 CLKS.t3 VSUBS 0.015465f
C5271 CLKS.n236 VSUBS 0.035221f
C5272 CLKS.t5 VSUBS 0.023792f
C5273 CLKS.t7 VSUBS 0.023792f
C5274 CLKS.n237 VSUBS 0.052889f
C5275 CLKS.t11 VSUBS 0.023792f
C5276 CLKS.t10 VSUBS 0.023792f
C5277 CLKS.n238 VSUBS 0.052889f
C5278 CLKS.t2 VSUBS 0.023792f
C5279 CLKS.t12 VSUBS 0.023792f
C5280 CLKS.n239 VSUBS 0.052889f
C5281 CLKS.n240 VSUBS 0.138083f
C5282 CLKS.n241 VSUBS 0.138083f
C5283 CLKS.n242 VSUBS 0.152876f
C5284 CLKS.n243 VSUBS 0.111675f
C5285 CLKS.n244 VSUBS 0.10547f
C5286 CLKS.n245 VSUBS 0.10547f
C5287 CLKS.n246 VSUBS 0.111023f
C5288 CLKS.n247 VSUBS 0.04555f
C5289 CLKS.n248 VSUBS 0.147446f
C5290 CLKS.n249 VSUBS 6.39492f
C5291 CLKS.t101 VSUBS 0.016321f
C5292 CLKS.t98 VSUBS 0.038238f
C5293 CLKS.n250 VSUBS 0.067899f
C5294 CLKS.n251 VSUBS 0.092719f
C5295 CLKS.n252 VSUBS 0.029282f
C5296 CLKS.t50 VSUBS 0.020962f
C5297 CLKS.t100 VSUBS 0.033285f
C5298 CLKS.n253 VSUBS 0.064926f
C5299 CLKS.n254 VSUBS 0.034408f
C5300 CLKS.n255 VSUBS 0.014012f
C5301 CLKS.n257 VSUBS 0.808301f
C5302 CLKS.t129 VSUBS 0.016321f
C5303 CLKS.t125 VSUBS 0.038238f
C5304 CLKS.n258 VSUBS 0.067899f
C5305 CLKS.n259 VSUBS 0.092719f
C5306 CLKS.n260 VSUBS 0.029282f
C5307 CLKS.t83 VSUBS 0.020962f
C5308 CLKS.t140 VSUBS 0.033285f
C5309 CLKS.n261 VSUBS 0.064926f
C5310 CLKS.n262 VSUBS 0.034408f
C5311 CLKS.n263 VSUBS 0.014012f
C5312 CLKS.n265 VSUBS 0.876118f
C5313 CLKS.t118 VSUBS 0.016321f
C5314 CLKS.t113 VSUBS 0.038238f
C5315 CLKS.n266 VSUBS 0.067899f
C5316 CLKS.n267 VSUBS 0.092719f
C5317 CLKS.n268 VSUBS 0.029282f
C5318 CLKS.t105 VSUBS 0.020962f
C5319 CLKS.t42 VSUBS 0.033285f
C5320 CLKS.n269 VSUBS 0.064926f
C5321 CLKS.n270 VSUBS 0.034408f
C5322 CLKS.n271 VSUBS 0.014012f
C5323 CLKS.n273 VSUBS 0.876118f
C5324 CLKS.t34 VSUBS 0.016321f
C5325 CLKS.t30 VSUBS 0.038238f
C5326 CLKS.n274 VSUBS 0.067899f
C5327 CLKS.n275 VSUBS 0.092719f
C5328 CLKS.n276 VSUBS 0.029282f
C5329 CLKS.t24 VSUBS 0.020962f
C5330 CLKS.t70 VSUBS 0.033285f
C5331 CLKS.n277 VSUBS 0.064926f
C5332 CLKS.n278 VSUBS 0.034408f
C5333 CLKS.n279 VSUBS 0.014012f
C5334 CLKS.n281 VSUBS 0.863268f
C5335 CLKS.t91 VSUBS 0.016321f
C5336 CLKS.t87 VSUBS 0.038238f
C5337 CLKS.n282 VSUBS 0.067899f
C5338 CLKS.n283 VSUBS 0.092719f
C5339 CLKS.n284 VSUBS 0.029282f
C5340 CLKS.t60 VSUBS 0.020962f
C5341 CLKS.t116 VSUBS 0.033285f
C5342 CLKS.n285 VSUBS 0.064926f
C5343 CLKS.n286 VSUBS 0.034408f
C5344 CLKS.n287 VSUBS 0.014012f
C5345 CLKS.n289 VSUBS 0.533763f
C5346 CLKS.n290 VSUBS 0.020694f
C5347 CLKS.t53 VSUBS 0.038238f
C5348 CLKS.t45 VSUBS 0.016321f
C5349 CLKS.n291 VSUBS 0.067818f
C5350 CLKS.n292 VSUBS 0.076076f
C5351 CLKS.n293 VSUBS 0.095185f
C5352 CLKS.t27 VSUBS 0.033285f
C5353 CLKS.t54 VSUBS 0.020962f
C5354 CLKS.n294 VSUBS 0.064926f
C5355 CLKS.n295 VSUBS 0.01402f
C5356 CLKS.n296 VSUBS 0.010759f
C5357 CLKS.n297 VSUBS 0.02555f
C5358 CLKS.n298 VSUBS 0.027322f
C5359 CLKS.n299 VSUBS 0.249115f
C5360 CLKS.n300 VSUBS 0.020694f
C5361 CLKS.t61 VSUBS 0.038238f
C5362 CLKS.t77 VSUBS 0.016321f
C5363 CLKS.n301 VSUBS 0.067818f
C5364 CLKS.n302 VSUBS 0.076076f
C5365 CLKS.n303 VSUBS 0.095185f
C5366 CLKS.t92 VSUBS 0.033285f
C5367 CLKS.t48 VSUBS 0.020962f
C5368 CLKS.n304 VSUBS 0.064926f
C5369 CLKS.n305 VSUBS 0.01402f
C5370 CLKS.n306 VSUBS 0.010759f
C5371 CLKS.n307 VSUBS 0.02555f
C5372 CLKS.n308 VSUBS 0.027322f
C5373 CLKS.n309 VSUBS 0.022907f
C5374 CLKS.n310 VSUBS 1.0953f
C5375 CLKS.n311 VSUBS 0.020694f
C5376 CLKS.t17 VSUBS 0.038238f
C5377 CLKS.t68 VSUBS 0.016321f
C5378 CLKS.n312 VSUBS 0.067818f
C5379 CLKS.n313 VSUBS 0.076076f
C5380 CLKS.n314 VSUBS 0.095185f
C5381 CLKS.t21 VSUBS 0.033285f
C5382 CLKS.t79 VSUBS 0.020962f
C5383 CLKS.n315 VSUBS 0.064926f
C5384 CLKS.n316 VSUBS 0.01402f
C5385 CLKS.n317 VSUBS 0.010759f
C5386 CLKS.n318 VSUBS 0.02555f
C5387 CLKS.n319 VSUBS 0.027322f
C5388 CLKS.n320 VSUBS 0.022907f
C5389 CLKS.n321 VSUBS 0.876118f
C5390 CLKS.n322 VSUBS 0.020694f
C5391 CLKS.t59 VSUBS 0.038238f
C5392 CLKS.t102 VSUBS 0.016321f
C5393 CLKS.n323 VSUBS 0.067818f
C5394 CLKS.n324 VSUBS 0.076076f
C5395 CLKS.n325 VSUBS 0.095185f
C5396 CLKS.t32 VSUBS 0.033285f
C5397 CLKS.t28 VSUBS 0.020962f
C5398 CLKS.n326 VSUBS 0.064926f
C5399 CLKS.n327 VSUBS 0.01402f
C5400 CLKS.n328 VSUBS 0.010759f
C5401 CLKS.n329 VSUBS 0.02555f
C5402 CLKS.n330 VSUBS 0.027322f
C5403 CLKS.n331 VSUBS 0.022907f
C5404 CLKS.n332 VSUBS 0.876118f
C5405 CLKS.n333 VSUBS 0.020694f
C5406 CLKS.t23 VSUBS 0.038238f
C5407 CLKS.t133 VSUBS 0.016321f
C5408 CLKS.n334 VSUBS 0.067818f
C5409 CLKS.n335 VSUBS 0.076076f
C5410 CLKS.n336 VSUBS 0.095185f
C5411 CLKS.t99 VSUBS 0.033285f
C5412 CLKS.t20 VSUBS 0.020962f
C5413 CLKS.n337 VSUBS 0.064926f
C5414 CLKS.n338 VSUBS 0.01402f
C5415 CLKS.n339 VSUBS 0.010759f
C5416 CLKS.n340 VSUBS 0.02555f
C5417 CLKS.n341 VSUBS 0.027322f
C5418 CLKS.n342 VSUBS 0.022907f
C5419 CLKS.n343 VSUBS 0.664878f
C5420 CLKS.n344 VSUBS 0.437142f
C5421 CLKS.n345 VSUBS 7.10874f
C5422 CLKS.t66 VSUBS 0.018228f
C5423 CLKS.t106 VSUBS 0.026476f
C5424 CLKS.n346 VSUBS 0.063031f
C5425 CLKS.n347 VSUBS 0.046689f
C5426 CLKS.t139 VSUBS 0.026476f
C5427 CLKS.t120 VSUBS 0.018228f
C5428 CLKS.n348 VSUBS 0.062943f
C5429 CLKS.n349 VSUBS 0.026916f
C5430 CLKS.n350 VSUBS 0.439118f
C5431 CLKS.n351 VSUBS 10.450299f
C5432 VDDD.n0 VSUBS 1.48589f
C5433 VDDD.n1 VSUBS 10.4828f
C5434 VDDD.t1007 VSUBS 1.66443f
C5435 VDDD.t117 VSUBS 1.3672f
C5436 VDDD.t691 VSUBS 1.3672f
C5437 VDDD.t463 VSUBS 0.877942f
C5438 VDDD.t1009 VSUBS 0.877942f
C5439 VDDD.t234 VSUBS 0.777344f
C5440 VDDD.t950 VSUBS 0.845919f
C5441 VDDD.t1107 VSUBS 1.35346f
C5442 VDDD.t905 VSUBS 1.34432f
C5443 VDDD.t1355 VSUBS 1.08369f
C5444 VDDD.t947 VSUBS 1.09284f
C5445 VDDD.t374 VSUBS 0.873355f
C5446 VDDD.t1037 VSUBS 1.64155f
C5447 VDDD.t948 VSUBS 1.60497f
C5448 VDDD.t282 VSUBS 0.681305f
C5449 VDDD.t334 VSUBS 0.983097f
C5450 VDDD.t1386 VSUBS 1.3672f
C5451 VDDD.t731 VSUBS 1.3672f
C5452 VDDD.t502 VSUBS 0.877942f
C5453 VDDD.t336 VSUBS 0.877942f
C5454 VDDD.t519 VSUBS 0.777344f
C5455 VDDD.t1176 VSUBS 0.845919f
C5456 VDDD.t1195 VSUBS 1.35346f
C5457 VDDD.t1304 VSUBS 1.34432f
C5458 VDDD.t605 VSUBS 1.08369f
C5459 VDDD.t1173 VSUBS 1.09284f
C5460 VDDD.t933 VSUBS 0.873355f
C5461 VDDD.t705 VSUBS 1.64155f
C5462 VDDD.t1174 VSUBS 1.60497f
C5463 VDDD.t917 VSUBS 0.681305f
C5464 VDDD.t713 VSUBS 0.983097f
C5465 VDDD.t715 VSUBS 1.3672f
C5466 VDDD.t580 VSUBS 1.3672f
C5467 VDDD.t261 VSUBS 0.877942f
C5468 VDDD.t711 VSUBS 0.877942f
C5469 VDDD.t1190 VSUBS 0.777344f
C5470 VDDD.t497 VSUBS 0.845919f
C5471 VDDD.t332 VSUBS 1.35346f
C5472 VDDD.t613 VSUBS 1.34432f
C5473 VDDD.t808 VSUBS 1.08369f
C5474 VDDD.t273 VSUBS 1.09284f
C5475 VDDD.t1189 VSUBS 0.873355f
C5476 VDDD.t1120 VSUBS 1.64155f
C5477 VDDD.t274 VSUBS 1.60497f
C5478 VDDD.t241 VSUBS 0.681305f
C5479 VDDD.t80 VSUBS 0.983097f
C5480 VDDD.t770 VSUBS 1.3672f
C5481 VDDD.t603 VSUBS 1.3672f
C5482 VDDD.t851 VSUBS 0.877942f
C5483 VDDD.t725 VSUBS 0.877942f
C5484 VDDD.t735 VSUBS 0.777344f
C5485 VDDD.t1150 VSUBS 0.845919f
C5486 VDDD.t193 VSUBS 1.35346f
C5487 VDDD.t1312 VSUBS 1.34432f
C5488 VDDD.t999 VSUBS 1.08369f
C5489 VDDD.t1151 VSUBS 1.09284f
C5490 VDDD.t524 VSUBS 0.873355f
C5491 VDDD.t707 VSUBS 1.64155f
C5492 VDDD.t1001 VSUBS 1.60497f
C5493 VDDD.t717 VSUBS 0.681305f
C5494 VDDD.t1035 VSUBS 0.983097f
C5495 VDDD.t1031 VSUBS 1.3672f
C5496 VDDD.t63 VSUBS 1.3672f
C5497 VDDD.t1274 VSUBS 0.877942f
C5498 VDDD.t1033 VSUBS 0.877942f
C5499 VDDD.t801 VSUBS 0.777344f
C5500 VDDD.t751 VSUBS 0.845919f
C5501 VDDD.t594 VSUBS 1.35346f
C5502 VDDD.t171 VSUBS 1.34432f
C5503 VDDD.t141 VSUBS 1.08369f
C5504 VDDD.t750 VSUBS 1.09284f
C5505 VDDD.t564 VSUBS 0.873355f
C5506 VDDD.t1122 VSUBS 1.64155f
C5507 VDDD.t752 VSUBS 1.60497f
C5508 VDDD.t535 VSUBS 0.681305f
C5509 VDDD.t183 VSUBS 0.983097f
C5510 VDDD.t146 VSUBS 1.3672f
C5511 VDDD.t301 VSUBS 1.3672f
C5512 VDDD.t490 VSUBS 0.877942f
C5513 VDDD.t370 VSUBS 0.877942f
C5514 VDDD.t741 VSUBS 0.777344f
C5515 VDDD.t310 VSUBS 0.845919f
C5516 VDDD.t587 VSUBS 1.35346f
C5517 VDDD.t634 VSUBS 1.34432f
C5518 VDDD.t298 VSUBS 1.08369f
C5519 VDDD.t307 VSUBS 1.09284f
C5520 VDDD.t742 VSUBS 0.873355f
C5521 VDDD.t1118 VSUBS 1.64155f
C5522 VDDD.t308 VSUBS 1.60497f
C5523 VDDD.t4 VSUBS 0.681305f
C5524 VDDD.t1357 VSUBS 0.983097f
C5525 VDDD.t1361 VSUBS 1.3672f
C5526 VDDD.t736 VSUBS 1.3672f
C5527 VDDD.t1314 VSUBS 0.877942f
C5528 VDDD.t1359 VSUBS 0.877942f
C5529 VDDD.t379 VSUBS 0.777344f
C5530 VDDD.t590 VSUBS 0.845919f
C5531 VDDD.t27 VSUBS 1.35346f
C5532 VDDD.t546 VSUBS 1.34432f
C5533 VDDD.t745 VSUBS 1.08369f
C5534 VDDD.t57 VSUBS 1.09284f
C5535 VDDD.t380 VSUBS 0.873355f
C5536 VDDD.t1039 VSUBS 1.64155f
C5537 VDDD.t591 VSUBS 1.60497f
C5538 VDDD.t1287 VSUBS 0.681305f
C5539 VDDD.t863 VSUBS 0.983097f
C5540 VDDD.t78 VSUBS 1.3672f
C5541 VDDD.t695 VSUBS 1.3672f
C5542 VDDD.t513 VSUBS 0.877942f
C5543 VDDD.t76 VSUBS 0.877942f
C5544 VDDD.t982 VSUBS 0.777344f
C5545 VDDD.t494 VSUBS 0.845919f
C5546 VDDD.t723 VSUBS 1.35346f
C5547 VDDD.t263 VSUBS 1.34432f
C5548 VDDD.t686 VSUBS 1.08369f
C5549 VDDD.t775 VSUBS 1.09284f
C5550 VDDD.t981 VSUBS 0.873355f
C5551 VDDD.t1185 VSUBS 1.64155f
C5552 VDDD.t773 VSUBS 1.60497f
C5553 VDDD.t853 VSUBS 0.681305f
C5554 VDDD.t319 VSUBS 0.983097f
C5555 VDDD.t317 VSUBS 1.3672f
C5556 VDDD.t1136 VSUBS 1.3672f
C5557 VDDD.t847 VSUBS 0.877942f
C5558 VDDD.t315 VSUBS 0.877942f
C5559 VDDD.t1168 VSUBS 0.777344f
C5560 VDDD.t638 VSUBS 0.845919f
C5561 VDDD.t1282 VSUBS 1.35346f
C5562 VDDD.t901 VSUBS 1.34432f
C5563 VDDD.t154 VSUBS 1.08369f
C5564 VDDD.t639 VSUBS 1.09284f
C5565 VDDD.t166 VSUBS 0.873355f
C5566 VDDD.t1041 VSUBS 1.64155f
C5567 VDDD.t6 VSUBS 1.60497f
C5568 VDDD.t1131 VSUBS 0.681305f
C5569 VDDD.t21 VSUBS 0.983097f
C5570 VDDD.t599 VSUBS 1.3672f
C5571 VDDD.t74 VSUBS 1.3672f
C5572 VDDD.t498 VSUBS 0.877942f
C5573 VDDD.t23 VSUBS 0.877942f
C5574 VDDD.t997 VSUBS 0.777344f
C5575 VDDD.t921 VSUBS 0.845919f
C5576 VDDD.t845 VSUBS 1.35346f
C5577 VDDD.t1213 VSUBS 1.34432f
C5578 VDDD.t355 VSUBS 1.08369f
C5579 VDDD.t1165 VSUBS 1.09284f
C5580 VDDD.t998 VSUBS 0.873355f
C5581 VDDD.t1183 VSUBS 1.64155f
C5582 VDDD.t922 VSUBS 1.60497f
C5583 VDDD.t977 VSUBS 0.681305f
C5584 VDDD.t384 VSUBS 1.29403f
C5585 VDDD.t399 VSUBS 0.768199f
C5586 VDDD.t401 VSUBS 0.768199f
C5587 VDDD.t386 VSUBS 0.768199f
C5588 VDDD.t390 VSUBS 0.768199f
C5589 VDDD.t1454 VSUBS 0.768199f
C5590 VDDD.t267 VSUBS 0.768199f
C5591 VDDD.t388 VSUBS 0.768199f
C5592 VDDD.t480 VSUBS 0.768199f
C5593 VDDD.t286 VSUBS 0.768199f
C5594 VDDD.t478 VSUBS 0.676747f
C5595 VDDD.n2 VSUBS 0.251622f
C5596 VDDD.t287 VSUBS 0.076922f
C5597 VDDD.t479 VSUBS 0.076922f
C5598 VDDD.n3 VSUBS 0.165125f
C5599 VDDD.t389 VSUBS 0.076922f
C5600 VDDD.t481 VSUBS 0.076922f
C5601 VDDD.n4 VSUBS 0.165125f
C5602 VDDD.n5 VSUBS 0.188262f
C5603 VDDD.n6 VSUBS 0.251622f
C5604 VDDD.n7 VSUBS 0.048917f
C5605 VDDD.n8 VSUBS 0.251622f
C5606 VDDD.t385 VSUBS 0.307526f
C5607 VDDD.n9 VSUBS 0.542325f
C5608 VDDD.t923 VSUBS 0.04923f
C5609 VDDD.t978 VSUBS 0.04923f
C5610 VDDD.n10 VSUBS 0.102503f
C5611 VDDD.n11 VSUBS 0.305072f
C5612 VDDD.n12 VSUBS 0.251622f
C5613 VDDD.n13 VSUBS 0.08621f
C5614 VDDD.t1184 VSUBS 0.118653f
C5615 VDDD.n14 VSUBS 0.251622f
C5616 VDDD.t1214 VSUBS 0.032307f
C5617 VDDD.t356 VSUBS 0.047863f
C5618 VDDD.n15 VSUBS 0.083298f
C5619 VDDD.n16 VSUBS 0.235104f
C5620 VDDD.n17 VSUBS 0.251622f
C5621 VDDD.n18 VSUBS 0.085726f
C5622 VDDD.t846 VSUBS 0.229702f
C5623 VDDD.n19 VSUBS 0.251622f
C5624 VDDD.n20 VSUBS 0.05037f
C5625 VDDD.t499 VSUBS 0.032307f
C5626 VDDD.t24 VSUBS 0.061025f
C5627 VDDD.n21 VSUBS 0.096588f
C5628 VDDD.n22 VSUBS 0.251622f
C5629 VDDD.t22 VSUBS 0.306728f
C5630 VDDD.n23 VSUBS 0.427682f
C5631 VDDD.n24 VSUBS 0.251622f
C5632 VDDD.n25 VSUBS 0.067806f
C5633 VDDD.n26 VSUBS 0.251622f
C5634 VDDD.n27 VSUBS 0.089116f
C5635 VDDD.n28 VSUBS 0.251622f
C5636 VDDD.t1283 VSUBS 0.229702f
C5637 VDDD.n29 VSUBS 0.3381f
C5638 VDDD.n30 VSUBS 0.251622f
C5639 VDDD.t848 VSUBS 0.032307f
C5640 VDDD.t316 VSUBS 0.061025f
C5641 VDDD.n31 VSUBS 0.096588f
C5642 VDDD.n32 VSUBS 0.24113f
C5643 VDDD.n33 VSUBS 0.251622f
C5644 VDDD.n34 VSUBS 0.057151f
C5645 VDDD.t318 VSUBS 0.337079f
C5646 VDDD.t774 VSUBS 0.04923f
C5647 VDDD.t854 VSUBS 0.04923f
C5648 VDDD.n35 VSUBS 0.102503f
C5649 VDDD.n36 VSUBS 0.305072f
C5650 VDDD.n37 VSUBS 0.251622f
C5651 VDDD.n38 VSUBS 0.08621f
C5652 VDDD.t1186 VSUBS 0.118653f
C5653 VDDD.n39 VSUBS 0.251622f
C5654 VDDD.t264 VSUBS 0.032307f
C5655 VDDD.t687 VSUBS 0.047863f
C5656 VDDD.n40 VSUBS 0.083298f
C5657 VDDD.n41 VSUBS 0.235104f
C5658 VDDD.n42 VSUBS 0.251622f
C5659 VDDD.n43 VSUBS 0.085726f
C5660 VDDD.t724 VSUBS 0.229702f
C5661 VDDD.n44 VSUBS 0.251622f
C5662 VDDD.n45 VSUBS 0.05037f
C5663 VDDD.t514 VSUBS 0.032307f
C5664 VDDD.t77 VSUBS 0.061025f
C5665 VDDD.n46 VSUBS 0.096588f
C5666 VDDD.n47 VSUBS 0.251622f
C5667 VDDD.t864 VSUBS 0.306728f
C5668 VDDD.n48 VSUBS 0.427682f
C5669 VDDD.n49 VSUBS 0.251622f
C5670 VDDD.n50 VSUBS 0.067806f
C5671 VDDD.n51 VSUBS 0.251622f
C5672 VDDD.n52 VSUBS 0.089116f
C5673 VDDD.n53 VSUBS 0.251622f
C5674 VDDD.t28 VSUBS 0.229702f
C5675 VDDD.n54 VSUBS 0.3381f
C5676 VDDD.n55 VSUBS 0.251622f
C5677 VDDD.t1315 VSUBS 0.032307f
C5678 VDDD.t1360 VSUBS 0.061025f
C5679 VDDD.n56 VSUBS 0.096588f
C5680 VDDD.n57 VSUBS 0.24113f
C5681 VDDD.n58 VSUBS 0.251622f
C5682 VDDD.n59 VSUBS 0.057151f
C5683 VDDD.t1362 VSUBS 0.337079f
C5684 VDDD.t309 VSUBS 0.04923f
C5685 VDDD.t5 VSUBS 0.04923f
C5686 VDDD.n60 VSUBS 0.102503f
C5687 VDDD.n61 VSUBS 0.305072f
C5688 VDDD.n62 VSUBS 0.251622f
C5689 VDDD.n63 VSUBS 0.08621f
C5690 VDDD.t1119 VSUBS 0.118653f
C5691 VDDD.n64 VSUBS 0.251622f
C5692 VDDD.t635 VSUBS 0.032307f
C5693 VDDD.t299 VSUBS 0.047863f
C5694 VDDD.n65 VSUBS 0.083298f
C5695 VDDD.n66 VSUBS 0.235104f
C5696 VDDD.n67 VSUBS 0.251622f
C5697 VDDD.n68 VSUBS 0.085726f
C5698 VDDD.t588 VSUBS 0.229702f
C5699 VDDD.n69 VSUBS 0.251622f
C5700 VDDD.n70 VSUBS 0.05037f
C5701 VDDD.t491 VSUBS 0.032307f
C5702 VDDD.t371 VSUBS 0.061025f
C5703 VDDD.n71 VSUBS 0.096588f
C5704 VDDD.n72 VSUBS 0.251622f
C5705 VDDD.t184 VSUBS 0.306728f
C5706 VDDD.n73 VSUBS 0.427682f
C5707 VDDD.n74 VSUBS 0.251622f
C5708 VDDD.n75 VSUBS 0.067806f
C5709 VDDD.n76 VSUBS 0.251622f
C5710 VDDD.n77 VSUBS 0.089116f
C5711 VDDD.n78 VSUBS 0.251622f
C5712 VDDD.t595 VSUBS 0.229702f
C5713 VDDD.n79 VSUBS 0.3381f
C5714 VDDD.n80 VSUBS 0.251622f
C5715 VDDD.t1275 VSUBS 0.032307f
C5716 VDDD.t1034 VSUBS 0.061025f
C5717 VDDD.n81 VSUBS 0.096588f
C5718 VDDD.n82 VSUBS 0.24113f
C5719 VDDD.n83 VSUBS 0.251622f
C5720 VDDD.n84 VSUBS 0.057151f
C5721 VDDD.t1032 VSUBS 0.337079f
C5722 VDDD.t1002 VSUBS 0.04923f
C5723 VDDD.t718 VSUBS 0.04923f
C5724 VDDD.n85 VSUBS 0.102503f
C5725 VDDD.n86 VSUBS 0.305072f
C5726 VDDD.n87 VSUBS 0.251622f
C5727 VDDD.n88 VSUBS 0.08621f
C5728 VDDD.t708 VSUBS 0.118653f
C5729 VDDD.n89 VSUBS 0.251622f
C5730 VDDD.t1313 VSUBS 0.032307f
C5731 VDDD.t1000 VSUBS 0.047863f
C5732 VDDD.n90 VSUBS 0.083298f
C5733 VDDD.n91 VSUBS 0.235104f
C5734 VDDD.n92 VSUBS 0.251622f
C5735 VDDD.n93 VSUBS 0.085726f
C5736 VDDD.t194 VSUBS 0.229702f
C5737 VDDD.n94 VSUBS 0.251622f
C5738 VDDD.n95 VSUBS 0.05037f
C5739 VDDD.t852 VSUBS 0.032307f
C5740 VDDD.t726 VSUBS 0.061025f
C5741 VDDD.n96 VSUBS 0.096588f
C5742 VDDD.n97 VSUBS 0.251622f
C5743 VDDD.t81 VSUBS 0.306728f
C5744 VDDD.n98 VSUBS 0.427682f
C5745 VDDD.n99 VSUBS 0.251622f
C5746 VDDD.n100 VSUBS 0.067806f
C5747 VDDD.n101 VSUBS 0.251622f
C5748 VDDD.n102 VSUBS 0.089116f
C5749 VDDD.n103 VSUBS 0.251622f
C5750 VDDD.t333 VSUBS 0.229702f
C5751 VDDD.n104 VSUBS 0.3381f
C5752 VDDD.n105 VSUBS 0.251622f
C5753 VDDD.t262 VSUBS 0.032307f
C5754 VDDD.t712 VSUBS 0.061025f
C5755 VDDD.n106 VSUBS 0.096588f
C5756 VDDD.n107 VSUBS 0.24113f
C5757 VDDD.n108 VSUBS 0.251622f
C5758 VDDD.n109 VSUBS 0.057151f
C5759 VDDD.t716 VSUBS 0.337079f
C5760 VDDD.t1175 VSUBS 0.04923f
C5761 VDDD.t918 VSUBS 0.04923f
C5762 VDDD.n110 VSUBS 0.102503f
C5763 VDDD.n111 VSUBS 0.305072f
C5764 VDDD.n112 VSUBS 0.251622f
C5765 VDDD.n113 VSUBS 0.08621f
C5766 VDDD.t706 VSUBS 0.118653f
C5767 VDDD.n114 VSUBS 0.251622f
C5768 VDDD.t1305 VSUBS 0.032307f
C5769 VDDD.t606 VSUBS 0.047863f
C5770 VDDD.n115 VSUBS 0.083298f
C5771 VDDD.n116 VSUBS 0.235104f
C5772 VDDD.n117 VSUBS 0.251622f
C5773 VDDD.n118 VSUBS 0.085726f
C5774 VDDD.t1196 VSUBS 0.229702f
C5775 VDDD.n119 VSUBS 0.251622f
C5776 VDDD.n120 VSUBS 0.05037f
C5777 VDDD.t503 VSUBS 0.032307f
C5778 VDDD.t337 VSUBS 0.061025f
C5779 VDDD.n121 VSUBS 0.096588f
C5780 VDDD.n122 VSUBS 0.251622f
C5781 VDDD.t335 VSUBS 0.306728f
C5782 VDDD.n123 VSUBS 0.427682f
C5783 VDDD.n124 VSUBS 0.251622f
C5784 VDDD.n125 VSUBS 0.067806f
C5785 VDDD.n126 VSUBS 0.251622f
C5786 VDDD.n127 VSUBS 0.089116f
C5787 VDDD.n128 VSUBS 0.251622f
C5788 VDDD.t1108 VSUBS 0.229702f
C5789 VDDD.n129 VSUBS 0.3381f
C5790 VDDD.n130 VSUBS 0.251622f
C5791 VDDD.t464 VSUBS 0.032307f
C5792 VDDD.t1010 VSUBS 0.061025f
C5793 VDDD.n131 VSUBS 0.096588f
C5794 VDDD.n132 VSUBS 0.24113f
C5795 VDDD.n133 VSUBS 0.251622f
C5796 VDDD.n134 VSUBS 0.057151f
C5797 VDDD.t118 VSUBS 0.337079f
C5798 VDDD.n135 VSUBS 0.251622f
C5799 VDDD.n136 VSUBS 0.032934f
C5800 VDDD.n137 VSUBS 0.251622f
C5801 VDDD.t1111 VSUBS 0.121884f
C5802 VDDD.n138 VSUBS 0.226774f
C5803 VDDD.n139 VSUBS 0.089116f
C5804 VDDD.n140 VSUBS 0.251622f
C5805 VDDD.n141 VSUBS 0.049401f
C5806 VDDD.n142 VSUBS 0.251622f
C5807 VDDD.t1220 VSUBS 0.032307f
C5808 VDDD.t541 VSUBS 0.047863f
C5809 VDDD.n143 VSUBS 0.083298f
C5810 VDDD.n144 VSUBS 0.235104f
C5811 VDDD.n145 VSUBS 0.08621f
C5812 VDDD.n146 VSUBS 0.251622f
C5813 VDDD.t20 VSUBS 0.04923f
C5814 VDDD.t285 VSUBS 0.04923f
C5815 VDDD.n147 VSUBS 0.102503f
C5816 VDDD.n148 VSUBS 0.305072f
C5817 VDDD.n149 VSUBS 0.057151f
C5818 VDDD.n150 VSUBS 0.251622f
C5819 VDDD.t312 VSUBS 0.032307f
C5820 VDDD.t898 VSUBS 0.061025f
C5821 VDDD.n151 VSUBS 0.096588f
C5822 VDDD.n152 VSUBS 0.24113f
C5823 VDDD.n153 VSUBS 0.251622f
C5824 VDDD.t1082 VSUBS 0.229702f
C5825 VDDD.n154 VSUBS 0.3381f
C5826 VDDD.n155 VSUBS 0.251622f
C5827 VDDD.n156 VSUBS 0.089116f
C5828 VDDD.n157 VSUBS 0.251622f
C5829 VDDD.n158 VSUBS 0.067806f
C5830 VDDD.n159 VSUBS 0.251622f
C5831 VDDD.t755 VSUBS 0.306728f
C5832 VDDD.n160 VSUBS 0.427682f
C5833 VDDD.n161 VSUBS 0.251622f
C5834 VDDD.t256 VSUBS 0.121884f
C5835 VDDD.n162 VSUBS 0.226774f
C5836 VDDD.n163 VSUBS 0.251622f
C5837 VDDD.n164 VSUBS 0.089116f
C5838 VDDD.n165 VSUBS 0.251622f
C5839 VDDD.n166 VSUBS 0.049401f
C5840 VDDD.n167 VSUBS 0.251622f
C5841 VDDD.t501 VSUBS 0.032307f
C5842 VDDD.t1299 VSUBS 0.047863f
C5843 VDDD.n168 VSUBS 0.083298f
C5844 VDDD.n169 VSUBS 0.235104f
C5845 VDDD.n170 VSUBS 0.08621f
C5846 VDDD.n171 VSUBS 0.251622f
C5847 VDDD.t153 VSUBS 0.04923f
C5848 VDDD.t984 VSUBS 0.04923f
C5849 VDDD.n172 VSUBS 0.102503f
C5850 VDDD.n173 VSUBS 0.305072f
C5851 VDDD.n174 VSUBS 0.057151f
C5852 VDDD.n175 VSUBS 0.251622f
C5853 VDDD.t820 VSUBS 0.032307f
C5854 VDDD.t33 VSUBS 0.061025f
C5855 VDDD.n176 VSUBS 0.096588f
C5856 VDDD.n177 VSUBS 0.24113f
C5857 VDDD.n178 VSUBS 0.251622f
C5858 VDDD.t260 VSUBS 0.229702f
C5859 VDDD.n179 VSUBS 0.3381f
C5860 VDDD.n180 VSUBS 0.251622f
C5861 VDDD.n181 VSUBS 0.089116f
C5862 VDDD.n182 VSUBS 0.251622f
C5863 VDDD.n183 VSUBS 0.067806f
C5864 VDDD.n184 VSUBS 0.251622f
C5865 VDDD.t1424 VSUBS 0.306728f
C5866 VDDD.n185 VSUBS 0.427682f
C5867 VDDD.n186 VSUBS 0.251622f
C5868 VDDD.t1160 VSUBS 0.121884f
C5869 VDDD.n187 VSUBS 0.226774f
C5870 VDDD.n188 VSUBS 0.251622f
C5871 VDDD.n189 VSUBS 0.089116f
C5872 VDDD.n190 VSUBS 0.251622f
C5873 VDDD.n191 VSUBS 0.049401f
C5874 VDDD.n192 VSUBS 0.251622f
C5875 VDDD.t466 VSUBS 0.032307f
C5876 VDDD.t1338 VSUBS 0.047863f
C5877 VDDD.n193 VSUBS 0.083298f
C5878 VDDD.n194 VSUBS 0.235104f
C5879 VDDD.n195 VSUBS 0.08621f
C5880 VDDD.n196 VSUBS 0.251622f
C5881 VDDD.t1404 VSUBS 0.04923f
C5882 VDDD.t538 VSUBS 0.04923f
C5883 VDDD.n197 VSUBS 0.102503f
C5884 VDDD.n198 VSUBS 0.305072f
C5885 VDDD.n199 VSUBS 0.057151f
C5886 VDDD.n200 VSUBS 0.251622f
C5887 VDDD.t1218 VSUBS 0.032307f
C5888 VDDD.t910 VSUBS 0.061025f
C5889 VDDD.n201 VSUBS 0.096588f
C5890 VDDD.n202 VSUBS 0.24113f
C5891 VDDD.n203 VSUBS 0.251622f
C5892 VDDD.t435 VSUBS 0.229702f
C5893 VDDD.n204 VSUBS 0.3381f
C5894 VDDD.n205 VSUBS 0.251622f
C5895 VDDD.n206 VSUBS 0.089116f
C5896 VDDD.n207 VSUBS 0.251622f
C5897 VDDD.n208 VSUBS 0.067806f
C5898 VDDD.n209 VSUBS 0.251622f
C5899 VDDD.t93 VSUBS 0.306728f
C5900 VDDD.n210 VSUBS 0.427682f
C5901 VDDD.n211 VSUBS 0.251622f
C5902 VDDD.t992 VSUBS 0.121884f
C5903 VDDD.n212 VSUBS 0.226774f
C5904 VDDD.n213 VSUBS 0.251622f
C5905 VDDD.n214 VSUBS 0.089116f
C5906 VDDD.n215 VSUBS 0.251622f
C5907 VDDD.n216 VSUBS 0.049401f
C5908 VDDD.n217 VSUBS 0.251622f
C5909 VDDD.t1317 VSUBS 0.032307f
C5910 VDDD.t530 VSUBS 0.047863f
C5911 VDDD.n218 VSUBS 0.083298f
C5912 VDDD.n219 VSUBS 0.235104f
C5913 VDDD.n220 VSUBS 0.08621f
C5914 VDDD.n221 VSUBS 0.251622f
C5915 VDDD.t59 VSUBS 0.04923f
C5916 VDDD.t1292 VSUBS 0.04923f
C5917 VDDD.n222 VSUBS 0.102503f
C5918 VDDD.n223 VSUBS 0.305072f
C5919 VDDD.n224 VSUBS 0.057151f
C5920 VDDD.n225 VSUBS 0.251622f
C5921 VDDD.t487 VSUBS 0.032307f
C5922 VDDD.t398 VSUBS 0.061025f
C5923 VDDD.n226 VSUBS 0.096588f
C5924 VDDD.n227 VSUBS 0.24113f
C5925 VDDD.n228 VSUBS 0.251622f
C5926 VDDD.t1074 VSUBS 0.229702f
C5927 VDDD.n229 VSUBS 0.3381f
C5928 VDDD.n230 VSUBS 0.251622f
C5929 VDDD.n231 VSUBS 0.089116f
C5930 VDDD.n232 VSUBS 0.251622f
C5931 VDDD.n233 VSUBS 0.067806f
C5932 VDDD.n234 VSUBS 0.251622f
C5933 VDDD.t749 VSUBS 0.306728f
C5934 VDDD.n235 VSUBS 0.427682f
C5935 VDDD.n236 VSUBS 0.251622f
C5936 VDDD.t1458 VSUBS 0.121884f
C5937 VDDD.n237 VSUBS 0.226774f
C5938 VDDD.n238 VSUBS 0.251622f
C5939 VDDD.n239 VSUBS 0.089116f
C5940 VDDD.n240 VSUBS 0.251622f
C5941 VDDD.n241 VSUBS 0.049401f
C5942 VDDD.n242 VSUBS 0.251622f
C5943 VDDD.t904 VSUBS 0.032307f
C5944 VDDD.t1379 VSUBS 0.047863f
C5945 VDDD.n243 VSUBS 0.083298f
C5946 VDDD.n244 VSUBS 0.235104f
C5947 VDDD.n245 VSUBS 0.08621f
C5948 VDDD.n246 VSUBS 0.251622f
C5949 VDDD.t807 VSUBS 0.04923f
C5950 VDDD.t85 VSUBS 0.04923f
C5951 VDDD.n247 VSUBS 0.102503f
C5952 VDDD.n248 VSUBS 0.305072f
C5953 VDDD.n249 VSUBS 0.057151f
C5954 VDDD.n250 VSUBS 0.251622f
C5955 VDDD.t785 VSUBS 0.032307f
C5956 VDDD.t1246 VSUBS 0.061025f
C5957 VDDD.n251 VSUBS 0.096588f
C5958 VDDD.n252 VSUBS 0.24113f
C5959 VDDD.n253 VSUBS 0.251622f
C5960 VDDD.t382 VSUBS 0.229702f
C5961 VDDD.n254 VSUBS 0.3381f
C5962 VDDD.n255 VSUBS 0.251622f
C5963 VDDD.n256 VSUBS 0.089116f
C5964 VDDD.n257 VSUBS 0.251622f
C5965 VDDD.n258 VSUBS 0.067806f
C5966 VDDD.n259 VSUBS 0.251622f
C5967 VDDD.n260 VSUBS 0.06829f
C5968 VDDD.n261 VSUBS 0.251622f
C5969 VDDD.n262 VSUBS 0.049401f
C5970 VDDD.n263 VSUBS 0.251622f
C5971 VDDD.t272 VSUBS 0.076922f
C5972 VDDD.t186 VSUBS 0.076922f
C5973 VDDD.n264 VSUBS 0.168898f
C5974 VDDD.n265 VSUBS 0.362323f
C5975 VDDD.n266 VSUBS 0.053276f
C5976 VDDD.n267 VSUBS 0.251622f
C5977 VDDD.t188 VSUBS 0.076922f
C5978 VDDD.t666 VSUBS 0.076922f
C5979 VDDD.n268 VSUBS 0.165125f
C5980 VDDD.n269 VSUBS 0.188262f
C5981 VDDD.t927 VSUBS 0.076922f
C5982 VDDD.t925 VSUBS 0.076922f
C5983 VDDD.n270 VSUBS 0.165125f
C5984 VDDD.n271 VSUBS 0.216855f
C5985 VDDD.n272 VSUBS 0.207246f
C5986 VDDD.n273 VSUBS 0.045527f
C5987 VDDD.n274 VSUBS 0.080398f
C5988 VDDD.n275 VSUBS 0.251622f
C5989 VDDD.n276 VSUBS 0.251622f
C5990 VDDD.n277 VSUBS 0.251622f
C5991 VDDD.n278 VSUBS 0.056666f
C5992 VDDD.t212 VSUBS 0.076922f
C5993 VDDD.t886 VSUBS 0.076922f
C5994 VDDD.n279 VSUBS 0.168898f
C5995 VDDD.n280 VSUBS 0.362323f
C5996 VDDD.n281 VSUBS 0.045042f
C5997 VDDD.n282 VSUBS 0.048917f
C5998 VDDD.n283 VSUBS 0.251622f
C5999 VDDD.n284 VSUBS 0.251622f
C6000 VDDD.n285 VSUBS 0.251622f
C6001 VDDD.t888 VSUBS 0.076922f
C6002 VDDD.t411 VSUBS 0.076922f
C6003 VDDD.n286 VSUBS 0.168898f
C6004 VDDD.n287 VSUBS 0.406881f
C6005 VDDD.n288 VSUBS 0.049401f
C6006 VDDD.t270 VSUBS 0.307526f
C6007 VDDD.n289 VSUBS 0.542325f
C6008 VDDD.n290 VSUBS 0.251622f
C6009 VDDD.n291 VSUBS 0.188716f
C6010 VDDD.n292 VSUBS 0.149059f
C6011 VDDD.n293 VSUBS 0.072165f
C6012 VDDD.t126 VSUBS 0.04923f
C6013 VDDD.t976 VSUBS 0.04923f
C6014 VDDD.n294 VSUBS 0.102503f
C6015 VDDD.n295 VSUBS 0.305072f
C6016 VDDD.n296 VSUBS 0.074102f
C6017 VDDD.n297 VSUBS 0.251622f
C6018 VDDD.n298 VSUBS 0.251622f
C6019 VDDD.n299 VSUBS 0.251622f
C6020 VDDD.t1453 VSUBS 0.118653f
C6021 VDDD.n300 VSUBS 0.250175f
C6022 VDDD.n301 VSUBS 0.08621f
C6023 VDDD.n302 VSUBS 0.089116f
C6024 VDDD.n303 VSUBS 0.251622f
C6025 VDDD.n304 VSUBS 0.251622f
C6026 VDDD.n305 VSUBS 0.251622f
C6027 VDDD.n306 VSUBS 0.052307f
C6028 VDDD.t631 VSUBS 0.032307f
C6029 VDDD.t1238 VSUBS 0.047863f
C6030 VDDD.n307 VSUBS 0.083298f
C6031 VDDD.n308 VSUBS 0.235104f
C6032 VDDD.n309 VSUBS 0.049401f
C6033 VDDD.n310 VSUBS 0.056666f
C6034 VDDD.n311 VSUBS 0.251622f
C6035 VDDD.n312 VSUBS 0.251622f
C6036 VDDD.n313 VSUBS 0.251622f
C6037 VDDD.n314 VSUBS 0.085726f
C6038 VDDD.n315 VSUBS 0.089116f
C6039 VDDD.n316 VSUBS 0.070712f
C6040 VDDD.n317 VSUBS 0.251622f
C6041 VDDD.n318 VSUBS 0.251622f
C6042 VDDD.n319 VSUBS 0.251622f
C6043 VDDD.n320 VSUBS 0.05037f
C6044 VDDD.t289 VSUBS 0.121884f
C6045 VDDD.n321 VSUBS 0.226774f
C6046 VDDD.n322 VSUBS 0.032934f
C6047 VDDD.t1248 VSUBS 0.337079f
C6048 VDDD.n323 VSUBS 0.521062f
C6049 VDDD.n324 VSUBS 0.251622f
C6050 VDDD.n325 VSUBS 0.251622f
C6051 VDDD.n326 VSUBS 0.188716f
C6052 VDDD.t161 VSUBS 0.306728f
C6053 VDDD.n327 VSUBS 0.427682f
C6054 VDDD.n328 VSUBS 0.062962f
C6055 VDDD.n329 VSUBS 0.149059f
C6056 VDDD.n330 VSUBS 0.251622f
C6057 VDDD.n331 VSUBS 0.251622f
C6058 VDDD.n332 VSUBS 0.074102f
C6059 VDDD.n333 VSUBS 0.067806f
C6060 VDDD.t661 VSUBS 0.118653f
C6061 VDDD.n334 VSUBS 0.250175f
C6062 VDDD.n335 VSUBS 0.251622f
C6063 VDDD.n336 VSUBS 0.251622f
C6064 VDDD.n337 VSUBS 0.251622f
C6065 VDDD.n338 VSUBS 0.089116f
C6066 VDDD.n339 VSUBS 0.089116f
C6067 VDDD.n340 VSUBS 0.052307f
C6068 VDDD.n341 VSUBS 0.251622f
C6069 VDDD.n342 VSUBS 0.251622f
C6070 VDDD.n343 VSUBS 0.251622f
C6071 VDDD.n344 VSUBS 0.056666f
C6072 VDDD.t459 VSUBS 0.229702f
C6073 VDDD.n345 VSUBS 0.3381f
C6074 VDDD.n346 VSUBS 0.085726f
C6075 VDDD.n347 VSUBS 0.251622f
C6076 VDDD.n348 VSUBS 0.251622f
C6077 VDDD.n349 VSUBS 0.251622f
C6078 VDDD.n350 VSUBS 0.070712f
C6079 VDDD.t493 VSUBS 0.032307f
C6080 VDDD.t929 VSUBS 0.061025f
C6081 VDDD.n351 VSUBS 0.096588f
C6082 VDDD.n352 VSUBS 0.24113f
C6083 VDDD.n353 VSUBS 0.05037f
C6084 VDDD.n354 VSUBS 0.251622f
C6085 VDDD.n355 VSUBS 0.251622f
C6086 VDDD.n356 VSUBS 0.032934f
C6087 VDDD.t862 VSUBS 0.337079f
C6088 VDDD.n357 VSUBS 0.521062f
C6089 VDDD.n358 VSUBS 0.057151f
C6090 VDDD.n359 VSUBS 0.251622f
C6091 VDDD.n360 VSUBS 0.188716f
C6092 VDDD.n361 VSUBS 0.149059f
C6093 VDDD.n362 VSUBS 0.062962f
C6094 VDDD.t834 VSUBS 0.04923f
C6095 VDDD.t668 VSUBS 0.04923f
C6096 VDDD.n363 VSUBS 0.102503f
C6097 VDDD.n364 VSUBS 0.305072f
C6098 VDDD.n365 VSUBS 0.074102f
C6099 VDDD.n366 VSUBS 0.251622f
C6100 VDDD.n367 VSUBS 0.251622f
C6101 VDDD.n368 VSUBS 0.251622f
C6102 VDDD.t37 VSUBS 0.118653f
C6103 VDDD.n369 VSUBS 0.250175f
C6104 VDDD.n370 VSUBS 0.08621f
C6105 VDDD.n371 VSUBS 0.089116f
C6106 VDDD.n372 VSUBS 0.251622f
C6107 VDDD.n373 VSUBS 0.251622f
C6108 VDDD.n374 VSUBS 0.251622f
C6109 VDDD.n375 VSUBS 0.052307f
C6110 VDDD.t900 VSUBS 0.032307f
C6111 VDDD.t798 VSUBS 0.047863f
C6112 VDDD.n376 VSUBS 0.083298f
C6113 VDDD.n377 VSUBS 0.235104f
C6114 VDDD.n378 VSUBS 0.049401f
C6115 VDDD.n379 VSUBS 0.056666f
C6116 VDDD.n380 VSUBS 0.251622f
C6117 VDDD.n381 VSUBS 0.251622f
C6118 VDDD.n382 VSUBS 0.251622f
C6119 VDDD.n383 VSUBS 0.085726f
C6120 VDDD.n384 VSUBS 0.089116f
C6121 VDDD.n385 VSUBS 0.070712f
C6122 VDDD.n386 VSUBS 0.251622f
C6123 VDDD.n387 VSUBS 0.251622f
C6124 VDDD.n388 VSUBS 0.251622f
C6125 VDDD.n389 VSUBS 0.05037f
C6126 VDDD.t1155 VSUBS 0.121884f
C6127 VDDD.n390 VSUBS 0.226774f
C6128 VDDD.n391 VSUBS 0.032934f
C6129 VDDD.t1336 VSUBS 0.337079f
C6130 VDDD.n392 VSUBS 0.521062f
C6131 VDDD.n393 VSUBS 0.251622f
C6132 VDDD.n394 VSUBS 0.251622f
C6133 VDDD.n395 VSUBS 0.188716f
C6134 VDDD.t1350 VSUBS 0.306728f
C6135 VDDD.n396 VSUBS 0.427682f
C6136 VDDD.n397 VSUBS 0.062962f
C6137 VDDD.n398 VSUBS 0.149059f
C6138 VDDD.n399 VSUBS 0.251622f
C6139 VDDD.n400 VSUBS 0.251622f
C6140 VDDD.n401 VSUBS 0.074102f
C6141 VDDD.n402 VSUBS 0.067806f
C6142 VDDD.t236 VSUBS 0.118653f
C6143 VDDD.n403 VSUBS 0.250175f
C6144 VDDD.n404 VSUBS 0.251622f
C6145 VDDD.n405 VSUBS 0.251622f
C6146 VDDD.n406 VSUBS 0.251622f
C6147 VDDD.n407 VSUBS 0.089116f
C6148 VDDD.n408 VSUBS 0.089116f
C6149 VDDD.n409 VSUBS 0.052307f
C6150 VDDD.n410 VSUBS 0.251622f
C6151 VDDD.n411 VSUBS 0.251622f
C6152 VDDD.n412 VSUBS 0.251622f
C6153 VDDD.n413 VSUBS 0.056666f
C6154 VDDD.t62 VSUBS 0.229702f
C6155 VDDD.n414 VSUBS 0.3381f
C6156 VDDD.n415 VSUBS 0.085726f
C6157 VDDD.n416 VSUBS 0.251622f
C6158 VDDD.n417 VSUBS 0.251622f
C6159 VDDD.n418 VSUBS 0.251622f
C6160 VDDD.n419 VSUBS 0.070712f
C6161 VDDD.t915 VSUBS 0.032307f
C6162 VDDD.t244 VSUBS 0.061025f
C6163 VDDD.n420 VSUBS 0.096588f
C6164 VDDD.n421 VSUBS 0.24113f
C6165 VDDD.n422 VSUBS 0.05037f
C6166 VDDD.n423 VSUBS 0.251622f
C6167 VDDD.n424 VSUBS 0.251622f
C6168 VDDD.n425 VSUBS 0.032934f
C6169 VDDD.t91 VSUBS 0.337079f
C6170 VDDD.n426 VSUBS 0.521062f
C6171 VDDD.n427 VSUBS 0.057151f
C6172 VDDD.n428 VSUBS 0.251622f
C6173 VDDD.n429 VSUBS 0.188716f
C6174 VDDD.n430 VSUBS 0.149059f
C6175 VDDD.n431 VSUBS 0.062962f
C6176 VDDD.t761 VSUBS 0.04923f
C6177 VDDD.t3 VSUBS 0.04923f
C6178 VDDD.n432 VSUBS 0.102503f
C6179 VDDD.n433 VSUBS 0.305072f
C6180 VDDD.n434 VSUBS 0.074102f
C6181 VDDD.n435 VSUBS 0.251622f
C6182 VDDD.n436 VSUBS 0.251622f
C6183 VDDD.n437 VSUBS 0.251622f
C6184 VDDD.t100 VSUBS 0.118653f
C6185 VDDD.n438 VSUBS 0.250175f
C6186 VDDD.n439 VSUBS 0.08621f
C6187 VDDD.n440 VSUBS 0.089116f
C6188 VDDD.n441 VSUBS 0.251622f
C6189 VDDD.n442 VSUBS 0.251622f
C6190 VDDD.n443 VSUBS 0.251622f
C6191 VDDD.n444 VSUBS 0.052307f
C6192 VDDD.t1216 VSUBS 0.032307f
C6193 VDDD.t890 VSUBS 0.047863f
C6194 VDDD.n445 VSUBS 0.083298f
C6195 VDDD.n446 VSUBS 0.235104f
C6196 VDDD.n447 VSUBS 0.049401f
C6197 VDDD.n448 VSUBS 0.056666f
C6198 VDDD.n449 VSUBS 0.251622f
C6199 VDDD.n450 VSUBS 0.251622f
C6200 VDDD.n451 VSUBS 0.251622f
C6201 VDDD.n452 VSUBS 0.085726f
C6202 VDDD.n453 VSUBS 0.089116f
C6203 VDDD.n454 VSUBS 0.070712f
C6204 VDDD.n455 VSUBS 0.251622f
C6205 VDDD.n456 VSUBS 0.251622f
C6206 VDDD.n457 VSUBS 0.251622f
C6207 VDDD.n458 VSUBS 0.05037f
C6208 VDDD.t551 VSUBS 0.121884f
C6209 VDDD.n459 VSUBS 0.226774f
C6210 VDDD.n460 VSUBS 0.032934f
C6211 VDDD.t218 VSUBS 0.337079f
C6212 VDDD.n461 VSUBS 0.521062f
C6213 VDDD.n462 VSUBS 0.251622f
C6214 VDDD.n463 VSUBS 0.251622f
C6215 VDDD.n464 VSUBS 0.188716f
C6216 VDDD.t220 VSUBS 0.306728f
C6217 VDDD.n465 VSUBS 0.427682f
C6218 VDDD.n466 VSUBS 0.062962f
C6219 VDDD.n467 VSUBS 0.149059f
C6220 VDDD.n468 VSUBS 0.251622f
C6221 VDDD.n469 VSUBS 0.251622f
C6222 VDDD.n470 VSUBS 0.074102f
C6223 VDDD.n471 VSUBS 0.067806f
C6224 VDDD.t417 VSUBS 0.118653f
C6225 VDDD.n472 VSUBS 0.250175f
C6226 VDDD.n473 VSUBS 0.251622f
C6227 VDDD.n474 VSUBS 0.251622f
C6228 VDDD.n475 VSUBS 0.251622f
C6229 VDDD.n476 VSUBS 0.089116f
C6230 VDDD.n477 VSUBS 0.089116f
C6231 VDDD.n478 VSUBS 0.052307f
C6232 VDDD.n479 VSUBS 0.251622f
C6233 VDDD.n480 VSUBS 0.251622f
C6234 VDDD.n481 VSUBS 0.251622f
C6235 VDDD.n482 VSUBS 0.056666f
C6236 VDDD.t1067 VSUBS 0.229702f
C6237 VDDD.n483 VSUBS 0.3381f
C6238 VDDD.n484 VSUBS 0.085726f
C6239 VDDD.n485 VSUBS 0.251622f
C6240 VDDD.n486 VSUBS 0.251622f
C6241 VDDD.n487 VSUBS 0.251622f
C6242 VDDD.n488 VSUBS 0.070712f
C6243 VDDD.t1188 VSUBS 0.032307f
C6244 VDDD.t1014 VSUBS 0.061025f
C6245 VDDD.n489 VSUBS 0.096588f
C6246 VDDD.n490 VSUBS 0.24113f
C6247 VDDD.n491 VSUBS 0.05037f
C6248 VDDD.n492 VSUBS 0.251622f
C6249 VDDD.n493 VSUBS 0.251622f
C6250 VDDD.n494 VSUBS 0.032934f
C6251 VDDD.t1012 VSUBS 0.337079f
C6252 VDDD.n495 VSUBS 0.521062f
C6253 VDDD.n496 VSUBS 0.057151f
C6254 VDDD.n497 VSUBS 0.251622f
C6255 VDDD.n498 VSUBS 0.188716f
C6256 VDDD.n499 VSUBS 0.149059f
C6257 VDDD.n500 VSUBS 0.062962f
C6258 VDDD.t210 VSUBS 0.04923f
C6259 VDDD.t132 VSUBS 0.04923f
C6260 VDDD.n501 VSUBS 0.102503f
C6261 VDDD.n502 VSUBS 0.305072f
C6262 VDDD.n503 VSUBS 0.074102f
C6263 VDDD.n504 VSUBS 0.251622f
C6264 VDDD.n505 VSUBS 0.251622f
C6265 VDDD.n506 VSUBS 0.251622f
C6266 VDDD.t238 VSUBS 0.118653f
C6267 VDDD.n507 VSUBS 0.250175f
C6268 VDDD.n508 VSUBS 0.08621f
C6269 VDDD.n509 VSUBS 0.089116f
C6270 VDDD.n510 VSUBS 0.251622f
C6271 VDDD.n511 VSUBS 0.251622f
C6272 VDDD.n512 VSUBS 0.251622f
C6273 VDDD.n513 VSUBS 0.052307f
C6274 VDDD.t824 VSUBS 0.032307f
C6275 VDDD.t836 VSUBS 0.047863f
C6276 VDDD.n514 VSUBS 0.083298f
C6277 VDDD.n515 VSUBS 0.235104f
C6278 VDDD.n516 VSUBS 0.049401f
C6279 VDDD.n517 VSUBS 0.056666f
C6280 VDDD.n518 VSUBS 0.251622f
C6281 VDDD.n519 VSUBS 0.251622f
C6282 VDDD.n520 VSUBS 0.251622f
C6283 VDDD.n521 VSUBS 0.085726f
C6284 VDDD.n522 VSUBS 0.089116f
C6285 VDDD.n523 VSUBS 0.070712f
C6286 VDDD.n524 VSUBS 0.251622f
C6287 VDDD.n525 VSUBS 0.251622f
C6288 VDDD.n526 VSUBS 0.251622f
C6289 VDDD.n527 VSUBS 0.05037f
C6290 VDDD.t563 VSUBS 0.121884f
C6291 VDDD.n528 VSUBS 0.226774f
C6292 VDDD.n529 VSUBS 0.032934f
C6293 VDDD.t35 VSUBS 0.337079f
C6294 VDDD.n530 VSUBS 0.521062f
C6295 VDDD.n531 VSUBS 0.251622f
C6296 VDDD.n532 VSUBS 0.251622f
C6297 VDDD.n533 VSUBS 0.188716f
C6298 VDDD.t1385 VSUBS 0.306728f
C6299 VDDD.n534 VSUBS 0.427682f
C6300 VDDD.n535 VSUBS 0.062962f
C6301 VDDD.n536 VSUBS 0.149059f
C6302 VDDD.n537 VSUBS 0.251622f
C6303 VDDD.n538 VSUBS 0.251622f
C6304 VDDD.n539 VSUBS 0.074102f
C6305 VDDD.n540 VSUBS 0.067806f
C6306 VDDD.t663 VSUBS 0.118653f
C6307 VDDD.n541 VSUBS 0.250175f
C6308 VDDD.n542 VSUBS 0.251622f
C6309 VDDD.n543 VSUBS 0.251622f
C6310 VDDD.n544 VSUBS 0.251622f
C6311 VDDD.n545 VSUBS 0.089116f
C6312 VDDD.n546 VSUBS 0.089116f
C6313 VDDD.n547 VSUBS 0.052307f
C6314 VDDD.n548 VSUBS 0.251622f
C6315 VDDD.n549 VSUBS 0.251622f
C6316 VDDD.n550 VSUBS 0.251622f
C6317 VDDD.n551 VSUBS 0.056666f
C6318 VDDD.t1228 VSUBS 0.229702f
C6319 VDDD.n552 VSUBS 0.3381f
C6320 VDDD.n553 VSUBS 0.085726f
C6321 VDDD.n554 VSUBS 0.251622f
C6322 VDDD.n555 VSUBS 0.251622f
C6323 VDDD.n556 VSUBS 0.251622f
C6324 VDDD.n557 VSUBS 0.070712f
C6325 VDDD.t1269 VSUBS 0.032307f
C6326 VDDD.t702 VSUBS 0.061025f
C6327 VDDD.n558 VSUBS 0.096588f
C6328 VDDD.n559 VSUBS 0.24113f
C6329 VDDD.n560 VSUBS 0.05037f
C6330 VDDD.n561 VSUBS 0.251622f
C6331 VDDD.n562 VSUBS 0.251622f
C6332 VDDD.n563 VSUBS 0.032934f
C6333 VDDD.t700 VSUBS 0.337079f
C6334 VDDD.n564 VSUBS 0.521062f
C6335 VDDD.n565 VSUBS 0.057151f
C6336 VDDD.n566 VSUBS 0.251622f
C6337 VDDD.n567 VSUBS 0.188716f
C6338 VDDD.n568 VSUBS 0.149059f
C6339 VDDD.n569 VSUBS 0.062962f
C6340 VDDD.t1103 VSUBS 0.04923f
C6341 VDDD.t645 VSUBS 0.04923f
C6342 VDDD.n570 VSUBS 0.102503f
C6343 VDDD.n571 VSUBS 0.305072f
C6344 VDDD.n572 VSUBS 0.074102f
C6345 VDDD.n573 VSUBS 0.251622f
C6346 VDDD.n574 VSUBS 0.251622f
C6347 VDDD.n575 VSUBS 0.251622f
C6348 VDDD.t98 VSUBS 0.118653f
C6349 VDDD.n576 VSUBS 0.250175f
C6350 VDDD.n577 VSUBS 0.08621f
C6351 VDDD.n578 VSUBS 0.089116f
C6352 VDDD.n579 VSUBS 0.251622f
C6353 VDDD.n580 VSUBS 0.251622f
C6354 VDDD.n581 VSUBS 0.251622f
C6355 VDDD.n582 VSUBS 0.052307f
C6356 VDDD.t616 VSUBS 0.032307f
C6357 VDDD.t612 VSUBS 0.047863f
C6358 VDDD.n583 VSUBS 0.083298f
C6359 VDDD.n584 VSUBS 0.235104f
C6360 VDDD.n585 VSUBS 0.049401f
C6361 VDDD.n586 VSUBS 0.056666f
C6362 VDDD.n587 VSUBS 0.251622f
C6363 VDDD.n588 VSUBS 0.251622f
C6364 VDDD.n589 VSUBS 0.251622f
C6365 VDDD.n590 VSUBS 0.085726f
C6366 VDDD.n591 VSUBS 0.089116f
C6367 VDDD.n592 VSUBS 0.070712f
C6368 VDDD.n593 VSUBS 0.251622f
C6369 VDDD.n594 VSUBS 0.251622f
C6370 VDDD.n595 VSUBS 0.251622f
C6371 VDDD.n596 VSUBS 0.05037f
C6372 VDDD.t932 VSUBS 0.121884f
C6373 VDDD.n597 VSUBS 0.226774f
C6374 VDDD.n598 VSUBS 0.032934f
C6375 VDDD.t1145 VSUBS 0.337079f
C6376 VDDD.n599 VSUBS 0.521062f
C6377 VDDD.n600 VSUBS 0.251622f
C6378 VDDD.n601 VSUBS 0.251622f
C6379 VDDD.n602 VSUBS 0.188716f
C6380 VDDD.t1147 VSUBS 0.306728f
C6381 VDDD.n603 VSUBS 0.427682f
C6382 VDDD.n604 VSUBS 0.062962f
C6383 VDDD.n605 VSUBS 0.149059f
C6384 VDDD.n606 VSUBS 0.251622f
C6385 VDDD.n607 VSUBS 0.251622f
C6386 VDDD.n608 VSUBS 0.074102f
C6387 VDDD.n609 VSUBS 0.067806f
C6388 VDDD.t1451 VSUBS 0.118653f
C6389 VDDD.n610 VSUBS 0.250175f
C6390 VDDD.n611 VSUBS 0.251622f
C6391 VDDD.n612 VSUBS 0.251622f
C6392 VDDD.n613 VSUBS 0.251622f
C6393 VDDD.n614 VSUBS 0.089116f
C6394 VDDD.n615 VSUBS 0.089116f
C6395 VDDD.n616 VSUBS 0.052307f
C6396 VDDD.n617 VSUBS 0.251622f
C6397 VDDD.n618 VSUBS 0.251622f
C6398 VDDD.n619 VSUBS 0.251622f
C6399 VDDD.n620 VSUBS 0.056666f
C6400 VDDD.t1236 VSUBS 0.229702f
C6401 VDDD.n621 VSUBS 0.3381f
C6402 VDDD.n622 VSUBS 0.085726f
C6403 VDDD.n623 VSUBS 0.251622f
C6404 VDDD.n624 VSUBS 0.251622f
C6405 VDDD.n625 VSUBS 0.251622f
C6406 VDDD.n626 VSUBS 0.070712f
C6407 VDDD.t489 VSUBS 0.032307f
C6408 VDDD.t602 VSUBS 0.061025f
C6409 VDDD.n627 VSUBS 0.096588f
C6410 VDDD.n628 VSUBS 0.24113f
C6411 VDDD.n629 VSUBS 0.05037f
C6412 VDDD.n630 VSUBS 0.251622f
C6413 VDDD.n631 VSUBS 0.251622f
C6414 VDDD.n632 VSUBS 0.251622f
C6415 VDDD.t1372 VSUBS 0.337079f
C6416 VDDD.n633 VSUBS 0.521062f
C6417 VDDD.n634 VSUBS 0.057151f
C6418 VDDD.t1370 VSUBS 0.306728f
C6419 VDDD.n635 VSUBS 0.366172f
C6420 VDDD.n636 VSUBS 2.02392f
C6421 VDDD.t1008 VSUBS 0.306728f
C6422 VDDD.n637 VSUBS 0.366173f
C6423 VDDD.n638 VSUBS 2.02392f
C6424 VDDD.n639 VSUBS 0.251622f
C6425 VDDD.n640 VSUBS 0.251622f
C6426 VDDD.n641 VSUBS 0.521063f
C6427 VDDD.n642 VSUBS 0.032934f
C6428 VDDD.t692 VSUBS 0.121884f
C6429 VDDD.n643 VSUBS 0.226774f
C6430 VDDD.n644 VSUBS 0.05037f
C6431 VDDD.n645 VSUBS 0.251622f
C6432 VDDD.n646 VSUBS 0.251622f
C6433 VDDD.n647 VSUBS 0.251622f
C6434 VDDD.n648 VSUBS 0.070712f
C6435 VDDD.n649 VSUBS 0.089116f
C6436 VDDD.n650 VSUBS 0.085726f
C6437 VDDD.n651 VSUBS 0.251622f
C6438 VDDD.n652 VSUBS 0.251622f
C6439 VDDD.n653 VSUBS 0.251622f
C6440 VDDD.n654 VSUBS 0.056666f
C6441 VDDD.n655 VSUBS 0.049401f
C6442 VDDD.t906 VSUBS 0.032307f
C6443 VDDD.t1356 VSUBS 0.047863f
C6444 VDDD.n656 VSUBS 0.083298f
C6445 VDDD.n657 VSUBS 0.235104f
C6446 VDDD.n658 VSUBS 0.052307f
C6447 VDDD.n659 VSUBS 0.251622f
C6448 VDDD.n660 VSUBS 0.251622f
C6449 VDDD.n661 VSUBS 0.251622f
C6450 VDDD.n662 VSUBS 0.089116f
C6451 VDDD.n663 VSUBS 0.08621f
C6452 VDDD.t1038 VSUBS 0.118653f
C6453 VDDD.n664 VSUBS 0.250175f
C6454 VDDD.n665 VSUBS 0.251622f
C6455 VDDD.n666 VSUBS 0.251622f
C6456 VDDD.n667 VSUBS 0.251622f
C6457 VDDD.n668 VSUBS 0.074102f
C6458 VDDD.t949 VSUBS 0.04923f
C6459 VDDD.t283 VSUBS 0.04923f
C6460 VDDD.n669 VSUBS 0.102503f
C6461 VDDD.n670 VSUBS 0.305072f
C6462 VDDD.n671 VSUBS 0.062962f
C6463 VDDD.n672 VSUBS 0.149059f
C6464 VDDD.n673 VSUBS 0.188716f
C6465 VDDD.n674 VSUBS 0.251622f
C6466 VDDD.n675 VSUBS 0.057151f
C6467 VDDD.t1387 VSUBS 0.337079f
C6468 VDDD.n676 VSUBS 0.521063f
C6469 VDDD.t732 VSUBS 0.121884f
C6470 VDDD.n677 VSUBS 0.226774f
C6471 VDDD.n678 VSUBS 0.032934f
C6472 VDDD.n679 VSUBS 0.251622f
C6473 VDDD.n680 VSUBS 0.251622f
C6474 VDDD.n681 VSUBS 0.251622f
C6475 VDDD.n682 VSUBS 0.24113f
C6476 VDDD.n683 VSUBS 0.070712f
C6477 VDDD.n684 VSUBS 0.089116f
C6478 VDDD.n685 VSUBS 0.251622f
C6479 VDDD.n686 VSUBS 0.251622f
C6480 VDDD.n687 VSUBS 0.251622f
C6481 VDDD.n688 VSUBS 0.3381f
C6482 VDDD.n689 VSUBS 0.056666f
C6483 VDDD.n690 VSUBS 0.049401f
C6484 VDDD.n691 VSUBS 0.251622f
C6485 VDDD.n692 VSUBS 0.251622f
C6486 VDDD.n693 VSUBS 0.052307f
C6487 VDDD.n694 VSUBS 0.089116f
C6488 VDDD.n695 VSUBS 0.089116f
C6489 VDDD.n696 VSUBS 0.251622f
C6490 VDDD.n697 VSUBS 0.251622f
C6491 VDDD.n698 VSUBS 0.251622f
C6492 VDDD.n699 VSUBS 0.250175f
C6493 VDDD.n700 VSUBS 0.067806f
C6494 VDDD.n701 VSUBS 0.074102f
C6495 VDDD.n702 VSUBS 0.251622f
C6496 VDDD.n703 VSUBS 0.251622f
C6497 VDDD.n704 VSUBS 0.149059f
C6498 VDDD.n705 VSUBS 0.062962f
C6499 VDDD.t714 VSUBS 0.306728f
C6500 VDDD.n706 VSUBS 0.427682f
C6501 VDDD.n707 VSUBS 0.188716f
C6502 VDDD.n708 VSUBS 0.251622f
C6503 VDDD.n709 VSUBS 0.251622f
C6504 VDDD.n710 VSUBS 0.521063f
C6505 VDDD.n711 VSUBS 0.032934f
C6506 VDDD.t581 VSUBS 0.121884f
C6507 VDDD.n712 VSUBS 0.226774f
C6508 VDDD.n713 VSUBS 0.05037f
C6509 VDDD.n714 VSUBS 0.251622f
C6510 VDDD.n715 VSUBS 0.251622f
C6511 VDDD.n716 VSUBS 0.251622f
C6512 VDDD.n717 VSUBS 0.070712f
C6513 VDDD.n718 VSUBS 0.089116f
C6514 VDDD.n719 VSUBS 0.085726f
C6515 VDDD.n720 VSUBS 0.251622f
C6516 VDDD.n721 VSUBS 0.251622f
C6517 VDDD.n722 VSUBS 0.251622f
C6518 VDDD.n723 VSUBS 0.056666f
C6519 VDDD.n724 VSUBS 0.049401f
C6520 VDDD.t614 VSUBS 0.032307f
C6521 VDDD.t809 VSUBS 0.047863f
C6522 VDDD.n725 VSUBS 0.083298f
C6523 VDDD.n726 VSUBS 0.235104f
C6524 VDDD.n727 VSUBS 0.052307f
C6525 VDDD.n728 VSUBS 0.251622f
C6526 VDDD.n729 VSUBS 0.251622f
C6527 VDDD.n730 VSUBS 0.251622f
C6528 VDDD.n731 VSUBS 0.089116f
C6529 VDDD.n732 VSUBS 0.08621f
C6530 VDDD.t1121 VSUBS 0.118653f
C6531 VDDD.n733 VSUBS 0.250175f
C6532 VDDD.n734 VSUBS 0.251622f
C6533 VDDD.n735 VSUBS 0.251622f
C6534 VDDD.n736 VSUBS 0.251622f
C6535 VDDD.n737 VSUBS 0.074102f
C6536 VDDD.t275 VSUBS 0.04923f
C6537 VDDD.t242 VSUBS 0.04923f
C6538 VDDD.n738 VSUBS 0.102503f
C6539 VDDD.n739 VSUBS 0.305072f
C6540 VDDD.n740 VSUBS 0.062962f
C6541 VDDD.n741 VSUBS 0.149059f
C6542 VDDD.n742 VSUBS 0.188716f
C6543 VDDD.n743 VSUBS 0.251622f
C6544 VDDD.n744 VSUBS 0.057151f
C6545 VDDD.t771 VSUBS 0.337079f
C6546 VDDD.n745 VSUBS 0.521063f
C6547 VDDD.t604 VSUBS 0.121884f
C6548 VDDD.n746 VSUBS 0.226774f
C6549 VDDD.n747 VSUBS 0.032934f
C6550 VDDD.n748 VSUBS 0.251622f
C6551 VDDD.n749 VSUBS 0.251622f
C6552 VDDD.n750 VSUBS 0.251622f
C6553 VDDD.n751 VSUBS 0.24113f
C6554 VDDD.n752 VSUBS 0.070712f
C6555 VDDD.n753 VSUBS 0.089116f
C6556 VDDD.n754 VSUBS 0.251622f
C6557 VDDD.n755 VSUBS 0.251622f
C6558 VDDD.n756 VSUBS 0.251622f
C6559 VDDD.n757 VSUBS 0.3381f
C6560 VDDD.n758 VSUBS 0.056666f
C6561 VDDD.n759 VSUBS 0.049401f
C6562 VDDD.n760 VSUBS 0.251622f
C6563 VDDD.n761 VSUBS 0.251622f
C6564 VDDD.n762 VSUBS 0.052307f
C6565 VDDD.n763 VSUBS 0.089116f
C6566 VDDD.n764 VSUBS 0.089116f
C6567 VDDD.n765 VSUBS 0.251622f
C6568 VDDD.n766 VSUBS 0.251622f
C6569 VDDD.n767 VSUBS 0.251622f
C6570 VDDD.n768 VSUBS 0.250175f
C6571 VDDD.n769 VSUBS 0.067806f
C6572 VDDD.n770 VSUBS 0.074102f
C6573 VDDD.n771 VSUBS 0.251622f
C6574 VDDD.n772 VSUBS 0.251622f
C6575 VDDD.n773 VSUBS 0.149059f
C6576 VDDD.n774 VSUBS 0.062962f
C6577 VDDD.t1036 VSUBS 0.306728f
C6578 VDDD.n775 VSUBS 0.427682f
C6579 VDDD.n776 VSUBS 0.188716f
C6580 VDDD.n777 VSUBS 0.251622f
C6581 VDDD.n778 VSUBS 0.251622f
C6582 VDDD.n779 VSUBS 0.521063f
C6583 VDDD.n780 VSUBS 0.032934f
C6584 VDDD.t64 VSUBS 0.121884f
C6585 VDDD.n781 VSUBS 0.226774f
C6586 VDDD.n782 VSUBS 0.05037f
C6587 VDDD.n783 VSUBS 0.251622f
C6588 VDDD.n784 VSUBS 0.251622f
C6589 VDDD.n785 VSUBS 0.251622f
C6590 VDDD.n786 VSUBS 0.070712f
C6591 VDDD.n787 VSUBS 0.089116f
C6592 VDDD.n788 VSUBS 0.085726f
C6593 VDDD.n789 VSUBS 0.251622f
C6594 VDDD.n790 VSUBS 0.251622f
C6595 VDDD.n791 VSUBS 0.251622f
C6596 VDDD.n792 VSUBS 0.056666f
C6597 VDDD.n793 VSUBS 0.049401f
C6598 VDDD.t172 VSUBS 0.032307f
C6599 VDDD.t142 VSUBS 0.047863f
C6600 VDDD.n794 VSUBS 0.083298f
C6601 VDDD.n795 VSUBS 0.235104f
C6602 VDDD.n796 VSUBS 0.052307f
C6603 VDDD.n797 VSUBS 0.251622f
C6604 VDDD.n798 VSUBS 0.251622f
C6605 VDDD.n799 VSUBS 0.251622f
C6606 VDDD.n800 VSUBS 0.089116f
C6607 VDDD.n801 VSUBS 0.08621f
C6608 VDDD.t1123 VSUBS 0.118653f
C6609 VDDD.n802 VSUBS 0.250175f
C6610 VDDD.n803 VSUBS 0.251622f
C6611 VDDD.n804 VSUBS 0.251622f
C6612 VDDD.n805 VSUBS 0.251622f
C6613 VDDD.n806 VSUBS 0.074102f
C6614 VDDD.t753 VSUBS 0.04923f
C6615 VDDD.t536 VSUBS 0.04923f
C6616 VDDD.n807 VSUBS 0.102503f
C6617 VDDD.n808 VSUBS 0.305072f
C6618 VDDD.n809 VSUBS 0.062962f
C6619 VDDD.n810 VSUBS 0.149059f
C6620 VDDD.n811 VSUBS 0.188716f
C6621 VDDD.n812 VSUBS 0.251622f
C6622 VDDD.n813 VSUBS 0.057151f
C6623 VDDD.t147 VSUBS 0.337079f
C6624 VDDD.n814 VSUBS 0.521063f
C6625 VDDD.t302 VSUBS 0.121884f
C6626 VDDD.n815 VSUBS 0.226774f
C6627 VDDD.n816 VSUBS 0.032934f
C6628 VDDD.n817 VSUBS 0.251622f
C6629 VDDD.n818 VSUBS 0.251622f
C6630 VDDD.n819 VSUBS 0.251622f
C6631 VDDD.n820 VSUBS 0.24113f
C6632 VDDD.n821 VSUBS 0.070712f
C6633 VDDD.n822 VSUBS 0.089116f
C6634 VDDD.n823 VSUBS 0.251622f
C6635 VDDD.n824 VSUBS 0.251622f
C6636 VDDD.n825 VSUBS 0.251622f
C6637 VDDD.n826 VSUBS 0.3381f
C6638 VDDD.n827 VSUBS 0.056666f
C6639 VDDD.n828 VSUBS 0.049401f
C6640 VDDD.n829 VSUBS 0.251622f
C6641 VDDD.n830 VSUBS 0.251622f
C6642 VDDD.n831 VSUBS 0.052307f
C6643 VDDD.n832 VSUBS 0.089116f
C6644 VDDD.n833 VSUBS 0.089116f
C6645 VDDD.n834 VSUBS 0.251622f
C6646 VDDD.n835 VSUBS 0.251622f
C6647 VDDD.n836 VSUBS 0.251622f
C6648 VDDD.n837 VSUBS 0.250175f
C6649 VDDD.n838 VSUBS 0.067806f
C6650 VDDD.n839 VSUBS 0.074102f
C6651 VDDD.n840 VSUBS 0.251622f
C6652 VDDD.n841 VSUBS 0.251622f
C6653 VDDD.n842 VSUBS 0.149059f
C6654 VDDD.n843 VSUBS 0.062962f
C6655 VDDD.t1358 VSUBS 0.306728f
C6656 VDDD.n844 VSUBS 0.427682f
C6657 VDDD.n845 VSUBS 0.188716f
C6658 VDDD.n846 VSUBS 0.251622f
C6659 VDDD.n847 VSUBS 0.251622f
C6660 VDDD.n848 VSUBS 0.521063f
C6661 VDDD.n849 VSUBS 0.032934f
C6662 VDDD.t737 VSUBS 0.121884f
C6663 VDDD.n850 VSUBS 0.226774f
C6664 VDDD.n851 VSUBS 0.05037f
C6665 VDDD.n852 VSUBS 0.251622f
C6666 VDDD.n853 VSUBS 0.251622f
C6667 VDDD.n854 VSUBS 0.251622f
C6668 VDDD.n855 VSUBS 0.070712f
C6669 VDDD.n856 VSUBS 0.089116f
C6670 VDDD.n857 VSUBS 0.085726f
C6671 VDDD.n858 VSUBS 0.251622f
C6672 VDDD.n859 VSUBS 0.251622f
C6673 VDDD.n860 VSUBS 0.251622f
C6674 VDDD.n861 VSUBS 0.056666f
C6675 VDDD.n862 VSUBS 0.049401f
C6676 VDDD.t547 VSUBS 0.032307f
C6677 VDDD.t746 VSUBS 0.047863f
C6678 VDDD.n863 VSUBS 0.083298f
C6679 VDDD.n864 VSUBS 0.235104f
C6680 VDDD.n865 VSUBS 0.052307f
C6681 VDDD.n866 VSUBS 0.251622f
C6682 VDDD.n867 VSUBS 0.251622f
C6683 VDDD.n868 VSUBS 0.251622f
C6684 VDDD.n869 VSUBS 0.089116f
C6685 VDDD.n870 VSUBS 0.08621f
C6686 VDDD.t1040 VSUBS 0.118653f
C6687 VDDD.n871 VSUBS 0.250175f
C6688 VDDD.n872 VSUBS 0.251622f
C6689 VDDD.n873 VSUBS 0.251622f
C6690 VDDD.n874 VSUBS 0.251622f
C6691 VDDD.n875 VSUBS 0.074102f
C6692 VDDD.t592 VSUBS 0.04923f
C6693 VDDD.t1288 VSUBS 0.04923f
C6694 VDDD.n876 VSUBS 0.102503f
C6695 VDDD.n877 VSUBS 0.305072f
C6696 VDDD.n878 VSUBS 0.062962f
C6697 VDDD.n879 VSUBS 0.149059f
C6698 VDDD.n880 VSUBS 0.188716f
C6699 VDDD.n881 VSUBS 0.251622f
C6700 VDDD.n882 VSUBS 0.057151f
C6701 VDDD.t79 VSUBS 0.337079f
C6702 VDDD.n883 VSUBS 0.521063f
C6703 VDDD.t696 VSUBS 0.121884f
C6704 VDDD.n884 VSUBS 0.226774f
C6705 VDDD.n885 VSUBS 0.032934f
C6706 VDDD.n886 VSUBS 0.251622f
C6707 VDDD.n887 VSUBS 0.251622f
C6708 VDDD.n888 VSUBS 0.251622f
C6709 VDDD.n889 VSUBS 0.24113f
C6710 VDDD.n890 VSUBS 0.070712f
C6711 VDDD.n891 VSUBS 0.089116f
C6712 VDDD.n892 VSUBS 0.251622f
C6713 VDDD.n893 VSUBS 0.251622f
C6714 VDDD.n894 VSUBS 0.251622f
C6715 VDDD.n895 VSUBS 0.3381f
C6716 VDDD.n896 VSUBS 0.056666f
C6717 VDDD.n897 VSUBS 0.049401f
C6718 VDDD.n898 VSUBS 0.251622f
C6719 VDDD.n899 VSUBS 0.251622f
C6720 VDDD.n900 VSUBS 0.052307f
C6721 VDDD.n901 VSUBS 0.089116f
C6722 VDDD.n902 VSUBS 0.089116f
C6723 VDDD.n903 VSUBS 0.251622f
C6724 VDDD.n904 VSUBS 0.251622f
C6725 VDDD.n905 VSUBS 0.251622f
C6726 VDDD.n906 VSUBS 0.250175f
C6727 VDDD.n907 VSUBS 0.067806f
C6728 VDDD.n908 VSUBS 0.074102f
C6729 VDDD.n909 VSUBS 0.251622f
C6730 VDDD.n910 VSUBS 0.251622f
C6731 VDDD.n911 VSUBS 0.149059f
C6732 VDDD.n912 VSUBS 0.062962f
C6733 VDDD.t320 VSUBS 0.306728f
C6734 VDDD.n913 VSUBS 0.427682f
C6735 VDDD.n914 VSUBS 0.188716f
C6736 VDDD.n915 VSUBS 0.251622f
C6737 VDDD.n916 VSUBS 0.251622f
C6738 VDDD.n917 VSUBS 0.521063f
C6739 VDDD.n918 VSUBS 0.032934f
C6740 VDDD.t1137 VSUBS 0.121884f
C6741 VDDD.n919 VSUBS 0.226774f
C6742 VDDD.n920 VSUBS 0.05037f
C6743 VDDD.n921 VSUBS 0.251622f
C6744 VDDD.n922 VSUBS 0.251622f
C6745 VDDD.n923 VSUBS 0.251622f
C6746 VDDD.n924 VSUBS 0.070712f
C6747 VDDD.n925 VSUBS 0.089116f
C6748 VDDD.n926 VSUBS 0.085726f
C6749 VDDD.n927 VSUBS 0.251622f
C6750 VDDD.n928 VSUBS 0.251622f
C6751 VDDD.n929 VSUBS 0.251622f
C6752 VDDD.n930 VSUBS 0.056666f
C6753 VDDD.n931 VSUBS 0.049401f
C6754 VDDD.t902 VSUBS 0.032307f
C6755 VDDD.t155 VSUBS 0.047863f
C6756 VDDD.n932 VSUBS 0.083298f
C6757 VDDD.n933 VSUBS 0.235104f
C6758 VDDD.n934 VSUBS 0.052307f
C6759 VDDD.n935 VSUBS 0.251622f
C6760 VDDD.n936 VSUBS 0.251622f
C6761 VDDD.n937 VSUBS 0.251622f
C6762 VDDD.n938 VSUBS 0.089116f
C6763 VDDD.n939 VSUBS 0.08621f
C6764 VDDD.t1042 VSUBS 0.118653f
C6765 VDDD.n940 VSUBS 0.250175f
C6766 VDDD.n941 VSUBS 0.251622f
C6767 VDDD.n942 VSUBS 0.251622f
C6768 VDDD.n943 VSUBS 0.251622f
C6769 VDDD.n944 VSUBS 0.074102f
C6770 VDDD.t7 VSUBS 0.04923f
C6771 VDDD.t1132 VSUBS 0.04923f
C6772 VDDD.n945 VSUBS 0.102503f
C6773 VDDD.n946 VSUBS 0.305072f
C6774 VDDD.n947 VSUBS 0.062962f
C6775 VDDD.n948 VSUBS 0.149059f
C6776 VDDD.n949 VSUBS 0.188716f
C6777 VDDD.n950 VSUBS 0.251622f
C6778 VDDD.n951 VSUBS 0.057151f
C6779 VDDD.t600 VSUBS 0.337079f
C6780 VDDD.n952 VSUBS 0.521063f
C6781 VDDD.t75 VSUBS 0.121884f
C6782 VDDD.n953 VSUBS 0.226774f
C6783 VDDD.n954 VSUBS 0.032934f
C6784 VDDD.n955 VSUBS 0.251622f
C6785 VDDD.n956 VSUBS 0.251622f
C6786 VDDD.n957 VSUBS 0.251622f
C6787 VDDD.n958 VSUBS 0.24113f
C6788 VDDD.n959 VSUBS 0.070712f
C6789 VDDD.n960 VSUBS 0.089116f
C6790 VDDD.n961 VSUBS 0.251622f
C6791 VDDD.n962 VSUBS 0.251622f
C6792 VDDD.n963 VSUBS 0.251622f
C6793 VDDD.n964 VSUBS 0.3381f
C6794 VDDD.n965 VSUBS 0.056666f
C6795 VDDD.n966 VSUBS 0.049401f
C6796 VDDD.n967 VSUBS 0.251622f
C6797 VDDD.n968 VSUBS 0.251622f
C6798 VDDD.n969 VSUBS 0.052307f
C6799 VDDD.n970 VSUBS 0.089116f
C6800 VDDD.n971 VSUBS 0.089116f
C6801 VDDD.n972 VSUBS 0.251622f
C6802 VDDD.n973 VSUBS 0.251622f
C6803 VDDD.n974 VSUBS 0.251622f
C6804 VDDD.n975 VSUBS 0.250175f
C6805 VDDD.n976 VSUBS 0.067806f
C6806 VDDD.n977 VSUBS 0.074102f
C6807 VDDD.n978 VSUBS 0.251622f
C6808 VDDD.n979 VSUBS 0.251622f
C6809 VDDD.n980 VSUBS 0.149059f
C6810 VDDD.n981 VSUBS 0.072165f
C6811 VDDD.n982 VSUBS 0.06829f
C6812 VDDD.n983 VSUBS 0.188716f
C6813 VDDD.n984 VSUBS 0.251622f
C6814 VDDD.n985 VSUBS 0.251622f
C6815 VDDD.n986 VSUBS 0.049401f
C6816 VDDD.t400 VSUBS 0.076922f
C6817 VDDD.t402 VSUBS 0.076922f
C6818 VDDD.n987 VSUBS 0.168897f
C6819 VDDD.n988 VSUBS 0.406881f
C6820 VDDD.t387 VSUBS 0.076922f
C6821 VDDD.t391 VSUBS 0.076922f
C6822 VDDD.n989 VSUBS 0.168897f
C6823 VDDD.n990 VSUBS 0.362323f
C6824 VDDD.n991 VSUBS 0.049401f
C6825 VDDD.n992 VSUBS 0.251622f
C6826 VDDD.n993 VSUBS 0.251622f
C6827 VDDD.n994 VSUBS 0.251622f
C6828 VDDD.n995 VSUBS 0.045042f
C6829 VDDD.t1455 VSUBS 0.076922f
C6830 VDDD.t268 VSUBS 0.076922f
C6831 VDDD.n996 VSUBS 0.168897f
C6832 VDDD.n997 VSUBS 0.362323f
C6833 VDDD.n998 VSUBS 0.056666f
C6834 VDDD.n999 VSUBS 0.053276f
C6835 VDDD.n1000 VSUBS 0.251622f
C6836 VDDD.n1001 VSUBS 0.251622f
C6837 VDDD.n1002 VSUBS 0.080398f
C6838 VDDD.n1003 VSUBS 0.045527f
C6839 VDDD.n1004 VSUBS 0.207246f
C6840 VDDD.n1005 VSUBS 0.216855f
C6841 VDDD.n1006 VSUBS 6.74323f
C6842 VDDD.n1007 VSUBS 16.1901f
C6843 VDDD.n1008 VSUBS 6.56975f
C6844 VDDD.n1009 VSUBS 0.251622f
C6845 VDDD.t811 VSUBS 0.306728f
C6846 VDDD.t71 VSUBS 0.04923f
C6847 VDDD.t69 VSUBS 0.04923f
C6848 VDDD.n1010 VSUBS 0.102503f
C6849 VDDD.n1011 VSUBS 0.048917f
C6850 VDDD.t815 VSUBS 0.337079f
C6851 VDDD.n1012 VSUBS 0.251622f
C6852 VDDD.n1013 VSUBS 0.089116f
C6853 VDDD.n1014 VSUBS 0.251622f
C6854 VDDD.t878 VSUBS 0.229702f
C6855 VDDD.n1015 VSUBS 0.298385f
C6856 VDDD.n1016 VSUBS 0.251622f
C6857 VDDD.t1419 VSUBS 0.032307f
C6858 VDDD.t1101 VSUBS 0.061025f
C6859 VDDD.n1017 VSUBS 0.096588f
C6860 VDDD.n1018 VSUBS 0.24113f
C6861 VDDD.n1019 VSUBS 0.251622f
C6862 VDDD.t1267 VSUBS 0.117676f
C6863 VDDD.t954 VSUBS 0.12106f
C6864 VDDD.t1393 VSUBS 0.04923f
C6865 VDDD.t1178 VSUBS 0.04923f
C6866 VDDD.n1020 VSUBS 0.102503f
C6867 VDDD.n1021 VSUBS 0.273106f
C6868 VDDD.t347 VSUBS 0.337079f
C6869 VDDD.t940 VSUBS 0.04923f
C6870 VDDD.t67 VSUBS 0.04923f
C6871 VDDD.n1022 VSUBS 0.102503f
C6872 VDDD.n1023 VSUBS 0.273106f
C6873 VDDD.n1024 VSUBS 0.251622f
C6874 VDDD.t1194 VSUBS 0.12106f
C6875 VDDD.t43 VSUBS 0.117676f
C6876 VDDD.t722 VSUBS 0.061025f
C6877 VDDD.t202 VSUBS 0.032307f
C6878 VDDD.n1025 VSUBS 0.096588f
C6879 VDDD.n1026 VSUBS 0.24113f
C6880 VDDD.n1027 VSUBS 0.251622f
C6881 VDDD.t297 VSUBS 0.032307f
C6882 VDDD.t216 VSUBS 0.047863f
C6883 VDDD.n1028 VSUBS 0.083298f
C6884 VDDD.n1029 VSUBS 0.231714f
C6885 VDDD.n1030 VSUBS 0.251622f
C6886 VDDD.t47 VSUBS 0.047863f
C6887 VDDD.t200 VSUBS 0.032307f
C6888 VDDD.n1031 VSUBS 0.083298f
C6889 VDDD.n1032 VSUBS 0.231714f
C6890 VDDD.t1016 VSUBS 0.229702f
C6891 VDDD.n1033 VSUBS 0.251622f
C6892 VDDD.t779 VSUBS 0.032307f
C6893 VDDD.t415 VSUBS 0.061025f
C6894 VDDD.n1034 VSUBS 0.096588f
C6895 VDDD.n1035 VSUBS 0.24113f
C6896 VDDD.n1036 VSUBS 0.251622f
C6897 VDDD.t1389 VSUBS 0.117676f
C6898 VDDD.t1294 VSUBS 0.12106f
C6899 VDDD.t1341 VSUBS 0.04923f
C6900 VDDD.t1149 VSUBS 0.04923f
C6901 VDDD.n1037 VSUBS 0.102503f
C6902 VDDD.n1038 VSUBS 0.273106f
C6903 VDDD.t413 VSUBS 0.337079f
C6904 VDDD.t426 VSUBS 0.04923f
C6905 VDDD.t1437 VSUBS 0.04923f
C6906 VDDD.n1039 VSUBS 0.102503f
C6907 VDDD.n1040 VSUBS 0.273106f
C6908 VDDD.n1041 VSUBS 0.251622f
C6909 VDDD.t744 VSUBS 0.12106f
C6910 VDDD.t796 VSUBS 0.117676f
C6911 VDDD.t839 VSUBS 0.061025f
C6912 VDDD.t1061 VSUBS 0.032307f
C6913 VDDD.n1042 VSUBS 0.096588f
C6914 VDDD.n1043 VSUBS 0.24113f
C6915 VDDD.n1044 VSUBS 0.251622f
C6916 VDDD.t894 VSUBS 0.032307f
C6917 VDDD.t892 VSUBS 0.047863f
C6918 VDDD.n1045 VSUBS 0.083298f
C6919 VDDD.n1046 VSUBS 0.231714f
C6920 VDDD.n1047 VSUBS 0.251622f
C6921 VDDD.t873 VSUBS 0.047863f
C6922 VDDD.t1059 VSUBS 0.032307f
C6923 VDDD.n1048 VSUBS 0.083298f
C6924 VDDD.n1049 VSUBS 0.231714f
C6925 VDDD.t429 VSUBS 0.229702f
C6926 VDDD.n1050 VSUBS 0.251622f
C6927 VDDD.t176 VSUBS 0.032307f
C6928 VDDD.t496 VSUBS 0.061025f
C6929 VDDD.n1051 VSUBS 0.096588f
C6930 VDDD.n1052 VSUBS 0.24113f
C6931 VDDD.n1053 VSUBS 0.251622f
C6932 VDDD.t112 VSUBS 0.117676f
C6933 VDDD.t1078 VSUBS 0.12106f
C6934 VDDD.t1435 VSUBS 0.04923f
C6935 VDDD.t446 VSUBS 0.04923f
C6936 VDDD.n1054 VSUBS 0.102503f
C6937 VDDD.n1055 VSUBS 0.273106f
C6938 VDDD.t1244 VSUBS 0.337079f
C6939 VDDD.t758 VSUBS 0.04923f
C6940 VDDD.t1439 VSUBS 0.04923f
C6941 VDDD.n1056 VSUBS 0.102503f
C6942 VDDD.n1057 VSUBS 0.273106f
C6943 VDDD.n1058 VSUBS 0.251622f
C6944 VDDD.t228 VSUBS 0.12106f
C6945 VDDD.t1279 VSUBS 0.117676f
C6946 VDDD.t306 VSUBS 0.061025f
C6947 VDDD.t178 VSUBS 0.032307f
C6948 VDDD.n1059 VSUBS 0.096588f
C6949 VDDD.n1060 VSUBS 0.24113f
C6950 VDDD.n1061 VSUBS 0.251622f
C6951 VDDD.t1409 VSUBS 0.032307f
C6952 VDDD.t1057 VSUBS 0.047863f
C6953 VDDD.n1062 VSUBS 0.083298f
C6954 VDDD.n1063 VSUBS 0.231714f
C6955 VDDD.n1064 VSUBS 0.251622f
C6956 VDDD.t957 VSUBS 0.047863f
C6957 VDDD.t1321 VSUBS 0.032307f
C6958 VDDD.n1065 VSUBS 0.083298f
C6959 VDDD.n1066 VSUBS 0.231714f
C6960 VDDD.t1334 VSUBS 0.229702f
C6961 VDDD.n1067 VSUBS 0.251622f
C6962 VDDD.t1407 VSUBS 0.032307f
C6963 VDDD.t291 VSUBS 0.061025f
C6964 VDDD.n1068 VSUBS 0.096588f
C6965 VDDD.n1069 VSUBS 0.24113f
C6966 VDDD.n1070 VSUBS 0.251622f
C6967 VDDD.t832 VSUBS 0.117676f
C6968 VDDD.t393 VSUBS 0.12106f
C6969 VDDD.t224 VSUBS 0.04923f
C6970 VDDD.t766 VSUBS 0.04923f
C6971 VDDD.n1071 VSUBS 0.102503f
C6972 VDDD.n1072 VSUBS 0.273106f
C6973 VDDD.t655 VSUBS 0.337079f
C6974 VDDD.t884 VSUBS 0.04923f
C6975 VDDD.t1153 VSUBS 0.04923f
C6976 VDDD.n1073 VSUBS 0.102503f
C6977 VDDD.n1074 VSUBS 0.273106f
C6978 VDDD.n1075 VSUBS 0.251622f
C6979 VDDD.t163 VSUBS 0.12106f
C6980 VDDD.t959 VSUBS 0.117676f
C6981 VDDD.t150 VSUBS 0.061025f
C6982 VDDD.t1411 VSUBS 0.032307f
C6983 VDDD.n1076 VSUBS 0.096588f
C6984 VDDD.n1077 VSUBS 0.24113f
C6985 VDDD.n1078 VSUBS 0.251622f
C6986 VDDD.t373 VSUBS 0.032307f
C6987 VDDD.t120 VSUBS 0.047863f
C6988 VDDD.n1079 VSUBS 0.083298f
C6989 VDDD.n1080 VSUBS 0.231714f
C6990 VDDD.n1081 VSUBS 0.251622f
C6991 VDDD.t39 VSUBS 0.047863f
C6992 VDDD.t1325 VSUBS 0.032307f
C6993 VDDD.n1082 VSUBS 0.083298f
C6994 VDDD.n1083 VSUBS 0.231714f
C6995 VDDD.t570 VSUBS 0.229702f
C6996 VDDD.n1084 VSUBS 0.251622f
C6997 VDDD.t627 VSUBS 0.032307f
C6998 VDDD.t942 VSUBS 0.061025f
C6999 VDDD.n1085 VSUBS 0.096588f
C7000 VDDD.n1086 VSUBS 0.24113f
C7001 VDDD.n1087 VSUBS 0.251622f
C7002 VDDD.t1222 VSUBS 0.117676f
C7003 VDDD.t254 VSUBS 0.12106f
C7004 VDDD.t1391 VSUBS 0.04923f
C7005 VDDD.t168 VSUBS 0.04923f
C7006 VDDD.n1088 VSUBS 0.102503f
C7007 VDDD.n1089 VSUBS 0.273106f
C7008 VDDD.t579 VSUBS 0.337079f
C7009 VDDD.n1090 VSUBS 0.048917f
C7010 VDDD.n1091 VSUBS 0.228374f
C7011 VDDD.n1092 VSUBS 0.123295f
C7012 VDDD.n1093 VSUBS 0.11352f
C7013 VDDD.n1094 VSUBS 0.118956f
C7014 VDDD.n1095 VSUBS 0.427239f
C7015 VDDD.t68 VSUBS 0.588571f
C7016 VDDD.t810 VSUBS 0.677259f
C7017 VDDD.t70 VSUBS 0.677259f
C7018 VDDD.t814 VSUBS 1.79796f
C7019 VDDD.t788 VSUBS 2.08822f
C7020 VDDD.t1124 VSUBS 0.677259f
C7021 VDDD.t1201 VSUBS 0.74176f
C7022 VDDD.t1276 VSUBS 0.870762f
C7023 VDDD.t812 VSUBS 0.798199f
C7024 VDDD.t73 VSUBS 0.677259f
C7025 VDDD.t207 VSUBS 1.02395f
C7026 VDDD.t1179 VSUBS 0.798199f
C7027 VDDD.t1126 VSUBS 0.798199f
C7028 VDDD.t1376 VSUBS 0.782073f
C7029 VDDD.t1344 VSUBS 1.58833f
C7030 VDDD.t203 VSUBS 1.58833f
C7031 VDDD.t877 VSUBS 0.782073f
C7032 VDDD.t993 VSUBS 0.798199f
C7033 VDDD.t72 VSUBS 0.798199f
C7034 VDDD.t698 VSUBS 1.02395f
C7035 VDDD.t1094 VSUBS 0.677259f
C7036 VDDD.t1100 VSUBS 0.798199f
C7037 VDDD.t208 VSUBS 0.870762f
C7038 VDDD.t1418 VSUBS 0.74176f
C7039 VDDD.t1266 VSUBS 0.677259f
C7040 VDDD.t953 VSUBS 2.08822f
C7041 VDDD.t346 VSUBS 1.79796f
C7042 VDDD.t1177 VSUBS 0.677259f
C7043 VDDD.t348 VSUBS 0.677259f
C7044 VDDD.t1392 VSUBS 0.314442f
C7045 VDDD.t66 VSUBS 0.588571f
C7046 VDDD.t280 VSUBS 0.677259f
C7047 VDDD.t939 VSUBS 0.677259f
C7048 VDDD.t719 VSUBS 1.79796f
C7049 VDDD.t1193 VSUBS 2.08822f
C7050 VDDD.t42 VSUBS 0.677259f
C7051 VDDD.t201 VSUBS 0.74176f
C7052 VDDD.t1109 VSUBS 0.870762f
C7053 VDDD.t721 VSUBS 0.798199f
C7054 VDDD.t507 VSUBS 0.677259f
C7055 VDDD.t1083 VSUBS 1.02395f
C7056 VDDD.t629 VSUBS 0.798199f
C7057 VDDD.t215 VSUBS 0.798199f
C7058 VDDD.t164 VSUBS 0.782073f
C7059 VDDD.t296 VSUBS 1.58833f
C7060 VDDD.t199 VSUBS 1.58833f
C7061 VDDD.t1015 VSUBS 0.782073f
C7062 VDDD.t46 VSUBS 0.798199f
C7063 VDDD.t938 VSUBS 0.798199f
C7064 VDDD.t539 VSUBS 1.02395f
C7065 VDDD.t628 VSUBS 0.677259f
C7066 VDDD.t414 VSUBS 0.798199f
C7067 VDDD.t1422 VSUBS 0.870762f
C7068 VDDD.t778 VSUBS 0.74176f
C7069 VDDD.t1388 VSUBS 0.677259f
C7070 VDDD.t1293 VSUBS 2.08822f
C7071 VDDD.t412 VSUBS 1.79796f
C7072 VDDD.t1148 VSUBS 0.677259f
C7073 VDDD.t802 VSUBS 0.677259f
C7074 VDDD.t1340 VSUBS 0.314442f
C7075 VDDD.t1436 VSUBS 0.588571f
C7076 VDDD.t137 VSUBS 0.677259f
C7077 VDDD.t425 VSUBS 0.677259f
C7078 VDDD.t139 VSUBS 1.79796f
C7079 VDDD.t743 VSUBS 2.08822f
C7080 VDDD.t795 VSUBS 0.677259f
C7081 VDDD.t1060 VSUBS 0.74176f
C7082 VDDD.t792 VSUBS 0.870762f
C7083 VDDD.t838 VSUBS 0.798199f
C7084 VDDD.t427 VSUBS 0.677259f
C7085 VDDD.t874 VSUBS 1.02395f
C7086 VDDD.t1374 VSUBS 0.798199f
C7087 VDDD.t891 VSUBS 0.798199f
C7088 VDDD.t762 VSUBS 0.782073f
C7089 VDDD.t893 VSUBS 1.58833f
C7090 VDDD.t1058 VSUBS 1.58833f
C7091 VDDD.t428 VSUBS 0.782073f
C7092 VDDD.t872 VSUBS 0.798199f
C7093 VDDD.t424 VSUBS 0.798199f
C7094 VDDD.t911 VSUBS 1.02395f
C7095 VDDD.t1373 VSUBS 0.677259f
C7096 VDDD.t495 VSUBS 0.798199f
C7097 VDDD.t875 VSUBS 0.870762f
C7098 VDDD.t175 VSUBS 0.74176f
C7099 VDDD.t111 VSUBS 0.677259f
C7100 VDDD.t1077 VSUBS 2.08822f
C7101 VDDD.t1243 VSUBS 1.79796f
C7102 VDDD.t445 VSUBS 0.677259f
C7103 VDDD.t1241 VSUBS 0.677259f
C7104 VDDD.t1434 VSUBS 0.314442f
C7105 VDDD.t1438 VSUBS 0.588571f
C7106 VDDD.t1138 VSUBS 0.677259f
C7107 VDDD.t757 VSUBS 0.677259f
C7108 VDDD.t1140 VSUBS 1.79796f
C7109 VDDD.t227 VSUBS 2.08822f
C7110 VDDD.t1278 VSUBS 0.677259f
C7111 VDDD.t177 VSUBS 0.74176f
C7112 VDDD.t1401 VSUBS 0.870762f
C7113 VDDD.t305 VSUBS 0.798199f
C7114 VDDD.t756 VSUBS 0.677259f
C7115 VDDD.t1192 VSUBS 1.02395f
C7116 VDDD.t867 VSUBS 0.798199f
C7117 VDDD.t1056 VSUBS 0.798199f
C7118 VDDD.t585 VSUBS 0.782073f
C7119 VDDD.t1408 VSUBS 1.58833f
C7120 VDDD.t1320 VSUBS 1.58833f
C7121 VDDD.t1333 VSUBS 0.782073f
C7122 VDDD.t956 VSUBS 0.798199f
C7123 VDDD.t759 VSUBS 0.798199f
C7124 VDDD.t1400 VSUBS 1.02395f
C7125 VDDD.t955 VSUBS 0.677259f
C7126 VDDD.t290 VSUBS 0.798199f
C7127 VDDD.t1191 VSUBS 0.870762f
C7128 VDDD.t1406 VSUBS 0.74176f
C7129 VDDD.t831 VSUBS 0.677259f
C7130 VDDD.t392 VSUBS 2.08822f
C7131 VDDD.t654 VSUBS 1.79796f
C7132 VDDD.t765 VSUBS 0.677259f
C7133 VDDD.t652 VSUBS 0.677259f
C7134 VDDD.t223 VSUBS 0.314442f
C7135 VDDD.t1152 VSUBS 0.588571f
C7136 VDDD.t522 VSUBS 0.677259f
C7137 VDDD.t883 VSUBS 0.677259f
C7138 VDDD.t520 VSUBS 1.79796f
C7139 VDDD.t162 VSUBS 2.08822f
C7140 VDDD.t958 VSUBS 0.677259f
C7141 VDDD.t1410 VSUBS 0.74176f
C7142 VDDD.t952 VSUBS 0.870762f
C7143 VDDD.t149 VSUBS 0.798199f
C7144 VDDD.t325 VSUBS 0.677259f
C7145 VDDD.t1284 VSUBS 1.02395f
C7146 VDDD.t485 VSUBS 0.798199f
C7147 VDDD.t119 VSUBS 0.798199f
C7148 VDDD.t40 VSUBS 0.782073f
C7149 VDDD.t372 VSUBS 1.58833f
C7150 VDDD.t1324 VSUBS 1.58833f
C7151 VDDD.t569 VSUBS 0.782073f
C7152 VDDD.t38 VSUBS 0.798199f
C7153 VDDD.t462 VSUBS 0.798199f
C7154 VDDD.t951 VSUBS 1.02395f
C7155 VDDD.t484 VSUBS 0.677259f
C7156 VDDD.t941 VSUBS 0.798199f
C7157 VDDD.t300 VSUBS 0.870762f
C7158 VDDD.t626 VSUBS 0.74176f
C7159 VDDD.t1221 VSUBS 0.677259f
C7160 VDDD.t253 VSUBS 2.08822f
C7161 VDDD.t578 VSUBS 1.79796f
C7162 VDDD.t167 VSUBS 0.677259f
C7163 VDDD.t576 VSUBS 0.677259f
C7164 VDDD.t1390 VSUBS 0.314442f
C7165 VDDD.t542 VSUBS 2.48328f
C7166 VDDD.t912 VSUBS 1.54802f
C7167 VDDD.t945 VSUBS 1.21745f
C7168 VDDD.n1096 VSUBS 0.864566f
C7169 VDDD.n1097 VSUBS 0.11352f
C7170 VDDD.n1098 VSUBS 0.61245f
C7171 VDDD.n1100 VSUBS 0.11352f
C7172 VDDD.n1101 VSUBS 0.11352f
C7173 VDDD.n1102 VSUBS 0.118956f
C7174 VDDD.n1103 VSUBS 0.559076f
C7175 VDDD.n1104 VSUBS 0.175368f
C7176 VDDD.t1055 VSUBS 0.130341f
C7177 VDDD.t946 VSUBS 0.130341f
C7178 VDDD.n1105 VSUBS 0.541121f
C7179 VDDD.n1106 VSUBS 0.056666f
C7180 VDDD.t656 VSUBS 0.024112f
C7181 VDDD.t913 VSUBS 0.064644f
C7182 VDDD.n1107 VSUBS 0.297902f
C7183 VDDD.t543 VSUBS 0.024112f
C7184 VDDD.t1070 VSUBS 0.064644f
C7185 VDDD.n1108 VSUBS 0.297902f
C7186 VDDD.n1109 VSUBS 0.603939f
C7187 VDDD.n1110 VSUBS 0.052792f
C7188 VDDD.n1111 VSUBS 0.251622f
C7189 VDDD.n1112 VSUBS 0.251622f
C7190 VDDD.n1113 VSUBS 0.188716f
C7191 VDDD.n1114 VSUBS 0.07943f
C7192 VDDD.t577 VSUBS 0.306728f
C7193 VDDD.n1115 VSUBS 0.410246f
C7194 VDDD.n1116 VSUBS 0.084786f
C7195 VDDD.n1117 VSUBS 0.228374f
C7196 VDDD.n1118 VSUBS 0.251622f
C7197 VDDD.n1119 VSUBS 0.506049f
C7198 VDDD.n1120 VSUBS 0.048917f
C7199 VDDD.n1121 VSUBS 0.186431f
C7200 VDDD.n1122 VSUBS 0.165427f
C7201 VDDD.n1123 VSUBS 0.047948f
C7202 VDDD.n1124 VSUBS 0.251622f
C7203 VDDD.n1125 VSUBS 0.251622f
C7204 VDDD.n1126 VSUBS 0.251622f
C7205 VDDD.n1127 VSUBS 0.070712f
C7206 VDDD.n1128 VSUBS 0.089116f
C7207 VDDD.n1129 VSUBS 0.052307f
C7208 VDDD.n1130 VSUBS 0.251622f
C7209 VDDD.n1131 VSUBS 0.251622f
C7210 VDDD.n1132 VSUBS 0.298385f
C7211 VDDD.n1133 VSUBS 0.024216f
C7212 VDDD.t41 VSUBS 0.229702f
C7213 VDDD.n1134 VSUBS 0.298385f
C7214 VDDD.n1135 VSUBS 0.251622f
C7215 VDDD.n1136 VSUBS 0.251622f
C7216 VDDD.n1137 VSUBS 0.052307f
C7217 VDDD.n1138 VSUBS 0.089116f
C7218 VDDD.n1139 VSUBS 0.070712f
C7219 VDDD.n1140 VSUBS 0.251622f
C7220 VDDD.n1141 VSUBS 0.251622f
C7221 VDDD.n1142 VSUBS 0.251622f
C7222 VDDD.n1143 VSUBS 0.047948f
C7223 VDDD.n1144 VSUBS 0.165427f
C7224 VDDD.n1145 VSUBS 0.186431f
C7225 VDDD.n1146 VSUBS 0.048917f
C7226 VDDD.t521 VSUBS 0.337079f
C7227 VDDD.n1147 VSUBS 0.506048f
C7228 VDDD.n1148 VSUBS 0.251622f
C7229 VDDD.n1149 VSUBS 0.251622f
C7230 VDDD.n1150 VSUBS 0.149059f
C7231 VDDD.t523 VSUBS 0.306728f
C7232 VDDD.n1151 VSUBS 0.401528f
C7233 VDDD.t653 VSUBS 0.306728f
C7234 VDDD.n1152 VSUBS 0.401528f
C7235 VDDD.n1153 VSUBS 0.086153f
C7236 VDDD.n1154 VSUBS 0.228374f
C7237 VDDD.n1155 VSUBS 0.251622f
C7238 VDDD.n1156 VSUBS 0.506049f
C7239 VDDD.n1157 VSUBS 0.048917f
C7240 VDDD.n1158 VSUBS 0.186431f
C7241 VDDD.n1159 VSUBS 0.165427f
C7242 VDDD.n1160 VSUBS 0.047948f
C7243 VDDD.n1161 VSUBS 0.251622f
C7244 VDDD.n1162 VSUBS 0.251622f
C7245 VDDD.n1163 VSUBS 0.251622f
C7246 VDDD.n1164 VSUBS 0.070712f
C7247 VDDD.n1165 VSUBS 0.089116f
C7248 VDDD.n1166 VSUBS 0.052307f
C7249 VDDD.n1167 VSUBS 0.251622f
C7250 VDDD.n1168 VSUBS 0.251622f
C7251 VDDD.n1169 VSUBS 0.298385f
C7252 VDDD.n1170 VSUBS 0.024216f
C7253 VDDD.t586 VSUBS 0.229702f
C7254 VDDD.n1171 VSUBS 0.298385f
C7255 VDDD.n1172 VSUBS 0.251622f
C7256 VDDD.n1173 VSUBS 0.251622f
C7257 VDDD.n1174 VSUBS 0.052307f
C7258 VDDD.n1175 VSUBS 0.089116f
C7259 VDDD.n1176 VSUBS 0.070712f
C7260 VDDD.n1177 VSUBS 0.251622f
C7261 VDDD.n1178 VSUBS 0.251622f
C7262 VDDD.n1179 VSUBS 0.251622f
C7263 VDDD.n1180 VSUBS 0.047948f
C7264 VDDD.n1181 VSUBS 0.165427f
C7265 VDDD.n1182 VSUBS 0.186431f
C7266 VDDD.n1183 VSUBS 0.048917f
C7267 VDDD.t1141 VSUBS 0.337079f
C7268 VDDD.n1184 VSUBS 0.506048f
C7269 VDDD.n1185 VSUBS 0.251622f
C7270 VDDD.n1186 VSUBS 0.251622f
C7271 VDDD.n1187 VSUBS 0.149059f
C7272 VDDD.t1139 VSUBS 0.306728f
C7273 VDDD.n1188 VSUBS 0.401528f
C7274 VDDD.t1242 VSUBS 0.306728f
C7275 VDDD.n1189 VSUBS 0.401528f
C7276 VDDD.n1190 VSUBS 0.086153f
C7277 VDDD.n1191 VSUBS 0.228374f
C7278 VDDD.n1192 VSUBS 0.251622f
C7279 VDDD.n1193 VSUBS 0.506049f
C7280 VDDD.n1194 VSUBS 0.048917f
C7281 VDDD.n1195 VSUBS 0.186431f
C7282 VDDD.n1196 VSUBS 0.165427f
C7283 VDDD.n1197 VSUBS 0.047948f
C7284 VDDD.n1198 VSUBS 0.251622f
C7285 VDDD.n1199 VSUBS 0.251622f
C7286 VDDD.n1200 VSUBS 0.251622f
C7287 VDDD.n1201 VSUBS 0.070712f
C7288 VDDD.n1202 VSUBS 0.089116f
C7289 VDDD.n1203 VSUBS 0.052307f
C7290 VDDD.n1204 VSUBS 0.251622f
C7291 VDDD.n1205 VSUBS 0.251622f
C7292 VDDD.n1206 VSUBS 0.298385f
C7293 VDDD.n1207 VSUBS 0.024216f
C7294 VDDD.t763 VSUBS 0.229702f
C7295 VDDD.n1208 VSUBS 0.298385f
C7296 VDDD.n1209 VSUBS 0.251622f
C7297 VDDD.n1210 VSUBS 0.251622f
C7298 VDDD.n1211 VSUBS 0.052307f
C7299 VDDD.n1212 VSUBS 0.089116f
C7300 VDDD.n1213 VSUBS 0.070712f
C7301 VDDD.n1214 VSUBS 0.251622f
C7302 VDDD.n1215 VSUBS 0.251622f
C7303 VDDD.n1216 VSUBS 0.251622f
C7304 VDDD.n1217 VSUBS 0.047948f
C7305 VDDD.n1218 VSUBS 0.165427f
C7306 VDDD.n1219 VSUBS 0.186431f
C7307 VDDD.n1220 VSUBS 0.048917f
C7308 VDDD.t140 VSUBS 0.337079f
C7309 VDDD.n1221 VSUBS 0.506048f
C7310 VDDD.n1222 VSUBS 0.251622f
C7311 VDDD.n1223 VSUBS 0.251622f
C7312 VDDD.n1224 VSUBS 0.149059f
C7313 VDDD.t138 VSUBS 0.306728f
C7314 VDDD.n1225 VSUBS 0.401528f
C7315 VDDD.t803 VSUBS 0.306728f
C7316 VDDD.n1226 VSUBS 0.401528f
C7317 VDDD.n1227 VSUBS 0.086153f
C7318 VDDD.n1228 VSUBS 0.228374f
C7319 VDDD.n1229 VSUBS 0.251622f
C7320 VDDD.n1230 VSUBS 0.506049f
C7321 VDDD.n1231 VSUBS 0.048917f
C7322 VDDD.n1232 VSUBS 0.186431f
C7323 VDDD.n1233 VSUBS 0.165427f
C7324 VDDD.n1234 VSUBS 0.047948f
C7325 VDDD.n1235 VSUBS 0.251622f
C7326 VDDD.n1236 VSUBS 0.251622f
C7327 VDDD.n1237 VSUBS 0.251622f
C7328 VDDD.n1238 VSUBS 0.070712f
C7329 VDDD.n1239 VSUBS 0.089116f
C7330 VDDD.n1240 VSUBS 0.052307f
C7331 VDDD.n1241 VSUBS 0.251622f
C7332 VDDD.n1242 VSUBS 0.251622f
C7333 VDDD.n1243 VSUBS 0.298385f
C7334 VDDD.n1244 VSUBS 0.024216f
C7335 VDDD.t165 VSUBS 0.229702f
C7336 VDDD.n1245 VSUBS 0.298385f
C7337 VDDD.n1246 VSUBS 0.251622f
C7338 VDDD.n1247 VSUBS 0.251622f
C7339 VDDD.n1248 VSUBS 0.052307f
C7340 VDDD.n1249 VSUBS 0.089116f
C7341 VDDD.n1250 VSUBS 0.070712f
C7342 VDDD.n1251 VSUBS 0.251622f
C7343 VDDD.n1252 VSUBS 0.251622f
C7344 VDDD.n1253 VSUBS 0.251622f
C7345 VDDD.n1254 VSUBS 0.047948f
C7346 VDDD.n1255 VSUBS 0.165427f
C7347 VDDD.n1256 VSUBS 0.186431f
C7348 VDDD.n1257 VSUBS 0.048917f
C7349 VDDD.t720 VSUBS 0.337079f
C7350 VDDD.n1258 VSUBS 0.506048f
C7351 VDDD.n1259 VSUBS 0.251622f
C7352 VDDD.n1260 VSUBS 0.251622f
C7353 VDDD.n1261 VSUBS 0.149059f
C7354 VDDD.t281 VSUBS 0.306728f
C7355 VDDD.n1262 VSUBS 0.401528f
C7356 VDDD.t349 VSUBS 0.306728f
C7357 VDDD.n1263 VSUBS 0.401528f
C7358 VDDD.n1264 VSUBS 0.086153f
C7359 VDDD.n1265 VSUBS 0.228374f
C7360 VDDD.n1266 VSUBS 0.251622f
C7361 VDDD.n1267 VSUBS 0.506049f
C7362 VDDD.n1268 VSUBS 0.048917f
C7363 VDDD.n1269 VSUBS 0.186431f
C7364 VDDD.n1270 VSUBS 0.165427f
C7365 VDDD.n1271 VSUBS 0.047948f
C7366 VDDD.n1272 VSUBS 0.251622f
C7367 VDDD.n1273 VSUBS 0.251622f
C7368 VDDD.n1274 VSUBS 0.251622f
C7369 VDDD.n1275 VSUBS 0.070712f
C7370 VDDD.n1276 VSUBS 0.089116f
C7371 VDDD.t994 VSUBS 0.047863f
C7372 VDDD.t204 VSUBS 0.032307f
C7373 VDDD.n1277 VSUBS 0.083298f
C7374 VDDD.n1278 VSUBS 0.231714f
C7375 VDDD.n1279 VSUBS 0.052307f
C7376 VDDD.n1280 VSUBS 0.251622f
C7377 VDDD.n1281 VSUBS 0.251622f
C7378 VDDD.n1282 VSUBS 0.251622f
C7379 VDDD.n1283 VSUBS 0.024216f
C7380 VDDD.t1377 VSUBS 0.229702f
C7381 VDDD.n1284 VSUBS 0.298385f
C7382 VDDD.t1345 VSUBS 0.032307f
C7383 VDDD.t1127 VSUBS 0.047863f
C7384 VDDD.n1285 VSUBS 0.083298f
C7385 VDDD.n1286 VSUBS 0.231714f
C7386 VDDD.n1287 VSUBS 0.052307f
C7387 VDDD.n1288 VSUBS 0.251622f
C7388 VDDD.n1289 VSUBS 0.251622f
C7389 VDDD.n1290 VSUBS 0.251622f
C7390 VDDD.n1291 VSUBS 0.070712f
C7391 VDDD.t813 VSUBS 0.061025f
C7392 VDDD.t1202 VSUBS 0.032307f
C7393 VDDD.n1292 VSUBS 0.096588f
C7394 VDDD.n1293 VSUBS 0.24113f
C7395 VDDD.t1125 VSUBS 0.117676f
C7396 VDDD.t789 VSUBS 0.12106f
C7397 VDDD.n1294 VSUBS 0.186431f
C7398 VDDD.n1295 VSUBS 0.165427f
C7399 VDDD.n1296 VSUBS 0.047948f
C7400 VDDD.n1297 VSUBS 0.251622f
C7401 VDDD.n1298 VSUBS 0.251622f
C7402 VDDD.n1299 VSUBS 0.251622f
C7403 VDDD.n1300 VSUBS 0.506048f
C7404 VDDD.n1301 VSUBS 0.273106f
C7405 VDDD.n1302 VSUBS 0.349221f
C7406 VDDD.n1303 VSUBS 0.149059f
C7407 VDDD.n1304 VSUBS 21.3605f
C7408 VDDD.n1305 VSUBS 12.256599f
C7409 VDDD.n1306 VSUBS 7.0441f
C7410 VDDD.n1307 VSUBS 0.299607f
C7411 VDDD.t365 VSUBS 0.04923f
C7412 VDDD.t1054 VSUBS 0.04923f
C7413 VDDD.n1308 VSUBS 0.102503f
C7414 VDDD.t1204 VSUBS 0.118653f
C7415 VDDD.n1309 VSUBS 0.250175f
C7416 VDDD.n1310 VSUBS 0.251622f
C7417 VDDD.n1311 VSUBS 0.052307f
C7418 VDDD.n1312 VSUBS 0.251622f
C7419 VDDD.n1313 VSUBS 0.251622f
C7420 VDDD.t457 VSUBS 0.229702f
C7421 VDDD.n1314 VSUBS 0.089116f
C7422 VDDD.n1315 VSUBS 0.251622f
C7423 VDDD.t969 VSUBS 0.032307f
C7424 VDDD.t1309 VSUBS 0.061025f
C7425 VDDD.n1316 VSUBS 0.096588f
C7426 VDDD.t1212 VSUBS 0.121884f
C7427 VDDD.n1317 VSUBS 0.226774f
C7428 VDDD.n1318 VSUBS 0.251622f
C7429 VDDD.t230 VSUBS 0.337079f
C7430 VDDD.t1311 VSUBS 0.306728f
C7431 VDDD.n1319 VSUBS 0.427682f
C7432 VDDD.n1320 VSUBS 0.251622f
C7433 VDDD.t31 VSUBS 0.04923f
C7434 VDDD.t1022 VSUBS 0.04923f
C7435 VDDD.n1321 VSUBS 0.102503f
C7436 VDDD.n1322 VSUBS 0.067806f
C7437 VDDD.n1323 VSUBS 0.251622f
C7438 VDDD.t1381 VSUBS 0.118653f
C7439 VDDD.n1324 VSUBS 0.089116f
C7440 VDDD.n1325 VSUBS 0.251622f
C7441 VDDD.t1301 VSUBS 0.032307f
C7442 VDDD.t453 VSUBS 0.047863f
C7443 VDDD.n1326 VSUBS 0.083298f
C7444 VDDD.t882 VSUBS 0.229702f
C7445 VDDD.n1327 VSUBS 0.3381f
C7446 VDDD.n1328 VSUBS 0.251622f
C7447 VDDD.t1273 VSUBS 0.032307f
C7448 VDDD.t1368 VSUBS 0.061025f
C7449 VDDD.n1329 VSUBS 0.096588f
C7450 VDDD.n1330 VSUBS 0.24113f
C7451 VDDD.n1331 VSUBS 0.251622f
C7452 VDDD.t1135 VSUBS 0.121884f
C7453 VDDD.n1332 VSUBS 0.251622f
C7454 VDDD.t1366 VSUBS 0.337079f
C7455 VDDD.t378 VSUBS 0.306728f
C7456 VDDD.n1333 VSUBS 0.427682f
C7457 VDDD.n1334 VSUBS 0.251622f
C7458 VDDD.t122 VSUBS 0.04923f
C7459 VDDD.t828 VSUBS 0.04923f
C7460 VDDD.n1335 VSUBS 0.102503f
C7461 VDDD.n1336 VSUBS 0.067806f
C7462 VDDD.n1337 VSUBS 0.251622f
C7463 VDDD.t643 VSUBS 0.118653f
C7464 VDDD.n1338 VSUBS 0.089116f
C7465 VDDD.n1339 VSUBS 0.251622f
C7466 VDDD.t545 VSUBS 0.032307f
C7467 VDDD.t258 VSUBS 0.047863f
C7468 VDDD.n1340 VSUBS 0.083298f
C7469 VDDD.t214 VSUBS 0.229702f
C7470 VDDD.n1341 VSUBS 0.3381f
C7471 VDDD.n1342 VSUBS 0.251622f
C7472 VDDD.t633 VSUBS 0.032307f
C7473 VDDD.t677 VSUBS 0.061025f
C7474 VDDD.n1343 VSUBS 0.096588f
C7475 VDDD.n1344 VSUBS 0.24113f
C7476 VDDD.n1345 VSUBS 0.251622f
C7477 VDDD.t1106 VSUBS 0.121884f
C7478 VDDD.n1346 VSUBS 0.251622f
C7479 VDDD.t681 VSUBS 0.337079f
C7480 VDDD.t679 VSUBS 0.306728f
C7481 VDDD.n1347 VSUBS 0.427682f
C7482 VDDD.n1348 VSUBS 0.251622f
C7483 VDDD.t368 VSUBS 0.04923f
C7484 VDDD.t1024 VSUBS 0.04923f
C7485 VDDD.n1349 VSUBS 0.102503f
C7486 VDDD.n1350 VSUBS 0.067806f
C7487 VDDD.n1351 VSUBS 0.251622f
C7488 VDDD.t240 VSUBS 0.118653f
C7489 VDDD.n1352 VSUBS 0.089116f
C7490 VDDD.n1353 VSUBS 0.251622f
C7491 VDDD.t1303 VSUBS 0.032307f
C7492 VDDD.t1181 VSUBS 0.047863f
C7493 VDDD.n1354 VSUBS 0.083298f
C7494 VDDD.t518 VSUBS 0.229702f
C7495 VDDD.n1355 VSUBS 0.3381f
C7496 VDDD.n1356 VSUBS 0.251622f
C7497 VDDD.t850 VSUBS 0.032307f
C7498 VDDD.t1087 VSUBS 0.061025f
C7499 VDDD.n1357 VSUBS 0.096588f
C7500 VDDD.n1358 VSUBS 0.24113f
C7501 VDDD.n1359 VSUBS 0.251622f
C7502 VDDD.t1069 VSUBS 0.121884f
C7503 VDDD.n1360 VSUBS 0.251622f
C7504 VDDD.t1089 VSUBS 0.337079f
C7505 VDDD.t1085 VSUBS 0.306728f
C7506 VDDD.n1361 VSUBS 0.427682f
C7507 VDDD.n1362 VSUBS 0.251622f
C7508 VDDD.t1260 VSUBS 0.04923f
C7509 VDDD.t1048 VSUBS 0.04923f
C7510 VDDD.n1363 VSUBS 0.102503f
C7511 VDDD.n1364 VSUBS 0.067806f
C7512 VDDD.n1365 VSUBS 0.251622f
C7513 VDDD.t134 VSUBS 0.118653f
C7514 VDDD.n1366 VSUBS 0.089116f
C7515 VDDD.n1367 VSUBS 0.251622f
C7516 VDDD.t908 VSUBS 0.032307f
C7517 VDDD.t449 VSUBS 0.047863f
C7518 VDDD.n1368 VSUBS 0.083298f
C7519 VDDD.t455 VSUBS 0.229702f
C7520 VDDD.n1369 VSUBS 0.3381f
C7521 VDDD.n1370 VSUBS 0.251622f
C7522 VDDD.t516 VSUBS 0.032307f
C7523 VDDD.t1232 VSUBS 0.061025f
C7524 VDDD.n1371 VSUBS 0.096588f
C7525 VDDD.n1372 VSUBS 0.24113f
C7526 VDDD.n1373 VSUBS 0.251622f
C7527 VDDD.t1240 VSUBS 0.121884f
C7528 VDDD.n1374 VSUBS 0.251622f
C7529 VDDD.t1230 VSUBS 0.337079f
C7530 VDDD.t322 VSUBS 0.306728f
C7531 VDDD.n1375 VSUBS 0.366172f
C7532 VDDD.t1052 VSUBS 0.04923f
C7533 VDDD.t441 VSUBS 0.04923f
C7534 VDDD.n1376 VSUBS 0.102503f
C7535 VDDD.n1377 VSUBS 0.228374f
C7536 VDDD.n1378 VSUBS 0.067806f
C7537 VDDD.n1379 VSUBS 0.251622f
C7538 VDDD.t534 VSUBS 0.118653f
C7539 VDDD.n1380 VSUBS 0.089116f
C7540 VDDD.n1381 VSUBS 0.251622f
C7541 VDDD.t329 VSUBS 0.047863f
C7542 VDDD.t266 VSUBS 0.032307f
C7543 VDDD.n1382 VSUBS 0.083298f
C7544 VDDD.t95 VSUBS 0.229702f
C7545 VDDD.n1383 VSUBS 0.3381f
C7546 VDDD.n1384 VSUBS 0.251622f
C7547 VDDD.t967 VSUBS 0.061025f
C7548 VDDD.t971 VSUBS 0.032307f
C7549 VDDD.n1385 VSUBS 0.096588f
C7550 VDDD.n1386 VSUBS 0.24113f
C7551 VDDD.n1387 VSUBS 0.251622f
C7552 VDDD.t1397 VSUBS 0.121884f
C7553 VDDD.t963 VSUBS 0.337079f
C7554 VDDD.n1388 VSUBS 0.251622f
C7555 VDDD.t965 VSUBS 0.306728f
C7556 VDDD.n1389 VSUBS 0.427682f
C7557 VDDD.t830 VSUBS 0.04923f
C7558 VDDD.t1426 VSUBS 0.04923f
C7559 VDDD.n1390 VSUBS 0.102503f
C7560 VDDD.n1391 VSUBS 0.228374f
C7561 VDDD.n1392 VSUBS 0.067806f
C7562 VDDD.n1393 VSUBS 0.251622f
C7563 VDDD.t1 VSUBS 0.118653f
C7564 VDDD.n1394 VSUBS 0.089116f
C7565 VDDD.n1395 VSUBS 0.251622f
C7566 VDDD.t651 VSUBS 0.047863f
C7567 VDDD.t483 VSUBS 0.032307f
C7568 VDDD.n1396 VSUBS 0.083298f
C7569 VDDD.t1234 VSUBS 0.229702f
C7570 VDDD.n1397 VSUBS 0.3381f
C7571 VDDD.n1398 VSUBS 0.251622f
C7572 VDDD.t1044 VSUBS 0.061025f
C7573 VDDD.t1072 VSUBS 0.032307f
C7574 VDDD.n1399 VSUBS 0.096588f
C7575 VDDD.n1400 VSUBS 0.24113f
C7576 VDDD.n1401 VSUBS 0.251622f
C7577 VDDD.t800 VSUBS 0.121884f
C7578 VDDD.t1046 VSUBS 0.337079f
C7579 VDDD.n1402 VSUBS 0.251622f
C7580 VDDD.t1076 VSUBS 0.306728f
C7581 VDDD.n1403 VSUBS 0.427682f
C7582 VDDD.t1115 VSUBS 0.04923f
C7583 VDDD.t246 VSUBS 0.04923f
C7584 VDDD.n1404 VSUBS 0.102503f
C7585 VDDD.n1405 VSUBS 0.228374f
C7586 VDDD.n1406 VSUBS 0.067806f
C7587 VDDD.n1407 VSUBS 0.251622f
C7588 VDDD.t1290 VSUBS 0.118653f
C7589 VDDD.n1408 VSUBS 0.089116f
C7590 VDDD.n1409 VSUBS 0.251622f
C7591 VDDD.t1098 VSUBS 0.047863f
C7592 VDDD.t314 VSUBS 0.032307f
C7593 VDDD.n1410 VSUBS 0.083298f
C7594 VDDD.t361 VSUBS 0.229702f
C7595 VDDD.n1411 VSUBS 0.3381f
C7596 VDDD.n1412 VSUBS 0.251622f
C7597 VDDD.t1254 VSUBS 0.061025f
C7598 VDDD.t618 VSUBS 0.032307f
C7599 VDDD.n1413 VSUBS 0.096588f
C7600 VDDD.n1414 VSUBS 0.24113f
C7601 VDDD.n1415 VSUBS 0.251622f
C7602 VDDD.t1296 VSUBS 0.121884f
C7603 VDDD.t1250 VSUBS 0.337079f
C7604 VDDD.n1416 VSUBS 0.251622f
C7605 VDDD.t1252 VSUBS 0.306728f
C7606 VDDD.n1417 VSUBS 0.427682f
C7607 VDDD.t826 VSUBS 0.04923f
C7608 VDDD.t1006 VSUBS 0.04923f
C7609 VDDD.n1418 VSUBS 0.102503f
C7610 VDDD.n1419 VSUBS 0.228374f
C7611 VDDD.n1420 VSUBS 0.067806f
C7612 VDDD.n1421 VSUBS 0.251622f
C7613 VDDD.t670 VSUBS 0.118653f
C7614 VDDD.n1422 VSUBS 0.089116f
C7615 VDDD.n1423 VSUBS 0.251622f
C7616 VDDD.t641 VSUBS 0.047863f
C7617 VDDD.t1271 VSUBS 0.032307f
C7618 VDDD.n1424 VSUBS 0.083298f
C7619 VDDD.t468 VSUBS 0.229702f
C7620 VDDD.n1425 VSUBS 0.3381f
C7621 VDDD.n1426 VSUBS 0.251622f
C7622 VDDD.t1265 VSUBS 0.061025f
C7623 VDDD.t116 VSUBS 0.032307f
C7624 VDDD.n1427 VSUBS 0.096588f
C7625 VDDD.n1428 VSUBS 0.24113f
C7626 VDDD.n1429 VSUBS 0.251622f
C7627 VDDD.t222 VSUBS 0.121884f
C7628 VDDD.t1262 VSUBS 0.337079f
C7629 VDDD.n1430 VSUBS 0.251622f
C7630 VDDD.t1332 VSUBS 0.306728f
C7631 VDDD.n1431 VSUBS 0.427682f
C7632 VDDD.t694 VSUBS 0.04923f
C7633 VDDD.t597 VSUBS 0.04923f
C7634 VDDD.n1432 VSUBS 0.102503f
C7635 VDDD.n1433 VSUBS 0.228374f
C7636 VDDD.n1434 VSUBS 0.067806f
C7637 VDDD.n1435 VSUBS 0.251622f
C7638 VDDD.t83 VSUBS 0.118653f
C7639 VDDD.n1436 VSUBS 0.089116f
C7640 VDDD.n1437 VSUBS 0.251622f
C7641 VDDD.t880 VSUBS 0.047863f
C7642 VDDD.t822 VSUBS 0.032307f
C7643 VDDD.n1438 VSUBS 0.083298f
C7644 VDDD.t1327 VSUBS 0.229702f
C7645 VDDD.n1439 VSUBS 0.3381f
C7646 VDDD.n1440 VSUBS 0.251622f
C7647 VDDD.t1143 VSUBS 0.061025f
C7648 VDDD.t170 VSUBS 0.032307f
C7649 VDDD.n1441 VSUBS 0.096588f
C7650 VDDD.n1442 VSUBS 0.24113f
C7651 VDDD.n1443 VSUBS 0.251622f
C7652 VDDD.t476 VSUBS 0.121884f
C7653 VDDD.t89 VSUBS 0.337079f
C7654 VDDD.n1444 VSUBS 0.251622f
C7655 VDDD.t87 VSUBS 0.306728f
C7656 VDDD.n1445 VSUBS 0.427198f
C7657 VDDD.t980 VSUBS 0.076922f
C7658 VDDD.t1421 VSUBS 0.076922f
C7659 VDDD.n1446 VSUBS 0.165125f
C7660 VDDD.n1447 VSUBS 0.080398f
C7661 VDDD.n1448 VSUBS 0.251622f
C7662 VDDD.t423 VSUBS 0.076922f
C7663 VDDD.t1091 VSUBS 0.076922f
C7664 VDDD.n1449 VSUBS 0.165125f
C7665 VDDD.n1450 VSUBS 0.188262f
C7666 VDDD.t1441 VSUBS 0.076922f
C7667 VDDD.t1093 VSUBS 0.076922f
C7668 VDDD.n1451 VSUBS 0.168897f
C7669 VDDD.n1452 VSUBS 0.048917f
C7670 VDDD.n1453 VSUBS 0.251622f
C7671 VDDD.t1447 VSUBS 0.076922f
C7672 VDDD.t1443 VSUBS 0.076922f
C7673 VDDD.n1454 VSUBS 0.168897f
C7674 VDDD.n1455 VSUBS 0.362323f
C7675 VDDD.t672 VSUBS 0.076922f
C7676 VDDD.t1449 VSUBS 0.076922f
C7677 VDDD.n1456 VSUBS 0.168897f
C7678 VDDD.t1445 VSUBS 0.307526f
C7679 VDDD.n1457 VSUBS 0.565214f
C7680 VDDD.n1458 VSUBS 0.294184f
C7681 VDDD.n1459 VSUBS 0.302652f
C7682 VDDD.n1460 VSUBS 0.049401f
C7683 VDDD.n1461 VSUBS 0.406881f
C7684 VDDD.n1462 VSUBS 0.049401f
C7685 VDDD.n1463 VSUBS 0.251622f
C7686 VDDD.n1464 VSUBS 0.251622f
C7687 VDDD.n1465 VSUBS 0.251622f
C7688 VDDD.n1466 VSUBS 0.045042f
C7689 VDDD.n1467 VSUBS 0.362323f
C7690 VDDD.n1468 VSUBS 0.056666f
C7691 VDDD.n1469 VSUBS 0.053276f
C7692 VDDD.n1470 VSUBS 0.251622f
C7693 VDDD.n1471 VSUBS 0.251622f
C7694 VDDD.n1472 VSUBS 0.227007f
C7695 VDDD.n1473 VSUBS 0.045527f
C7696 VDDD.n1474 VSUBS 0.188262f
C7697 VDDD.n1475 VSUBS 0.078461f
C7698 VDDD.n1476 VSUBS 0.086153f
C7699 VDDD.n1477 VSUBS 0.188716f
C7700 VDDD.n1478 VSUBS 0.251622f
C7701 VDDD.n1479 VSUBS 0.057151f
C7702 VDDD.n1480 VSUBS 0.521063f
C7703 VDDD.n1481 VSUBS 0.032934f
C7704 VDDD.n1482 VSUBS 0.226774f
C7705 VDDD.n1483 VSUBS 0.05037f
C7706 VDDD.n1484 VSUBS 0.251622f
C7707 VDDD.n1485 VSUBS 0.251622f
C7708 VDDD.n1486 VSUBS 0.251622f
C7709 VDDD.n1487 VSUBS 0.070712f
C7710 VDDD.n1488 VSUBS 0.089116f
C7711 VDDD.n1489 VSUBS 0.085726f
C7712 VDDD.n1490 VSUBS 0.251622f
C7713 VDDD.n1491 VSUBS 0.251622f
C7714 VDDD.n1492 VSUBS 0.251622f
C7715 VDDD.n1493 VSUBS 0.056666f
C7716 VDDD.n1494 VSUBS 0.049401f
C7717 VDDD.n1495 VSUBS 0.235104f
C7718 VDDD.n1496 VSUBS 0.052307f
C7719 VDDD.n1497 VSUBS 0.251622f
C7720 VDDD.n1498 VSUBS 0.251622f
C7721 VDDD.n1499 VSUBS 0.251622f
C7722 VDDD.n1500 VSUBS 0.089116f
C7723 VDDD.n1501 VSUBS 0.08621f
C7724 VDDD.n1502 VSUBS 0.250175f
C7725 VDDD.n1503 VSUBS 0.251622f
C7726 VDDD.n1504 VSUBS 0.251622f
C7727 VDDD.n1505 VSUBS 0.251622f
C7728 VDDD.n1506 VSUBS 0.074102f
C7729 VDDD.n1507 VSUBS 0.305072f
C7730 VDDD.n1508 VSUBS 0.062962f
C7731 VDDD.n1509 VSUBS 0.086153f
C7732 VDDD.n1510 VSUBS 0.188716f
C7733 VDDD.n1511 VSUBS 0.251622f
C7734 VDDD.n1512 VSUBS 0.057151f
C7735 VDDD.n1513 VSUBS 0.521063f
C7736 VDDD.n1514 VSUBS 0.032934f
C7737 VDDD.n1515 VSUBS 0.226774f
C7738 VDDD.n1516 VSUBS 0.05037f
C7739 VDDD.n1517 VSUBS 0.251622f
C7740 VDDD.n1518 VSUBS 0.251622f
C7741 VDDD.n1519 VSUBS 0.251622f
C7742 VDDD.n1520 VSUBS 0.070712f
C7743 VDDD.n1521 VSUBS 0.089116f
C7744 VDDD.n1522 VSUBS 0.085726f
C7745 VDDD.n1523 VSUBS 0.251622f
C7746 VDDD.n1524 VSUBS 0.251622f
C7747 VDDD.n1525 VSUBS 0.251622f
C7748 VDDD.n1526 VSUBS 0.056666f
C7749 VDDD.n1527 VSUBS 0.049401f
C7750 VDDD.n1528 VSUBS 0.235104f
C7751 VDDD.n1529 VSUBS 0.052307f
C7752 VDDD.n1530 VSUBS 0.251622f
C7753 VDDD.n1531 VSUBS 0.251622f
C7754 VDDD.n1532 VSUBS 0.251622f
C7755 VDDD.n1533 VSUBS 0.089116f
C7756 VDDD.n1534 VSUBS 0.08621f
C7757 VDDD.n1535 VSUBS 0.250175f
C7758 VDDD.n1536 VSUBS 0.251622f
C7759 VDDD.n1537 VSUBS 0.251622f
C7760 VDDD.n1538 VSUBS 0.251622f
C7761 VDDD.n1539 VSUBS 0.074102f
C7762 VDDD.n1540 VSUBS 0.305072f
C7763 VDDD.n1541 VSUBS 0.062962f
C7764 VDDD.n1542 VSUBS 0.086153f
C7765 VDDD.n1543 VSUBS 0.188716f
C7766 VDDD.n1544 VSUBS 0.251622f
C7767 VDDD.n1545 VSUBS 0.057151f
C7768 VDDD.n1546 VSUBS 0.521063f
C7769 VDDD.n1547 VSUBS 0.032934f
C7770 VDDD.n1548 VSUBS 0.226774f
C7771 VDDD.n1549 VSUBS 0.05037f
C7772 VDDD.n1550 VSUBS 0.251622f
C7773 VDDD.n1551 VSUBS 0.251622f
C7774 VDDD.n1552 VSUBS 0.251622f
C7775 VDDD.n1553 VSUBS 0.070712f
C7776 VDDD.n1554 VSUBS 0.089116f
C7777 VDDD.n1555 VSUBS 0.085726f
C7778 VDDD.n1556 VSUBS 0.251622f
C7779 VDDD.n1557 VSUBS 0.251622f
C7780 VDDD.n1558 VSUBS 0.251622f
C7781 VDDD.n1559 VSUBS 0.056666f
C7782 VDDD.n1560 VSUBS 0.049401f
C7783 VDDD.n1561 VSUBS 0.235104f
C7784 VDDD.n1562 VSUBS 0.052307f
C7785 VDDD.n1563 VSUBS 0.251622f
C7786 VDDD.n1564 VSUBS 0.251622f
C7787 VDDD.n1565 VSUBS 0.251622f
C7788 VDDD.n1566 VSUBS 0.089116f
C7789 VDDD.n1567 VSUBS 0.08621f
C7790 VDDD.n1568 VSUBS 0.250175f
C7791 VDDD.n1569 VSUBS 0.251622f
C7792 VDDD.n1570 VSUBS 0.251622f
C7793 VDDD.n1571 VSUBS 0.251622f
C7794 VDDD.n1572 VSUBS 0.074102f
C7795 VDDD.n1573 VSUBS 0.305072f
C7796 VDDD.n1574 VSUBS 0.062962f
C7797 VDDD.n1575 VSUBS 0.086153f
C7798 VDDD.n1576 VSUBS 0.188716f
C7799 VDDD.n1577 VSUBS 0.251622f
C7800 VDDD.n1578 VSUBS 0.057151f
C7801 VDDD.n1579 VSUBS 0.521063f
C7802 VDDD.n1580 VSUBS 0.032934f
C7803 VDDD.n1581 VSUBS 0.226774f
C7804 VDDD.n1582 VSUBS 0.05037f
C7805 VDDD.n1583 VSUBS 0.251622f
C7806 VDDD.n1584 VSUBS 0.251622f
C7807 VDDD.n1585 VSUBS 0.251622f
C7808 VDDD.n1586 VSUBS 0.070712f
C7809 VDDD.n1587 VSUBS 0.089116f
C7810 VDDD.n1588 VSUBS 0.085726f
C7811 VDDD.n1589 VSUBS 0.251622f
C7812 VDDD.n1590 VSUBS 0.251622f
C7813 VDDD.n1591 VSUBS 0.251622f
C7814 VDDD.n1592 VSUBS 0.056666f
C7815 VDDD.n1593 VSUBS 0.049401f
C7816 VDDD.n1594 VSUBS 0.235104f
C7817 VDDD.n1595 VSUBS 0.052307f
C7818 VDDD.n1596 VSUBS 0.251622f
C7819 VDDD.n1597 VSUBS 0.251622f
C7820 VDDD.n1598 VSUBS 0.251622f
C7821 VDDD.n1599 VSUBS 0.089116f
C7822 VDDD.n1600 VSUBS 0.08621f
C7823 VDDD.n1601 VSUBS 0.250175f
C7824 VDDD.n1602 VSUBS 0.251622f
C7825 VDDD.n1603 VSUBS 0.251622f
C7826 VDDD.n1604 VSUBS 0.251622f
C7827 VDDD.n1605 VSUBS 0.074102f
C7828 VDDD.n1606 VSUBS 0.305072f
C7829 VDDD.n1607 VSUBS 0.062962f
C7830 VDDD.n1608 VSUBS 0.086153f
C7831 VDDD.n1609 VSUBS 0.188716f
C7832 VDDD.n1610 VSUBS 0.251622f
C7833 VDDD.n1611 VSUBS 0.057151f
C7834 VDDD.n1612 VSUBS 0.521063f
C7835 VDDD.n1613 VSUBS 0.032934f
C7836 VDDD.n1614 VSUBS 0.226774f
C7837 VDDD.n1615 VSUBS 0.05037f
C7838 VDDD.n1616 VSUBS 0.251622f
C7839 VDDD.n1617 VSUBS 0.251622f
C7840 VDDD.n1618 VSUBS 0.251622f
C7841 VDDD.n1619 VSUBS 0.070712f
C7842 VDDD.n1620 VSUBS 0.089116f
C7843 VDDD.n1621 VSUBS 0.085726f
C7844 VDDD.n1622 VSUBS 0.251622f
C7845 VDDD.n1623 VSUBS 0.251622f
C7846 VDDD.n1624 VSUBS 0.251622f
C7847 VDDD.n1625 VSUBS 0.056666f
C7848 VDDD.n1626 VSUBS 0.049401f
C7849 VDDD.n1627 VSUBS 0.235104f
C7850 VDDD.n1628 VSUBS 0.052307f
C7851 VDDD.n1629 VSUBS 0.251622f
C7852 VDDD.n1630 VSUBS 0.251622f
C7853 VDDD.n1631 VSUBS 0.251622f
C7854 VDDD.n1632 VSUBS 0.089116f
C7855 VDDD.n1633 VSUBS 0.08621f
C7856 VDDD.n1634 VSUBS 0.250175f
C7857 VDDD.n1635 VSUBS 0.251622f
C7858 VDDD.n1636 VSUBS 0.251622f
C7859 VDDD.n1637 VSUBS 0.251622f
C7860 VDDD.n1638 VSUBS 0.074102f
C7861 VDDD.n1639 VSUBS 0.326891f
C7862 VDDD.n1640 VSUBS 0.263934f
C7863 VDDD.n1641 VSUBS 0.670393f
C7864 VDDD.n1642 VSUBS 0.118956f
C7865 VDDD.n1643 VSUBS 0.11352f
C7866 VDDD.n1644 VSUBS 0.11352f
C7867 VDDD.n1645 VSUBS 0.11352f
C7868 VDDD.n1646 VSUBS 0.427239f
C7869 VDDD.n1648 VSUBS 0.61245f
C7870 VDDD.t1444 VSUBS 2.28631f
C7871 VDDD.t1448 VSUBS 0.768199f
C7872 VDDD.t671 VSUBS 0.768199f
C7873 VDDD.t1442 VSUBS 0.768199f
C7874 VDDD.t1446 VSUBS 0.768199f
C7875 VDDD.t1092 VSUBS 0.768199f
C7876 VDDD.t1440 VSUBS 0.768199f
C7877 VDDD.t1090 VSUBS 0.768199f
C7878 VDDD.t422 VSUBS 0.768199f
C7879 VDDD.t1420 VSUBS 0.768199f
C7880 VDDD.t979 VSUBS 0.521278f
C7881 VDDD.t86 VSUBS 1.13857f
C7882 VDDD.t88 VSUBS 1.3672f
C7883 VDDD.t475 VSUBS 1.3672f
C7884 VDDD.t169 VSUBS 0.877942f
C7885 VDDD.t1142 VSUBS 0.877942f
C7886 VDDD.t1163 VSUBS 0.777344f
C7887 VDDD.t1156 VSUBS 0.845919f
C7888 VDDD.t1326 VSUBS 1.35346f
C7889 VDDD.t821 VSUBS 1.34432f
C7890 VDDD.t879 VSUBS 1.08369f
C7891 VDDD.t598 VSUBS 1.09284f
C7892 VDDD.t1164 VSUBS 0.873355f
C7893 VDDD.t82 VSUBS 1.64155f
C7894 VDDD.t596 VSUBS 1.60497f
C7895 VDDD.t693 VSUBS 0.525836f
C7896 VDDD.t1331 VSUBS 1.13857f
C7897 VDDD.t1261 VSUBS 1.3672f
C7898 VDDD.t221 VSUBS 1.3672f
C7899 VDDD.t115 VSUBS 0.877942f
C7900 VDDD.t1264 VSUBS 0.877942f
C7901 VDDD.t837 VSUBS 0.777344f
C7902 VDDD.t363 VSUBS 0.845919f
C7903 VDDD.t467 VSUBS 1.35346f
C7904 VDDD.t1270 VSUBS 1.34432f
C7905 VDDD.t640 VSUBS 1.08369f
C7906 VDDD.t362 VSUBS 1.09284f
C7907 VDDD.t842 VSUBS 0.873355f
C7908 VDDD.t669 VSUBS 1.64155f
C7909 VDDD.t1005 VSUBS 1.60497f
C7910 VDDD.t825 VSUBS 0.525836f
C7911 VDDD.t1251 VSUBS 1.13857f
C7912 VDDD.t1249 VSUBS 1.3672f
C7913 VDDD.t1295 VSUBS 1.3672f
C7914 VDDD.t617 VSUBS 0.877942f
C7915 VDDD.t1253 VSUBS 0.877942f
C7916 VDDD.t986 VSUBS 0.777344f
C7917 VDDD.t247 VSUBS 0.845919f
C7918 VDDD.t360 VSUBS 1.35346f
C7919 VDDD.t313 VSUBS 1.34432f
C7920 VDDD.t1097 VSUBS 1.08369f
C7921 VDDD.t1263 VSUBS 1.09284f
C7922 VDDD.t985 VSUBS 0.873355f
C7923 VDDD.t1289 VSUBS 1.64155f
C7924 VDDD.t245 VSUBS 1.60497f
C7925 VDDD.t1114 VSUBS 0.525836f
C7926 VDDD.t1075 VSUBS 1.13857f
C7927 VDDD.t1045 VSUBS 1.3672f
C7928 VDDD.t799 VSUBS 1.3672f
C7929 VDDD.t1071 VSUBS 0.877942f
C7930 VDDD.t1043 VSUBS 0.877942f
C7931 VDDD.t1095 VSUBS 0.777344f
C7932 VDDD.t697 VSUBS 0.845919f
C7933 VDDD.t1233 VSUBS 1.35346f
C7934 VDDD.t482 VSUBS 1.34432f
C7935 VDDD.t650 VSUBS 1.08369f
C7936 VDDD.t1427 VSUBS 1.09284f
C7937 VDDD.t1096 VSUBS 0.873355f
C7938 VDDD.t0 VSUBS 1.64155f
C7939 VDDD.t1425 VSUBS 1.60497f
C7940 VDDD.t829 VSUBS 0.525836f
C7941 VDDD.t964 VSUBS 1.13857f
C7942 VDDD.t962 VSUBS 1.3672f
C7943 VDDD.t1396 VSUBS 1.3672f
C7944 VDDD.t970 VSUBS 0.877942f
C7945 VDDD.t966 VSUBS 0.877942f
C7946 VDDD.t840 VSUBS 0.777344f
C7947 VDDD.t1329 VSUBS 0.845919f
C7948 VDDD.t94 VSUBS 1.35346f
C7949 VDDD.t265 VSUBS 1.34432f
C7950 VDDD.t328 VSUBS 1.08369f
C7951 VDDD.t1328 VSUBS 1.09284f
C7952 VDDD.t841 VSUBS 0.873355f
C7953 VDDD.t533 VSUBS 1.64155f
C7954 VDDD.t440 VSUBS 1.60497f
C7955 VDDD.t1051 VSUBS 0.525836f
C7956 VDDD.n1649 VSUBS 0.726149f
C7957 VDDD.n1650 VSUBS 0.118956f
C7958 VDDD.n1651 VSUBS 0.118956f
C7959 VDDD.n1652 VSUBS 0.11352f
C7960 VDDD.n1653 VSUBS 1.47234f
C7961 VDDD.n1654 VSUBS 1.47738f
C7962 VDDD.n1655 VSUBS 0.118956f
C7963 VDDD.n1656 VSUBS 0.11352f
C7964 VDDD.n1657 VSUBS 0.11352f
C7965 VDDD.n1658 VSUBS 0.11352f
C7966 VDDD.n1659 VSUBS 0.427239f
C7967 VDDD.n1661 VSUBS 0.61245f
C7968 VDDD.t1053 VSUBS 0.681305f
C7969 VDDD.t364 VSUBS 1.60497f
C7970 VDDD.t1203 VSUBS 1.64155f
C7971 VDDD.t1099 VSUBS 0.873355f
C7972 VDDD.t26 VSUBS 1.09284f
C7973 VDDD.t1027 VSUBS 1.08369f
C7974 VDDD.t636 VSUBS 1.34432f
C7975 VDDD.t456 VSUBS 1.35346f
C7976 VDDD.t25 VSUBS 0.845919f
C7977 VDDD.t930 VSUBS 0.777344f
C7978 VDDD.t1308 VSUBS 0.877942f
C7979 VDDD.t968 VSUBS 0.877942f
C7980 VDDD.t1211 VSUBS 1.3672f
C7981 VDDD.t229 VSUBS 1.3672f
C7982 VDDD.t1310 VSUBS 0.983097f
C7983 VDDD.t1021 VSUBS 0.681305f
C7984 VDDD.t30 VSUBS 1.60497f
C7985 VDDD.t1380 VSUBS 1.64155f
C7986 VDDD.t1339 VSUBS 0.873355f
C7987 VDDD.t791 VSUBS 1.09284f
C7988 VDDD.t452 VSUBS 1.08369f
C7989 VDDD.t1300 VSUBS 1.34432f
C7990 VDDD.t881 VSUBS 1.35346f
C7991 VDDD.t29 VSUBS 0.845919f
C7992 VDDD.t690 VSUBS 0.777344f
C7993 VDDD.t1367 VSUBS 0.877942f
C7994 VDDD.t1272 VSUBS 0.877942f
C7995 VDDD.t1134 VSUBS 1.3672f
C7996 VDDD.t1365 VSUBS 1.3672f
C7997 VDDD.t377 VSUBS 0.983097f
C7998 VDDD.t827 VSUBS 0.681305f
C7999 VDDD.t121 VSUBS 1.60497f
C8000 VDDD.t642 VSUBS 1.64155f
C8001 VDDD.t943 VSUBS 0.873355f
C8002 VDDD.t123 VSUBS 1.09284f
C8003 VDDD.t257 VSUBS 1.08369f
C8004 VDDD.t544 VSUBS 1.34432f
C8005 VDDD.t213 VSUBS 1.35346f
C8006 VDDD.t571 VSUBS 0.845919f
C8007 VDDD.t944 VSUBS 0.777344f
C8008 VDDD.t676 VSUBS 0.877942f
C8009 VDDD.t632 VSUBS 0.877942f
C8010 VDDD.t1105 VSUBS 1.3672f
C8011 VDDD.t680 VSUBS 1.3672f
C8012 VDDD.t678 VSUBS 0.983097f
C8013 VDDD.t1023 VSUBS 0.681305f
C8014 VDDD.t367 VSUBS 1.60497f
C8015 VDDD.t239 VSUBS 1.64155f
C8016 VDDD.t60 VSUBS 0.873355f
C8017 VDDD.t369 VSUBS 1.09284f
C8018 VDDD.t1180 VSUBS 1.08369f
C8019 VDDD.t1302 VSUBS 1.34432f
C8020 VDDD.t517 VSUBS 1.35346f
C8021 VDDD.t366 VSUBS 0.845919f
C8022 VDDD.t664 VSUBS 0.777344f
C8023 VDDD.t1086 VSUBS 0.877942f
C8024 VDDD.t849 VSUBS 0.877942f
C8025 VDDD.t1068 VSUBS 1.3672f
C8026 VDDD.t1088 VSUBS 1.3672f
C8027 VDDD.t1084 VSUBS 0.983097f
C8028 VDDD.t1047 VSUBS 0.681305f
C8029 VDDD.t1259 VSUBS 1.60497f
C8030 VDDD.t133 VSUBS 1.64155f
C8031 VDDD.t143 VSUBS 0.873355f
C8032 VDDD.t504 VSUBS 1.09284f
C8033 VDDD.t448 VSUBS 1.08369f
C8034 VDDD.t907 VSUBS 1.34432f
C8035 VDDD.t454 VSUBS 1.35346f
C8036 VDDD.t623 VSUBS 0.845919f
C8037 VDDD.t1208 VSUBS 0.777344f
C8038 VDDD.t1231 VSUBS 0.877942f
C8039 VDDD.t515 VSUBS 0.877942f
C8040 VDDD.t1239 VSUBS 1.3672f
C8041 VDDD.t1229 VSUBS 1.3672f
C8042 VDDD.t321 VSUBS 1.30317f
C8043 VDDD.n1662 VSUBS 0.889235f
C8044 VDDD.n1663 VSUBS 0.118956f
C8045 VDDD.n1664 VSUBS 0.118956f
C8046 VDDD.n1665 VSUBS 0.11352f
C8047 VDDD.n1666 VSUBS 0.676923f
C8048 VDDD.n1667 VSUBS 0.315547f
C8049 VDDD.n1668 VSUBS 0.251622f
C8050 VDDD.n1669 VSUBS 0.057151f
C8051 VDDD.n1670 VSUBS 0.521062f
C8052 VDDD.n1671 VSUBS 0.032934f
C8053 VDDD.n1672 VSUBS 0.226774f
C8054 VDDD.n1673 VSUBS 0.05037f
C8055 VDDD.n1674 VSUBS 0.251622f
C8056 VDDD.n1675 VSUBS 0.251622f
C8057 VDDD.n1676 VSUBS 0.251622f
C8058 VDDD.n1677 VSUBS 0.070712f
C8059 VDDD.n1678 VSUBS 0.089116f
C8060 VDDD.n1679 VSUBS 0.085726f
C8061 VDDD.n1680 VSUBS 0.251622f
C8062 VDDD.n1681 VSUBS 0.251622f
C8063 VDDD.n1682 VSUBS 0.251622f
C8064 VDDD.n1683 VSUBS 0.056666f
C8065 VDDD.n1684 VSUBS 0.049401f
C8066 VDDD.n1685 VSUBS 0.235104f
C8067 VDDD.n1686 VSUBS 0.052307f
C8068 VDDD.n1687 VSUBS 0.251622f
C8069 VDDD.n1688 VSUBS 0.251622f
C8070 VDDD.n1689 VSUBS 0.251622f
C8071 VDDD.n1690 VSUBS 0.089116f
C8072 VDDD.n1691 VSUBS 0.08621f
C8073 VDDD.n1692 VSUBS 0.250175f
C8074 VDDD.n1693 VSUBS 0.251622f
C8075 VDDD.n1694 VSUBS 0.251622f
C8076 VDDD.n1695 VSUBS 0.251622f
C8077 VDDD.n1696 VSUBS 0.074102f
C8078 VDDD.n1697 VSUBS 0.305072f
C8079 VDDD.n1698 VSUBS 0.062962f
C8080 VDDD.n1699 VSUBS 0.149059f
C8081 VDDD.n1700 VSUBS 0.188716f
C8082 VDDD.n1701 VSUBS 0.251622f
C8083 VDDD.n1702 VSUBS 0.057151f
C8084 VDDD.n1703 VSUBS 0.521062f
C8085 VDDD.n1704 VSUBS 0.032934f
C8086 VDDD.n1705 VSUBS 0.226774f
C8087 VDDD.n1706 VSUBS 0.05037f
C8088 VDDD.n1707 VSUBS 0.251622f
C8089 VDDD.n1708 VSUBS 0.251622f
C8090 VDDD.n1709 VSUBS 0.251622f
C8091 VDDD.n1710 VSUBS 0.070712f
C8092 VDDD.n1711 VSUBS 0.089116f
C8093 VDDD.n1712 VSUBS 0.085726f
C8094 VDDD.n1713 VSUBS 0.251622f
C8095 VDDD.n1714 VSUBS 0.251622f
C8096 VDDD.n1715 VSUBS 0.251622f
C8097 VDDD.n1716 VSUBS 0.056666f
C8098 VDDD.n1717 VSUBS 0.049401f
C8099 VDDD.n1718 VSUBS 0.235104f
C8100 VDDD.n1719 VSUBS 0.052307f
C8101 VDDD.n1720 VSUBS 0.251622f
C8102 VDDD.n1721 VSUBS 0.251622f
C8103 VDDD.n1722 VSUBS 0.251622f
C8104 VDDD.n1723 VSUBS 0.089116f
C8105 VDDD.n1724 VSUBS 0.08621f
C8106 VDDD.n1725 VSUBS 0.250175f
C8107 VDDD.n1726 VSUBS 0.251622f
C8108 VDDD.n1727 VSUBS 0.251622f
C8109 VDDD.n1728 VSUBS 0.251622f
C8110 VDDD.n1729 VSUBS 0.074102f
C8111 VDDD.n1730 VSUBS 0.305072f
C8112 VDDD.n1731 VSUBS 0.062962f
C8113 VDDD.n1732 VSUBS 0.149059f
C8114 VDDD.n1733 VSUBS 0.188716f
C8115 VDDD.n1734 VSUBS 0.251622f
C8116 VDDD.n1735 VSUBS 0.057151f
C8117 VDDD.n1736 VSUBS 0.521062f
C8118 VDDD.n1737 VSUBS 0.032934f
C8119 VDDD.n1738 VSUBS 0.226774f
C8120 VDDD.n1739 VSUBS 0.05037f
C8121 VDDD.n1740 VSUBS 0.251622f
C8122 VDDD.n1741 VSUBS 0.251622f
C8123 VDDD.n1742 VSUBS 0.251622f
C8124 VDDD.n1743 VSUBS 0.070712f
C8125 VDDD.n1744 VSUBS 0.089116f
C8126 VDDD.n1745 VSUBS 0.085726f
C8127 VDDD.n1746 VSUBS 0.251622f
C8128 VDDD.n1747 VSUBS 0.251622f
C8129 VDDD.n1748 VSUBS 0.251622f
C8130 VDDD.n1749 VSUBS 0.056666f
C8131 VDDD.n1750 VSUBS 0.049401f
C8132 VDDD.n1751 VSUBS 0.235104f
C8133 VDDD.n1752 VSUBS 0.052307f
C8134 VDDD.n1753 VSUBS 0.251622f
C8135 VDDD.n1754 VSUBS 0.251622f
C8136 VDDD.n1755 VSUBS 0.251622f
C8137 VDDD.n1756 VSUBS 0.089116f
C8138 VDDD.n1757 VSUBS 0.08621f
C8139 VDDD.n1758 VSUBS 0.250175f
C8140 VDDD.n1759 VSUBS 0.251622f
C8141 VDDD.n1760 VSUBS 0.251622f
C8142 VDDD.n1761 VSUBS 0.251622f
C8143 VDDD.n1762 VSUBS 0.074102f
C8144 VDDD.n1763 VSUBS 0.305072f
C8145 VDDD.n1764 VSUBS 0.062962f
C8146 VDDD.n1765 VSUBS 0.149059f
C8147 VDDD.n1766 VSUBS 0.188716f
C8148 VDDD.n1767 VSUBS 0.251622f
C8149 VDDD.n1768 VSUBS 0.057151f
C8150 VDDD.n1769 VSUBS 0.521062f
C8151 VDDD.n1770 VSUBS 0.032934f
C8152 VDDD.n1771 VSUBS 0.226774f
C8153 VDDD.n1772 VSUBS 0.05037f
C8154 VDDD.n1773 VSUBS 0.251622f
C8155 VDDD.n1774 VSUBS 0.251622f
C8156 VDDD.n1775 VSUBS 0.251622f
C8157 VDDD.n1776 VSUBS 0.070712f
C8158 VDDD.n1777 VSUBS 0.089116f
C8159 VDDD.n1778 VSUBS 0.085726f
C8160 VDDD.n1779 VSUBS 0.251622f
C8161 VDDD.n1780 VSUBS 0.251622f
C8162 VDDD.n1781 VSUBS 0.251622f
C8163 VDDD.n1782 VSUBS 0.056666f
C8164 VDDD.n1783 VSUBS 0.049401f
C8165 VDDD.n1784 VSUBS 0.235104f
C8166 VDDD.n1785 VSUBS 0.052307f
C8167 VDDD.n1786 VSUBS 0.251622f
C8168 VDDD.n1787 VSUBS 0.251622f
C8169 VDDD.n1788 VSUBS 0.251622f
C8170 VDDD.n1789 VSUBS 0.089116f
C8171 VDDD.n1790 VSUBS 0.08621f
C8172 VDDD.n1791 VSUBS 0.250175f
C8173 VDDD.n1792 VSUBS 0.251622f
C8174 VDDD.n1793 VSUBS 0.251622f
C8175 VDDD.n1794 VSUBS 0.251622f
C8176 VDDD.n1795 VSUBS 0.074102f
C8177 VDDD.n1796 VSUBS 0.305072f
C8178 VDDD.n1797 VSUBS 0.062962f
C8179 VDDD.n1798 VSUBS 0.149059f
C8180 VDDD.n1799 VSUBS 0.188716f
C8181 VDDD.n1800 VSUBS 0.251622f
C8182 VDDD.n1801 VSUBS 0.057151f
C8183 VDDD.n1802 VSUBS 0.521062f
C8184 VDDD.n1803 VSUBS 0.032934f
C8185 VDDD.n1804 VSUBS 0.251622f
C8186 VDDD.n1805 VSUBS 0.251622f
C8187 VDDD.n1806 VSUBS 0.05037f
C8188 VDDD.n1807 VSUBS 0.24113f
C8189 VDDD.n1808 VSUBS 0.070712f
C8190 VDDD.n1809 VSUBS 0.251622f
C8191 VDDD.n1810 VSUBS 0.251622f
C8192 VDDD.n1811 VSUBS 0.251622f
C8193 VDDD.n1812 VSUBS 0.085726f
C8194 VDDD.n1813 VSUBS 0.3381f
C8195 VDDD.n1814 VSUBS 0.056666f
C8196 VDDD.t637 VSUBS 0.032307f
C8197 VDDD.t1028 VSUBS 0.047863f
C8198 VDDD.n1815 VSUBS 0.083298f
C8199 VDDD.n1816 VSUBS 0.235104f
C8200 VDDD.n1817 VSUBS 0.049401f
C8201 VDDD.n1818 VSUBS 0.251622f
C8202 VDDD.n1819 VSUBS 0.251622f
C8203 VDDD.n1820 VSUBS 0.251622f
C8204 VDDD.n1821 VSUBS 0.089116f
C8205 VDDD.n1822 VSUBS 0.089116f
C8206 VDDD.n1823 VSUBS 0.08621f
C8207 VDDD.n1824 VSUBS 0.251622f
C8208 VDDD.n1825 VSUBS 0.251622f
C8209 VDDD.n1826 VSUBS 0.251622f
C8210 VDDD.n1827 VSUBS 0.067806f
C8211 VDDD.n1828 VSUBS 0.074102f
C8212 VDDD.n1829 VSUBS 0.326891f
C8213 VDDD.n1830 VSUBS 0.242239f
C8214 VDDD.n1831 VSUBS 0.118956f
C8215 VDDD.n1832 VSUBS 0.11352f
C8216 VDDD.n1833 VSUBS 0.11352f
C8217 VDDD.n1834 VSUBS 0.61245f
C8218 VDDD.t1306 VSUBS 2.12169f
C8219 VDDD.t1430 VSUBS 1.03341f
C8220 VDDD.t471 VSUBS 0.768199f
C8221 VDDD.t173 VSUBS 0.768199f
C8222 VDDD.t1428 VSUBS 0.768199f
C8223 VDDD.t572 VSUBS 0.768199f
C8224 VDDD.t473 VSUBS 0.768199f
C8225 VDDD.t225 VSUBS 0.768199f
C8226 VDDD.t469 VSUBS 0.832215f
C8227 VDDD.t129 VSUBS 0.992243f
C8228 VDDD.t189 VSUBS 0.768199f
C8229 VDDD.t1003 VSUBS 0.768199f
C8230 VDDD.t191 VSUBS 0.727031f
C8231 VDDD.t619 VSUBS 0.955662f
C8232 VDDD.t768 VSUBS 0.69045f
C8233 VDDD.n1835 VSUBS 0.564272f
C8234 VDDD.n1836 VSUBS 0.118956f
C8235 VDDD.n1837 VSUBS 0.11352f
C8236 VDDD.n1839 VSUBS 0.427239f
C8237 VDDD.n1840 VSUBS 0.118956f
C8238 VDDD.n1841 VSUBS 0.11364f
C8239 VDDD.n1842 VSUBS 0.251622f
C8240 VDDD.t769 VSUBS 0.3066f
C8241 VDDD.n1843 VSUBS 0.188716f
C8242 VDDD.t620 VSUBS 0.306452f
C8243 VDDD.n1844 VSUBS 0.149059f
C8244 VDDD.t192 VSUBS 0.306813f
C8245 VDDD.t190 VSUBS 0.076922f
C8246 VDDD.t1004 VSUBS 0.076922f
C8247 VDDD.n1845 VSUBS 0.165125f
C8248 VDDD.n1846 VSUBS 0.23282f
C8249 VDDD.n1847 VSUBS 0.188716f
C8250 VDDD.t130 VSUBS 0.269235f
C8251 VDDD.t470 VSUBS 0.292897f
C8252 VDDD.n1848 VSUBS 0.305132f
C8253 VDDD.n1849 VSUBS 0.251622f
C8254 VDDD.t474 VSUBS 0.076922f
C8255 VDDD.t226 VSUBS 0.076922f
C8256 VDDD.n1850 VSUBS 0.165125f
C8257 VDDD.n1851 VSUBS 0.047948f
C8258 VDDD.n1852 VSUBS 0.251622f
C8259 VDDD.t472 VSUBS 0.076922f
C8260 VDDD.t174 VSUBS 0.076922f
C8261 VDDD.n1853 VSUBS 0.165125f
C8262 VDDD.t1431 VSUBS 0.292867f
C8263 VDDD.n1854 VSUBS 0.398428f
C8264 VDDD.t1307 VSUBS 0.31498f
C8265 VDDD.n1855 VSUBS 0.658939f
C8266 VDDD.n1856 VSUBS 0.188716f
C8267 VDDD.n1857 VSUBS 0.251622f
C8268 VDDD.n1858 VSUBS 0.068774f
C8269 VDDD.n1859 VSUBS 0.048917f
C8270 VDDD.n1860 VSUBS 0.188262f
C8271 VDDD.t1429 VSUBS 0.076922f
C8272 VDDD.t573 VSUBS 0.076922f
C8273 VDDD.n1861 VSUBS 0.165125f
C8274 VDDD.n1862 VSUBS 0.188262f
C8275 VDDD.n1863 VSUBS 0.081367f
C8276 VDDD.n1864 VSUBS 0.251622f
C8277 VDDD.n1865 VSUBS 0.251622f
C8278 VDDD.n1866 VSUBS 0.251622f
C8279 VDDD.n1867 VSUBS 0.077977f
C8280 VDDD.n1868 VSUBS 0.188262f
C8281 VDDD.n1869 VSUBS 0.055697f
C8282 VDDD.n1870 VSUBS 0.061994f
C8283 VDDD.n1871 VSUBS 0.251622f
C8284 VDDD.n1872 VSUBS 0.149059f
C8285 VDDD.n1873 VSUBS 0.042621f
C8286 VDDD.n1874 VSUBS 0.246601f
C8287 VDDD.n1875 VSUBS 0.073133f
C8288 VDDD.n1876 VSUBS 0.251622f
C8289 VDDD.n1877 VSUBS 0.251622f
C8290 VDDD.n1878 VSUBS 0.251622f
C8291 VDDD.n1879 VSUBS 0.073133f
C8292 VDDD.n1880 VSUBS 0.440304f
C8293 VDDD.n1881 VSUBS 0.362431f
C8294 VDDD.n1882 VSUBS 0.0649f
C8295 VDDD.n1883 VSUBS 0.341286f
C8296 VDDD.n1884 VSUBS 0.149059f
C8297 VDDD.n1885 VSUBS 4.79262f
C8298 VDDD.n1886 VSUBS 0.299607f
C8299 VDDD.t1286 VSUBS 0.04923f
C8300 VDDD.t1050 VSUBS 0.04923f
C8301 VDDD.n1887 VSUBS 0.102503f
C8302 VDDD.t506 VSUBS 0.118653f
C8303 VDDD.n1888 VSUBS 0.250175f
C8304 VDDD.n1889 VSUBS 0.251622f
C8305 VDDD.n1890 VSUBS 0.052307f
C8306 VDDD.n1891 VSUBS 0.251622f
C8307 VDDD.n1892 VSUBS 0.251622f
C8308 VDDD.t549 VSUBS 0.229702f
C8309 VDDD.n1893 VSUBS 0.089116f
C8310 VDDD.n1894 VSUBS 0.251622f
C8311 VDDD.t304 VSUBS 0.032307f
C8312 VDDD.t1399 VSUBS 0.061025f
C8313 VDDD.n1895 VSUBS 0.096588f
C8314 VDDD.t433 VSUBS 0.121884f
C8315 VDDD.n1896 VSUBS 0.226774f
C8316 VDDD.n1897 VSUBS 0.251622f
C8317 VDDD.t196 VSUBS 0.337079f
C8318 VDDD.t198 VSUBS 0.306728f
C8319 VDDD.n1898 VSUBS 0.427682f
C8320 VDDD.n1899 VSUBS 0.251622f
C8321 VDDD.t395 VSUBS 0.04923f
C8322 VDDD.t568 VSUBS 0.04923f
C8323 VDDD.n1900 VSUBS 0.102503f
C8324 VDDD.n1901 VSUBS 0.067806f
C8325 VDDD.n1902 VSUBS 0.251622f
C8326 VDDD.t622 VSUBS 0.118653f
C8327 VDDD.n1903 VSUBS 0.089116f
C8328 VDDD.n1904 VSUBS 0.251622f
C8329 VDDD.t1415 VSUBS 0.032307f
C8330 VDDD.t559 VSUBS 0.047863f
C8331 VDDD.n1905 VSUBS 0.083298f
C8332 VDDD.t443 VSUBS 0.229702f
C8333 VDDD.n1906 VSUBS 0.3381f
C8334 VDDD.n1907 VSUBS 0.251622f
C8335 VDDD.t1200 VSUBS 0.032307f
C8336 VDDD.t45 VSUBS 0.061025f
C8337 VDDD.n1908 VSUBS 0.096588f
C8338 VDDD.n1909 VSUBS 0.24113f
C8339 VDDD.n1910 VSUBS 0.251622f
C8340 VDDD.t1258 VSUBS 0.121884f
C8341 VDDD.n1911 VSUBS 0.251622f
C8342 VDDD.t51 VSUBS 0.337079f
C8343 VDDD.t49 VSUBS 0.306728f
C8344 VDDD.n1912 VSUBS 0.427682f
C8345 VDDD.n1913 VSUBS 0.251622f
C8346 VDDD.t844 VSUBS 0.04923f
C8347 VDDD.t339 VSUBS 0.04923f
C8348 VDDD.n1914 VSUBS 0.102503f
C8349 VDDD.n1915 VSUBS 0.067806f
C8350 VDDD.n1916 VSUBS 0.251622f
C8351 VDDD.t1256 VSUBS 0.118653f
C8352 VDDD.n1917 VSUBS 0.089116f
C8353 VDDD.n1918 VSUBS 0.251622f
C8354 VDDD.t11 VSUBS 0.032307f
C8355 VDDD.t419 VSUBS 0.047863f
C8356 VDDD.n1919 VSUBS 0.083298f
C8357 VDDD.t1167 VSUBS 0.229702f
C8358 VDDD.n1920 VSUBS 0.3381f
C8359 VDDD.n1921 VSUBS 0.251622f
C8360 VDDD.t206 VSUBS 0.032307f
C8361 VDDD.t277 VSUBS 0.061025f
C8362 VDDD.n1922 VSUBS 0.096588f
C8363 VDDD.n1923 VSUBS 0.24113f
C8364 VDDD.n1924 VSUBS 0.251622f
C8365 VDDD.t649 VSUBS 0.121884f
C8366 VDDD.n1925 VSUBS 0.251622f
C8367 VDDD.t1030 VSUBS 0.337079f
C8368 VDDD.t279 VSUBS 0.306728f
C8369 VDDD.n1926 VSUBS 0.427682f
C8370 VDDD.n1927 VSUBS 0.251622f
C8371 VDDD.t511 VSUBS 0.04923f
C8372 VDDD.t1018 VSUBS 0.04923f
C8373 VDDD.n1928 VSUBS 0.102503f
C8374 VDDD.n1929 VSUBS 0.067806f
C8375 VDDD.n1930 VSUBS 0.251622f
C8376 VDDD.t866 VSUBS 0.118653f
C8377 VDDD.n1931 VSUBS 0.089116f
C8378 VDDD.n1932 VSUBS 0.251622f
C8379 VDDD.t1413 VSUBS 0.032307f
C8380 VDDD.t920 VSUBS 0.047863f
C8381 VDDD.n1933 VSUBS 0.083298f
C8382 VDDD.t860 VSUBS 0.229702f
C8383 VDDD.n1934 VSUBS 0.3381f
C8384 VDDD.n1935 VSUBS 0.251622f
C8385 VDDD.t896 VSUBS 0.032307f
C8386 VDDD.t157 VSUBS 0.061025f
C8387 VDDD.n1936 VSUBS 0.096588f
C8388 VDDD.n1937 VSUBS 0.24113f
C8389 VDDD.n1938 VSUBS 0.251622f
C8390 VDDD.t327 VSUBS 0.121884f
C8391 VDDD.n1939 VSUBS 0.251622f
C8392 VDDD.t461 VSUBS 0.337079f
C8393 VDDD.t159 VSUBS 0.306728f
C8394 VDDD.n1940 VSUBS 0.427682f
C8395 VDDD.n1941 VSUBS 0.251622f
C8396 VDDD.t359 VSUBS 0.04923f
C8397 VDDD.t1113 VSUBS 0.04923f
C8398 VDDD.n1942 VSUBS 0.102503f
C8399 VDDD.n1943 VSUBS 0.067806f
C8400 VDDD.n1944 VSUBS 0.251622f
C8401 VDDD.t1343 VSUBS 0.118653f
C8402 VDDD.n1945 VSUBS 0.089116f
C8403 VDDD.n1946 VSUBS 0.251622f
C8404 VDDD.t13 VSUBS 0.032307f
C8405 VDDD.t561 VSUBS 0.047863f
C8406 VDDD.n1947 VSUBS 0.083298f
C8407 VDDD.t16 VSUBS 0.229702f
C8408 VDDD.n1948 VSUBS 0.3381f
C8409 VDDD.n1949 VSUBS 0.251622f
C8410 VDDD.t1198 VSUBS 0.032307f
C8411 VDDD.t55 VSUBS 0.061025f
C8412 VDDD.n1950 VSUBS 0.096588f
C8413 VDDD.n1951 VSUBS 0.24113f
C8414 VDDD.n1952 VSUBS 0.251622f
C8415 VDDD.t787 VSUBS 0.121884f
C8416 VDDD.n1953 VSUBS 0.251622f
C8417 VDDD.t53 VSUBS 0.337079f
C8418 VDDD.t728 VSUBS 0.306728f
C8419 VDDD.n1954 VSUBS 0.427682f
C8420 VDDD.n1955 VSUBS 0.251622f
C8421 VDDD.t250 VSUBS 0.04923f
C8422 VDDD.t566 VSUBS 0.04923f
C8423 VDDD.n1956 VSUBS 0.102503f
C8424 VDDD.n1957 VSUBS 0.067806f
C8425 VDDD.n1958 VSUBS 0.251622f
C8426 VDDD.t128 VSUBS 0.118653f
C8427 VDDD.n1959 VSUBS 0.089116f
C8428 VDDD.n1960 VSUBS 0.251622f
C8429 VDDD.t1323 VSUBS 0.032307f
C8430 VDDD.t1281 VSUBS 0.047863f
C8431 VDDD.n1961 VSUBS 0.083298f
C8432 VDDD.t1170 VSUBS 0.229702f
C8433 VDDD.n1962 VSUBS 0.3381f
C8434 VDDD.n1963 VSUBS 0.251622f
C8435 VDDD.t1417 VSUBS 0.032307f
C8436 VDDD.t406 VSUBS 0.061025f
C8437 VDDD.n1964 VSUBS 0.096588f
C8438 VDDD.n1965 VSUBS 0.24113f
C8439 VDDD.n1966 VSUBS 0.251622f
C8440 VDDD.t685 VSUBS 0.121884f
C8441 VDDD.n1967 VSUBS 0.251622f
C8442 VDDD.t404 VSUBS 0.337079f
C8443 VDDD.t408 VSUBS 0.306728f
C8444 VDDD.n1968 VSUBS 0.366172f
C8445 VDDD.n1969 VSUBS 0.118956f
C8446 VDDD.n1970 VSUBS 0.11352f
C8447 VDDD.n1971 VSUBS 0.11352f
C8448 VDDD.n1972 VSUBS 0.11352f
C8449 VDDD.t1049 VSUBS 0.681305f
C8450 VDDD.t1285 VSUBS 1.60497f
C8451 VDDD.t505 VSUBS 1.64155f
C8452 VDDD.t431 VSUBS 0.873355f
C8453 VDDD.t1171 VSUBS 1.09284f
C8454 VDDD.t673 VSUBS 1.08369f
C8455 VDDD.t868 VSUBS 1.34432f
C8456 VDDD.t548 VSUBS 1.35346f
C8457 VDDD.t1172 VSUBS 0.845919f
C8458 VDDD.t430 VSUBS 0.777344f
C8459 VDDD.t1398 VSUBS 0.877942f
C8460 VDDD.t303 VSUBS 0.877942f
C8461 VDDD.t432 VSUBS 1.3672f
C8462 VDDD.t195 VSUBS 1.3672f
C8463 VDDD.t197 VSUBS 0.983097f
C8464 VDDD.t567 VSUBS 0.681305f
C8465 VDDD.t394 VSUBS 1.60497f
C8466 VDDD.t621 VSUBS 1.64155f
C8467 VDDD.t747 VSUBS 0.873355f
C8468 VDDD.t772 VSUBS 1.09284f
C8469 VDDD.t558 VSUBS 1.08369f
C8470 VDDD.t1414 VSUBS 1.34432f
C8471 VDDD.t442 VSUBS 1.35346f
C8472 VDDD.t396 VSUBS 0.845919f
C8473 VDDD.t876 VSUBS 0.777344f
C8474 VDDD.t44 VSUBS 0.877942f
C8475 VDDD.t1199 VSUBS 0.877942f
C8476 VDDD.t1257 VSUBS 1.3672f
C8477 VDDD.t50 VSUBS 1.3672f
C8478 VDDD.t48 VSUBS 0.983097f
C8479 VDDD.t338 VSUBS 0.681305f
C8480 VDDD.t843 VSUBS 1.60497f
C8481 VDDD.t1255 VSUBS 1.64155f
C8482 VDDD.t437 VSUBS 0.873355f
C8483 VDDD.t447 VSUBS 1.09284f
C8484 VDDD.t418 VSUBS 1.08369f
C8485 VDDD.t10 VSUBS 1.34432f
C8486 VDDD.t1166 VSUBS 1.35346f
C8487 VDDD.t1375 VSUBS 0.845919f
C8488 VDDD.t409 VSUBS 0.777344f
C8489 VDDD.t276 VSUBS 0.877942f
C8490 VDDD.t205 VSUBS 0.877942f
C8491 VDDD.t648 VSUBS 1.3672f
C8492 VDDD.t1029 VSUBS 1.3672f
C8493 VDDD.t278 VSUBS 0.983097f
C8494 VDDD.t1017 VSUBS 0.681305f
C8495 VDDD.t510 VSUBS 1.60497f
C8496 VDDD.t865 VSUBS 1.64155f
C8497 VDDD.t675 VSUBS 0.873355f
C8498 VDDD.t512 VSUBS 1.09284f
C8499 VDDD.t919 VSUBS 1.08369f
C8500 VDDD.t1412 VSUBS 1.34432f
C8501 VDDD.t859 VSUBS 1.35346f
C8502 VDDD.t477 VSUBS 0.845919f
C8503 VDDD.t972 VSUBS 0.777344f
C8504 VDDD.t156 VSUBS 0.877942f
C8505 VDDD.t895 VSUBS 0.877942f
C8506 VDDD.t326 VSUBS 1.3672f
C8507 VDDD.t460 VSUBS 1.3672f
C8508 VDDD.t158 VSUBS 0.983097f
C8509 VDDD.t1112 VSUBS 0.681305f
C8510 VDDD.t358 VSUBS 1.60497f
C8511 VDDD.t1342 VSUBS 1.64155f
C8512 VDDD.t56 VSUBS 0.873355f
C8513 VDDD.t357 VSUBS 1.09284f
C8514 VDDD.t560 VSUBS 1.08369f
C8515 VDDD.t12 VSUBS 1.34432f
C8516 VDDD.t15 VSUBS 1.35346f
C8517 VDDD.t14 VSUBS 0.845919f
C8518 VDDD.t9 VSUBS 0.777344f
C8519 VDDD.t54 VSUBS 0.877942f
C8520 VDDD.t1197 VSUBS 0.877942f
C8521 VDDD.t786 VSUBS 1.3672f
C8522 VDDD.t52 VSUBS 1.3672f
C8523 VDDD.t727 VSUBS 0.983097f
C8524 VDDD.t565 VSUBS 0.681305f
C8525 VDDD.t249 VSUBS 1.60497f
C8526 VDDD.t127 VSUBS 1.64155f
C8527 VDDD.t383 VSUBS 0.873355f
C8528 VDDD.t248 VSUBS 1.09284f
C8529 VDDD.t1280 VSUBS 1.08369f
C8530 VDDD.t1322 VSUBS 1.34432f
C8531 VDDD.t1169 VSUBS 1.35346f
C8532 VDDD.t251 VSUBS 0.845919f
C8533 VDDD.t110 VSUBS 0.777344f
C8534 VDDD.t405 VSUBS 0.877942f
C8535 VDDD.t1416 VSUBS 0.877942f
C8536 VDDD.t684 VSUBS 1.3672f
C8537 VDDD.t403 VSUBS 1.3672f
C8538 VDDD.t407 VSUBS 1.02427f
C8539 VDDD.n1973 VSUBS 0.427239f
C8540 VDDD.n1975 VSUBS 0.61245f
C8541 VDDD.n1976 VSUBS 0.833326f
C8542 VDDD.n1977 VSUBS 0.118956f
C8543 VDDD.n1978 VSUBS 0.118956f
C8544 VDDD.n1979 VSUBS 0.128942f
C8545 VDDD.n1980 VSUBS 1.07369f
C8546 VDDD.n1981 VSUBS 0.251622f
C8547 VDDD.n1982 VSUBS 0.057151f
C8548 VDDD.n1983 VSUBS 0.521062f
C8549 VDDD.n1984 VSUBS 0.032934f
C8550 VDDD.n1985 VSUBS 0.226774f
C8551 VDDD.n1986 VSUBS 0.05037f
C8552 VDDD.n1987 VSUBS 0.251622f
C8553 VDDD.n1988 VSUBS 0.251622f
C8554 VDDD.n1989 VSUBS 0.251622f
C8555 VDDD.n1990 VSUBS 0.070712f
C8556 VDDD.n1991 VSUBS 0.089116f
C8557 VDDD.n1992 VSUBS 0.085726f
C8558 VDDD.n1993 VSUBS 0.251622f
C8559 VDDD.n1994 VSUBS 0.251622f
C8560 VDDD.n1995 VSUBS 0.251622f
C8561 VDDD.n1996 VSUBS 0.056666f
C8562 VDDD.n1997 VSUBS 0.049401f
C8563 VDDD.n1998 VSUBS 0.235104f
C8564 VDDD.n1999 VSUBS 0.052307f
C8565 VDDD.n2000 VSUBS 0.251622f
C8566 VDDD.n2001 VSUBS 0.251622f
C8567 VDDD.n2002 VSUBS 0.251622f
C8568 VDDD.n2003 VSUBS 0.089116f
C8569 VDDD.n2004 VSUBS 0.08621f
C8570 VDDD.n2005 VSUBS 0.250175f
C8571 VDDD.n2006 VSUBS 0.251622f
C8572 VDDD.n2007 VSUBS 0.251622f
C8573 VDDD.n2008 VSUBS 0.251622f
C8574 VDDD.n2009 VSUBS 0.074102f
C8575 VDDD.n2010 VSUBS 0.305072f
C8576 VDDD.n2011 VSUBS 0.062962f
C8577 VDDD.n2012 VSUBS 0.149059f
C8578 VDDD.n2013 VSUBS 0.188716f
C8579 VDDD.n2014 VSUBS 0.251622f
C8580 VDDD.n2015 VSUBS 0.057151f
C8581 VDDD.n2016 VSUBS 0.521062f
C8582 VDDD.n2017 VSUBS 0.032934f
C8583 VDDD.n2018 VSUBS 0.226774f
C8584 VDDD.n2019 VSUBS 0.05037f
C8585 VDDD.n2020 VSUBS 0.251622f
C8586 VDDD.n2021 VSUBS 0.251622f
C8587 VDDD.n2022 VSUBS 0.251622f
C8588 VDDD.n2023 VSUBS 0.070712f
C8589 VDDD.n2024 VSUBS 0.089116f
C8590 VDDD.n2025 VSUBS 0.085726f
C8591 VDDD.n2026 VSUBS 0.251622f
C8592 VDDD.n2027 VSUBS 0.251622f
C8593 VDDD.n2028 VSUBS 0.251622f
C8594 VDDD.n2029 VSUBS 0.056666f
C8595 VDDD.n2030 VSUBS 0.049401f
C8596 VDDD.n2031 VSUBS 0.235104f
C8597 VDDD.n2032 VSUBS 0.052307f
C8598 VDDD.n2033 VSUBS 0.251622f
C8599 VDDD.n2034 VSUBS 0.251622f
C8600 VDDD.n2035 VSUBS 0.251622f
C8601 VDDD.n2036 VSUBS 0.089116f
C8602 VDDD.n2037 VSUBS 0.08621f
C8603 VDDD.n2038 VSUBS 0.250175f
C8604 VDDD.n2039 VSUBS 0.251622f
C8605 VDDD.n2040 VSUBS 0.251622f
C8606 VDDD.n2041 VSUBS 0.251622f
C8607 VDDD.n2042 VSUBS 0.074102f
C8608 VDDD.n2043 VSUBS 0.305072f
C8609 VDDD.n2044 VSUBS 0.062962f
C8610 VDDD.n2045 VSUBS 0.149059f
C8611 VDDD.n2046 VSUBS 0.188716f
C8612 VDDD.n2047 VSUBS 0.251622f
C8613 VDDD.n2048 VSUBS 0.057151f
C8614 VDDD.n2049 VSUBS 0.521062f
C8615 VDDD.n2050 VSUBS 0.032934f
C8616 VDDD.n2051 VSUBS 0.226774f
C8617 VDDD.n2052 VSUBS 0.05037f
C8618 VDDD.n2053 VSUBS 0.251622f
C8619 VDDD.n2054 VSUBS 0.251622f
C8620 VDDD.n2055 VSUBS 0.251622f
C8621 VDDD.n2056 VSUBS 0.070712f
C8622 VDDD.n2057 VSUBS 0.089116f
C8623 VDDD.n2058 VSUBS 0.085726f
C8624 VDDD.n2059 VSUBS 0.251622f
C8625 VDDD.n2060 VSUBS 0.251622f
C8626 VDDD.n2061 VSUBS 0.251622f
C8627 VDDD.n2062 VSUBS 0.056666f
C8628 VDDD.n2063 VSUBS 0.049401f
C8629 VDDD.n2064 VSUBS 0.235104f
C8630 VDDD.n2065 VSUBS 0.052307f
C8631 VDDD.n2066 VSUBS 0.251622f
C8632 VDDD.n2067 VSUBS 0.251622f
C8633 VDDD.n2068 VSUBS 0.251622f
C8634 VDDD.n2069 VSUBS 0.089116f
C8635 VDDD.n2070 VSUBS 0.08621f
C8636 VDDD.n2071 VSUBS 0.250175f
C8637 VDDD.n2072 VSUBS 0.251622f
C8638 VDDD.n2073 VSUBS 0.251622f
C8639 VDDD.n2074 VSUBS 0.251622f
C8640 VDDD.n2075 VSUBS 0.074102f
C8641 VDDD.n2076 VSUBS 0.305072f
C8642 VDDD.n2077 VSUBS 0.062962f
C8643 VDDD.n2078 VSUBS 0.149059f
C8644 VDDD.n2079 VSUBS 0.188716f
C8645 VDDD.n2080 VSUBS 0.251622f
C8646 VDDD.n2081 VSUBS 0.057151f
C8647 VDDD.n2082 VSUBS 0.521062f
C8648 VDDD.n2083 VSUBS 0.032934f
C8649 VDDD.n2084 VSUBS 0.226774f
C8650 VDDD.n2085 VSUBS 0.05037f
C8651 VDDD.n2086 VSUBS 0.251622f
C8652 VDDD.n2087 VSUBS 0.251622f
C8653 VDDD.n2088 VSUBS 0.251622f
C8654 VDDD.n2089 VSUBS 0.070712f
C8655 VDDD.n2090 VSUBS 0.089116f
C8656 VDDD.n2091 VSUBS 0.085726f
C8657 VDDD.n2092 VSUBS 0.251622f
C8658 VDDD.n2093 VSUBS 0.251622f
C8659 VDDD.n2094 VSUBS 0.251622f
C8660 VDDD.n2095 VSUBS 0.056666f
C8661 VDDD.n2096 VSUBS 0.049401f
C8662 VDDD.n2097 VSUBS 0.235104f
C8663 VDDD.n2098 VSUBS 0.052307f
C8664 VDDD.n2099 VSUBS 0.251622f
C8665 VDDD.n2100 VSUBS 0.251622f
C8666 VDDD.n2101 VSUBS 0.251622f
C8667 VDDD.n2102 VSUBS 0.089116f
C8668 VDDD.n2103 VSUBS 0.08621f
C8669 VDDD.n2104 VSUBS 0.250175f
C8670 VDDD.n2105 VSUBS 0.251622f
C8671 VDDD.n2106 VSUBS 0.251622f
C8672 VDDD.n2107 VSUBS 0.251622f
C8673 VDDD.n2108 VSUBS 0.074102f
C8674 VDDD.n2109 VSUBS 0.305072f
C8675 VDDD.n2110 VSUBS 0.062962f
C8676 VDDD.n2111 VSUBS 0.149059f
C8677 VDDD.n2112 VSUBS 0.188716f
C8678 VDDD.n2113 VSUBS 0.251622f
C8679 VDDD.n2114 VSUBS 0.057151f
C8680 VDDD.n2115 VSUBS 0.521062f
C8681 VDDD.n2116 VSUBS 0.032934f
C8682 VDDD.n2117 VSUBS 0.226774f
C8683 VDDD.n2118 VSUBS 0.05037f
C8684 VDDD.n2119 VSUBS 0.251622f
C8685 VDDD.n2120 VSUBS 0.251622f
C8686 VDDD.n2121 VSUBS 0.251622f
C8687 VDDD.n2122 VSUBS 0.070712f
C8688 VDDD.n2123 VSUBS 0.089116f
C8689 VDDD.n2124 VSUBS 0.085726f
C8690 VDDD.n2125 VSUBS 0.251622f
C8691 VDDD.n2126 VSUBS 0.251622f
C8692 VDDD.n2127 VSUBS 0.251622f
C8693 VDDD.n2128 VSUBS 0.056666f
C8694 VDDD.n2129 VSUBS 0.049401f
C8695 VDDD.n2130 VSUBS 0.235104f
C8696 VDDD.n2131 VSUBS 0.052307f
C8697 VDDD.n2132 VSUBS 0.251622f
C8698 VDDD.n2133 VSUBS 0.251622f
C8699 VDDD.n2134 VSUBS 0.251622f
C8700 VDDD.n2135 VSUBS 0.089116f
C8701 VDDD.n2136 VSUBS 0.08621f
C8702 VDDD.n2137 VSUBS 0.250175f
C8703 VDDD.n2138 VSUBS 0.251622f
C8704 VDDD.n2139 VSUBS 0.251622f
C8705 VDDD.n2140 VSUBS 0.251622f
C8706 VDDD.n2141 VSUBS 0.074102f
C8707 VDDD.n2142 VSUBS 0.305072f
C8708 VDDD.n2143 VSUBS 0.062962f
C8709 VDDD.n2144 VSUBS 0.149059f
C8710 VDDD.n2145 VSUBS 0.188716f
C8711 VDDD.n2146 VSUBS 0.251622f
C8712 VDDD.n2147 VSUBS 0.057151f
C8713 VDDD.n2148 VSUBS 0.521062f
C8714 VDDD.n2149 VSUBS 0.032934f
C8715 VDDD.n2150 VSUBS 0.251622f
C8716 VDDD.n2151 VSUBS 0.251622f
C8717 VDDD.n2152 VSUBS 0.05037f
C8718 VDDD.n2153 VSUBS 0.24113f
C8719 VDDD.n2154 VSUBS 0.070712f
C8720 VDDD.n2155 VSUBS 0.251622f
C8721 VDDD.n2156 VSUBS 0.251622f
C8722 VDDD.n2157 VSUBS 0.251622f
C8723 VDDD.n2158 VSUBS 0.085726f
C8724 VDDD.n2159 VSUBS 0.3381f
C8725 VDDD.n2160 VSUBS 0.056666f
C8726 VDDD.t869 VSUBS 0.032307f
C8727 VDDD.t674 VSUBS 0.047863f
C8728 VDDD.n2161 VSUBS 0.083298f
C8729 VDDD.n2162 VSUBS 0.235104f
C8730 VDDD.n2163 VSUBS 0.049401f
C8731 VDDD.n2164 VSUBS 0.251622f
C8732 VDDD.n2165 VSUBS 0.251622f
C8733 VDDD.n2166 VSUBS 0.251622f
C8734 VDDD.n2167 VSUBS 0.089116f
C8735 VDDD.n2168 VSUBS 0.089116f
C8736 VDDD.n2169 VSUBS 0.08621f
C8737 VDDD.n2170 VSUBS 0.251622f
C8738 VDDD.n2171 VSUBS 0.251622f
C8739 VDDD.n2172 VSUBS 0.251622f
C8740 VDDD.n2173 VSUBS 0.067806f
C8741 VDDD.n2174 VSUBS 0.074102f
C8742 VDDD.n2175 VSUBS 0.326891f
C8743 VDDD.n2176 VSUBS 0.242239f
C8744 VDDD.n2177 VSUBS 6.18301f
C8745 VDDD.n2178 VSUBS 0.299607f
C8746 VDDD.t1162 VSUBS 0.04923f
C8747 VDDD.t1026 VSUBS 0.04923f
C8748 VDDD.n2179 VSUBS 0.102503f
C8749 VDDD.t1433 VSUBS 0.118653f
C8750 VDDD.n2180 VSUBS 0.250175f
C8751 VDDD.n2181 VSUBS 0.251622f
C8752 VDDD.n2182 VSUBS 0.052307f
C8753 VDDD.n2183 VSUBS 0.251622f
C8754 VDDD.n2184 VSUBS 0.251622f
C8755 VDDD.t689 VSUBS 0.229702f
C8756 VDDD.n2185 VSUBS 0.089116f
C8757 VDDD.n2186 VSUBS 0.251622f
C8758 VDDD.t295 VSUBS 0.032307f
C8759 VDDD.t1130 VSUBS 0.061025f
C8760 VDDD.n2187 VSUBS 0.096588f
C8761 VDDD.t1383 VSUBS 0.121884f
C8762 VDDD.n2188 VSUBS 0.226774f
C8763 VDDD.n2189 VSUBS 0.251622f
C8764 VDDD.t1354 VSUBS 0.337079f
C8765 VDDD.t1352 VSUBS 0.306728f
C8766 VDDD.n2190 VSUBS 0.427682f
C8767 VDDD.n2191 VSUBS 0.251622f
C8768 VDDD.t974 VSUBS 0.04923f
C8769 VDDD.t343 VSUBS 0.04923f
C8770 VDDD.n2192 VSUBS 0.102503f
C8771 VDDD.n2193 VSUBS 0.067806f
C8772 VDDD.n2194 VSUBS 0.251622f
C8773 VDDD.t730 VSUBS 0.118653f
C8774 VDDD.n2195 VSUBS 0.089116f
C8775 VDDD.n2196 VSUBS 0.251622f
C8776 VDDD.t1065 VSUBS 0.032307f
C8777 VDDD.t710 VSUBS 0.047863f
C8778 VDDD.n2197 VSUBS 0.083298f
C8779 VDDD.t331 VSUBS 0.229702f
C8780 VDDD.n2198 VSUBS 0.3381f
C8781 VDDD.n2199 VSUBS 0.251622f
C8782 VDDD.t1319 VSUBS 0.032307f
C8783 VDDD.t557 VSUBS 0.061025f
C8784 VDDD.n2200 VSUBS 0.096588f
C8785 VDDD.n2201 VSUBS 0.24113f
C8786 VDDD.n2202 VSUBS 0.251622f
C8787 VDDD.t609 VSUBS 0.121884f
C8788 VDDD.n2203 VSUBS 0.251622f
C8789 VDDD.t555 VSUBS 0.337079f
C8790 VDDD.t553 VSUBS 0.306728f
C8791 VDDD.n2204 VSUBS 0.427682f
C8792 VDDD.n2205 VSUBS 0.251622f
C8793 VDDD.t659 VSUBS 0.04923f
C8794 VDDD.t345 VSUBS 0.04923f
C8795 VDDD.n2206 VSUBS 0.102503f
C8796 VDDD.n2207 VSUBS 0.067806f
C8797 VDDD.n2208 VSUBS 0.251622f
C8798 VDDD.t996 VSUBS 0.118653f
C8799 VDDD.n2209 VSUBS 0.089116f
C8800 VDDD.n2210 VSUBS 0.251622f
C8801 VDDD.t781 VSUBS 0.032307f
C8802 VDDD.t114 VSUBS 0.047863f
C8803 VDDD.n2211 VSUBS 0.083298f
C8804 VDDD.t351 VSUBS 0.229702f
C8805 VDDD.n2212 VSUBS 0.3381f
C8806 VDDD.n2213 VSUBS 0.251622f
C8807 VDDD.t783 VSUBS 0.032307f
C8808 VDDD.t988 VSUBS 0.061025f
C8809 VDDD.n2214 VSUBS 0.096588f
C8810 VDDD.n2215 VSUBS 0.24113f
C8811 VDDD.n2216 VSUBS 0.251622f
C8812 VDDD.t451 VSUBS 0.121884f
C8813 VDDD.n2217 VSUBS 0.251622f
C8814 VDDD.t1210 VSUBS 0.337079f
C8815 VDDD.t990 VSUBS 0.306728f
C8816 VDDD.n2218 VSUBS 0.427682f
C8817 VDDD.n2219 VSUBS 0.251622f
C8818 VDDD.t857 VSUBS 0.04923f
C8819 VDDD.t1020 VSUBS 0.04923f
C8820 VDDD.n2220 VSUBS 0.102503f
C8821 VDDD.n2221 VSUBS 0.067806f
C8822 VDDD.n2222 VSUBS 0.251622f
C8823 VDDD.t734 VSUBS 0.118653f
C8824 VDDD.n2223 VSUBS 0.089116f
C8825 VDDD.n2224 VSUBS 0.251622f
C8826 VDDD.t1347 VSUBS 0.032307f
C8827 VDDD.t871 VSUBS 0.047863f
C8828 VDDD.n2225 VSUBS 0.083298f
C8829 VDDD.t704 VSUBS 0.229702f
C8830 VDDD.n2226 VSUBS 0.3381f
C8831 VDDD.n2227 VSUBS 0.251622f
C8832 VDDD.t1063 VSUBS 0.032307f
C8833 VDDD.t575 VSUBS 0.061025f
C8834 VDDD.n2228 VSUBS 0.096588f
C8835 VDDD.n2229 VSUBS 0.24113f
C8836 VDDD.n2230 VSUBS 0.251622f
C8837 VDDD.t961 VSUBS 0.121884f
C8838 VDDD.n2231 VSUBS 0.251622f
C8839 VDDD.t584 VSUBS 0.337079f
C8840 VDDD.t937 VSUBS 0.306728f
C8841 VDDD.n2232 VSUBS 0.427682f
C8842 VDDD.n2233 VSUBS 0.251622f
C8843 VDDD.t354 VSUBS 0.04923f
C8844 VDDD.t1117 VSUBS 0.04923f
C8845 VDDD.n2234 VSUBS 0.102503f
C8846 VDDD.n2235 VSUBS 0.067806f
C8847 VDDD.n2236 VSUBS 0.251622f
C8848 VDDD.t817 VSUBS 0.118653f
C8849 VDDD.n2237 VSUBS 0.089116f
C8850 VDDD.n2238 VSUBS 0.251622f
C8851 VDDD.t625 VSUBS 0.032307f
C8852 VDDD.t647 VSUBS 0.047863f
C8853 VDDD.n2239 VSUBS 0.083298f
C8854 VDDD.t683 VSUBS 0.229702f
C8855 VDDD.n2240 VSUBS 0.3381f
C8856 VDDD.n2241 VSUBS 0.251622f
C8857 VDDD.t293 VSUBS 0.032307f
C8858 VDDD.t106 VSUBS 0.061025f
C8859 VDDD.n2242 VSUBS 0.096588f
C8860 VDDD.n2243 VSUBS 0.24113f
C8861 VDDD.n2244 VSUBS 0.251622f
C8862 VDDD.t102 VSUBS 0.121884f
C8863 VDDD.n2245 VSUBS 0.251622f
C8864 VDDD.t104 VSUBS 0.337079f
C8865 VDDD.t108 VSUBS 0.306728f
C8866 VDDD.n2246 VSUBS 0.427682f
C8867 VDDD.n2247 VSUBS 0.251622f
C8868 VDDD.t1206 VSUBS 0.04923f
C8869 VDDD.t341 VSUBS 0.04923f
C8870 VDDD.n2248 VSUBS 0.102503f
C8871 VDDD.n2249 VSUBS 0.067806f
C8872 VDDD.n2250 VSUBS 0.251622f
C8873 VDDD.t376 VSUBS 0.118653f
C8874 VDDD.n2251 VSUBS 0.089116f
C8875 VDDD.n2252 VSUBS 0.251622f
C8876 VDDD.t777 VSUBS 0.032307f
C8877 VDDD.t136 VSUBS 0.047863f
C8878 VDDD.n2253 VSUBS 0.083298f
C8879 VDDD.t421 VSUBS 0.229702f
C8880 VDDD.n2254 VSUBS 0.3381f
C8881 VDDD.n2255 VSUBS 0.251622f
C8882 VDDD.t180 VSUBS 0.032307f
C8883 VDDD.t526 VSUBS 0.061025f
C8884 VDDD.n2256 VSUBS 0.096588f
C8885 VDDD.n2257 VSUBS 0.24113f
C8886 VDDD.n2258 VSUBS 0.251622f
C8887 VDDD.t439 VSUBS 0.121884f
C8888 VDDD.n2259 VSUBS 0.251622f
C8889 VDDD.t232 VSUBS 0.337079f
C8890 VDDD.t528 VSUBS 0.306728f
C8891 VDDD.n2260 VSUBS 0.427682f
C8892 VDDD.n2261 VSUBS 0.118956f
C8893 VDDD.n2262 VSUBS 0.11352f
C8894 VDDD.n2263 VSUBS 0.11352f
C8895 VDDD.n2264 VSUBS 0.11352f
C8896 VDDD.t1025 VSUBS 0.681305f
C8897 VDDD.t1161 VSUBS 1.60497f
C8898 VDDD.t1432 VSUBS 1.64155f
C8899 VDDD.t252 VSUBS 0.873355f
C8900 VDDD.t1133 VSUBS 1.09284f
C8901 VDDD.t508 VSUBS 1.08369f
C8902 VDDD.t181 VSUBS 1.34432f
C8903 VDDD.t688 VSUBS 1.35346f
C8904 VDDD.t589 VSUBS 0.845919f
C8905 VDDD.t582 VSUBS 0.777344f
C8906 VDDD.t1129 VSUBS 0.877942f
C8907 VDDD.t294 VSUBS 0.877942f
C8908 VDDD.t1382 VSUBS 1.3672f
C8909 VDDD.t1353 VSUBS 1.3672f
C8910 VDDD.t1351 VSUBS 0.983097f
C8911 VDDD.t342 VSUBS 0.681305f
C8912 VDDD.t973 VSUBS 1.60497f
C8913 VDDD.t729 VSUBS 1.64155f
C8914 VDDD.t17 VSUBS 0.873355f
C8915 VDDD.t818 VSUBS 1.09284f
C8916 VDDD.t709 VSUBS 1.08369f
C8917 VDDD.t1064 VSUBS 1.34432f
C8918 VDDD.t330 VSUBS 1.35346f
C8919 VDDD.t1456 VSUBS 0.845919f
C8920 VDDD.t8 VSUBS 0.777344f
C8921 VDDD.t556 VSUBS 0.877942f
C8922 VDDD.t1318 VSUBS 0.877942f
C8923 VDDD.t608 VSUBS 1.3672f
C8924 VDDD.t554 VSUBS 1.3672f
C8925 VDDD.t552 VSUBS 0.983097f
C8926 VDDD.t344 VSUBS 0.681305f
C8927 VDDD.t658 VSUBS 1.60497f
C8928 VDDD.t995 VSUBS 1.64155f
C8929 VDDD.t1223 VSUBS 0.873355f
C8930 VDDD.t657 VSUBS 1.09284f
C8931 VDDD.t113 VSUBS 1.08369f
C8932 VDDD.t780 VSUBS 1.34432f
C8933 VDDD.t350 VSUBS 1.35346f
C8934 VDDD.t124 VSUBS 0.845919f
C8935 VDDD.t1224 VSUBS 0.777344f
C8936 VDDD.t987 VSUBS 0.877942f
C8937 VDDD.t782 VSUBS 0.877942f
C8938 VDDD.t450 VSUBS 1.3672f
C8939 VDDD.t1209 VSUBS 1.3672f
C8940 VDDD.t989 VSUBS 0.983097f
C8941 VDDD.t1019 VSUBS 0.681305f
C8942 VDDD.t856 VSUBS 1.60497f
C8943 VDDD.t733 VSUBS 1.64155f
C8944 VDDD.t444 VSUBS 0.873355f
C8945 VDDD.t855 VSUBS 1.09284f
C8946 VDDD.t870 VSUBS 1.08369f
C8947 VDDD.t1346 VSUBS 1.34432f
C8948 VDDD.t703 VSUBS 1.35346f
C8949 VDDD.t1348 VSUBS 0.845919f
C8950 VDDD.t607 VSUBS 0.777344f
C8951 VDDD.t574 VSUBS 0.877942f
C8952 VDDD.t1062 VSUBS 0.877942f
C8953 VDDD.t960 VSUBS 1.3672f
C8954 VDDD.t583 VSUBS 1.3672f
C8955 VDDD.t936 VSUBS 0.983097f
C8956 VDDD.t1116 VSUBS 0.681305f
C8957 VDDD.t353 VSUBS 1.60497f
C8958 VDDD.t816 VSUBS 1.64155f
C8959 VDDD.t532 VSUBS 0.873355f
C8960 VDDD.t352 VSUBS 1.09284f
C8961 VDDD.t646 VSUBS 1.08369f
C8962 VDDD.t624 VSUBS 1.34432f
C8963 VDDD.t682 VSUBS 1.35346f
C8964 VDDD.t764 VSUBS 0.845919f
C8965 VDDD.t531 VSUBS 0.777344f
C8966 VDDD.t105 VSUBS 0.877942f
C8967 VDDD.t292 VSUBS 0.877942f
C8968 VDDD.t101 VSUBS 1.3672f
C8969 VDDD.t103 VSUBS 1.3672f
C8970 VDDD.t107 VSUBS 0.983097f
C8971 VDDD.t340 VSUBS 0.681305f
C8972 VDDD.t1205 VSUBS 1.60497f
C8973 VDDD.t375 VSUBS 1.64155f
C8974 VDDD.t1363 VSUBS 0.873355f
C8975 VDDD.t1330 VSUBS 1.09284f
C8976 VDDD.t135 VSUBS 1.08369f
C8977 VDDD.t776 VSUBS 1.34432f
C8978 VDDD.t420 VSUBS 1.35346f
C8979 VDDD.t1207 VSUBS 0.845919f
C8980 VDDD.t1364 VSUBS 0.777344f
C8981 VDDD.t525 VSUBS 0.877942f
C8982 VDDD.t179 VSUBS 0.877942f
C8983 VDDD.t438 VSUBS 1.3672f
C8984 VDDD.t231 VSUBS 1.3672f
C8985 VDDD.t527 VSUBS 0.983097f
C8986 VDDD.t323 VSUBS 1.30318f
C8987 VDDD.n2265 VSUBS 0.427239f
C8988 VDDD.n2267 VSUBS 0.61245f
C8989 VDDD.n2268 VSUBS 1.01164f
C8990 VDDD.n2269 VSUBS 0.118956f
C8991 VDDD.n2270 VSUBS 0.118956f
C8992 VDDD.n2271 VSUBS 0.128849f
C8993 VDDD.n2272 VSUBS 1.00123f
C8994 VDDD.t324 VSUBS 0.306452f
C8995 VDDD.n2273 VSUBS 0.359955f
C8996 VDDD.n2274 VSUBS 0.046011f
C8997 VDDD.n2275 VSUBS 0.187166f
C8998 VDDD.n2276 VSUBS 0.188716f
C8999 VDDD.n2277 VSUBS 0.251622f
C9000 VDDD.n2278 VSUBS 0.057151f
C9001 VDDD.n2279 VSUBS 0.521062f
C9002 VDDD.n2280 VSUBS 0.032934f
C9003 VDDD.n2281 VSUBS 0.226774f
C9004 VDDD.n2282 VSUBS 0.05037f
C9005 VDDD.n2283 VSUBS 0.251622f
C9006 VDDD.n2284 VSUBS 0.251622f
C9007 VDDD.n2285 VSUBS 0.251622f
C9008 VDDD.n2286 VSUBS 0.070712f
C9009 VDDD.n2287 VSUBS 0.089116f
C9010 VDDD.n2288 VSUBS 0.085726f
C9011 VDDD.n2289 VSUBS 0.251622f
C9012 VDDD.n2290 VSUBS 0.251622f
C9013 VDDD.n2291 VSUBS 0.251622f
C9014 VDDD.n2292 VSUBS 0.056666f
C9015 VDDD.n2293 VSUBS 0.049401f
C9016 VDDD.n2294 VSUBS 0.235104f
C9017 VDDD.n2295 VSUBS 0.052307f
C9018 VDDD.n2296 VSUBS 0.251622f
C9019 VDDD.n2297 VSUBS 0.251622f
C9020 VDDD.n2298 VSUBS 0.251622f
C9021 VDDD.n2299 VSUBS 0.089116f
C9022 VDDD.n2300 VSUBS 0.08621f
C9023 VDDD.n2301 VSUBS 0.250175f
C9024 VDDD.n2302 VSUBS 0.251622f
C9025 VDDD.n2303 VSUBS 0.251622f
C9026 VDDD.n2304 VSUBS 0.251622f
C9027 VDDD.n2305 VSUBS 0.074102f
C9028 VDDD.n2306 VSUBS 0.305072f
C9029 VDDD.n2307 VSUBS 0.062962f
C9030 VDDD.n2308 VSUBS 0.149059f
C9031 VDDD.n2309 VSUBS 0.188716f
C9032 VDDD.n2310 VSUBS 0.251622f
C9033 VDDD.n2311 VSUBS 0.057151f
C9034 VDDD.n2312 VSUBS 0.521062f
C9035 VDDD.n2313 VSUBS 0.032934f
C9036 VDDD.n2314 VSUBS 0.226774f
C9037 VDDD.n2315 VSUBS 0.05037f
C9038 VDDD.n2316 VSUBS 0.251622f
C9039 VDDD.n2317 VSUBS 0.251622f
C9040 VDDD.n2318 VSUBS 0.251622f
C9041 VDDD.n2319 VSUBS 0.070712f
C9042 VDDD.n2320 VSUBS 0.089116f
C9043 VDDD.n2321 VSUBS 0.085726f
C9044 VDDD.n2322 VSUBS 0.251622f
C9045 VDDD.n2323 VSUBS 0.251622f
C9046 VDDD.n2324 VSUBS 0.251622f
C9047 VDDD.n2325 VSUBS 0.056666f
C9048 VDDD.n2326 VSUBS 0.049401f
C9049 VDDD.n2327 VSUBS 0.235104f
C9050 VDDD.n2328 VSUBS 0.052307f
C9051 VDDD.n2329 VSUBS 0.251622f
C9052 VDDD.n2330 VSUBS 0.251622f
C9053 VDDD.n2331 VSUBS 0.251622f
C9054 VDDD.n2332 VSUBS 0.089116f
C9055 VDDD.n2333 VSUBS 0.08621f
C9056 VDDD.n2334 VSUBS 0.250175f
C9057 VDDD.n2335 VSUBS 0.251622f
C9058 VDDD.n2336 VSUBS 0.251622f
C9059 VDDD.n2337 VSUBS 0.251622f
C9060 VDDD.n2338 VSUBS 0.074102f
C9061 VDDD.n2339 VSUBS 0.305072f
C9062 VDDD.n2340 VSUBS 0.062962f
C9063 VDDD.n2341 VSUBS 0.149059f
C9064 VDDD.n2342 VSUBS 0.188716f
C9065 VDDD.n2343 VSUBS 0.251622f
C9066 VDDD.n2344 VSUBS 0.057151f
C9067 VDDD.n2345 VSUBS 0.521062f
C9068 VDDD.n2346 VSUBS 0.032934f
C9069 VDDD.n2347 VSUBS 0.226774f
C9070 VDDD.n2348 VSUBS 0.05037f
C9071 VDDD.n2349 VSUBS 0.251622f
C9072 VDDD.n2350 VSUBS 0.251622f
C9073 VDDD.n2351 VSUBS 0.251622f
C9074 VDDD.n2352 VSUBS 0.070712f
C9075 VDDD.n2353 VSUBS 0.089116f
C9076 VDDD.n2354 VSUBS 0.085726f
C9077 VDDD.n2355 VSUBS 0.251622f
C9078 VDDD.n2356 VSUBS 0.251622f
C9079 VDDD.n2357 VSUBS 0.251622f
C9080 VDDD.n2358 VSUBS 0.056666f
C9081 VDDD.n2359 VSUBS 0.049401f
C9082 VDDD.n2360 VSUBS 0.235104f
C9083 VDDD.n2361 VSUBS 0.052307f
C9084 VDDD.n2362 VSUBS 0.251622f
C9085 VDDD.n2363 VSUBS 0.251622f
C9086 VDDD.n2364 VSUBS 0.251622f
C9087 VDDD.n2365 VSUBS 0.089116f
C9088 VDDD.n2366 VSUBS 0.08621f
C9089 VDDD.n2367 VSUBS 0.250175f
C9090 VDDD.n2368 VSUBS 0.251622f
C9091 VDDD.n2369 VSUBS 0.251622f
C9092 VDDD.n2370 VSUBS 0.251622f
C9093 VDDD.n2371 VSUBS 0.074102f
C9094 VDDD.n2372 VSUBS 0.305072f
C9095 VDDD.n2373 VSUBS 0.062962f
C9096 VDDD.n2374 VSUBS 0.149059f
C9097 VDDD.n2375 VSUBS 0.188716f
C9098 VDDD.n2376 VSUBS 0.251622f
C9099 VDDD.n2377 VSUBS 0.057151f
C9100 VDDD.n2378 VSUBS 0.521062f
C9101 VDDD.n2379 VSUBS 0.032934f
C9102 VDDD.n2380 VSUBS 0.226774f
C9103 VDDD.n2381 VSUBS 0.05037f
C9104 VDDD.n2382 VSUBS 0.251622f
C9105 VDDD.n2383 VSUBS 0.251622f
C9106 VDDD.n2384 VSUBS 0.251622f
C9107 VDDD.n2385 VSUBS 0.070712f
C9108 VDDD.n2386 VSUBS 0.089116f
C9109 VDDD.n2387 VSUBS 0.085726f
C9110 VDDD.n2388 VSUBS 0.251622f
C9111 VDDD.n2389 VSUBS 0.251622f
C9112 VDDD.n2390 VSUBS 0.251622f
C9113 VDDD.n2391 VSUBS 0.056666f
C9114 VDDD.n2392 VSUBS 0.049401f
C9115 VDDD.n2393 VSUBS 0.235104f
C9116 VDDD.n2394 VSUBS 0.052307f
C9117 VDDD.n2395 VSUBS 0.251622f
C9118 VDDD.n2396 VSUBS 0.251622f
C9119 VDDD.n2397 VSUBS 0.251622f
C9120 VDDD.n2398 VSUBS 0.089116f
C9121 VDDD.n2399 VSUBS 0.08621f
C9122 VDDD.n2400 VSUBS 0.250175f
C9123 VDDD.n2401 VSUBS 0.251622f
C9124 VDDD.n2402 VSUBS 0.251622f
C9125 VDDD.n2403 VSUBS 0.251622f
C9126 VDDD.n2404 VSUBS 0.074102f
C9127 VDDD.n2405 VSUBS 0.305072f
C9128 VDDD.n2406 VSUBS 0.062962f
C9129 VDDD.n2407 VSUBS 0.149059f
C9130 VDDD.n2408 VSUBS 0.188716f
C9131 VDDD.n2409 VSUBS 0.251622f
C9132 VDDD.n2410 VSUBS 0.057151f
C9133 VDDD.n2411 VSUBS 0.521062f
C9134 VDDD.n2412 VSUBS 0.032934f
C9135 VDDD.n2413 VSUBS 0.226774f
C9136 VDDD.n2414 VSUBS 0.05037f
C9137 VDDD.n2415 VSUBS 0.251622f
C9138 VDDD.n2416 VSUBS 0.251622f
C9139 VDDD.n2417 VSUBS 0.251622f
C9140 VDDD.n2418 VSUBS 0.070712f
C9141 VDDD.n2419 VSUBS 0.089116f
C9142 VDDD.n2420 VSUBS 0.085726f
C9143 VDDD.n2421 VSUBS 0.251622f
C9144 VDDD.n2422 VSUBS 0.251622f
C9145 VDDD.n2423 VSUBS 0.251622f
C9146 VDDD.n2424 VSUBS 0.056666f
C9147 VDDD.n2425 VSUBS 0.049401f
C9148 VDDD.n2426 VSUBS 0.235104f
C9149 VDDD.n2427 VSUBS 0.052307f
C9150 VDDD.n2428 VSUBS 0.251622f
C9151 VDDD.n2429 VSUBS 0.251622f
C9152 VDDD.n2430 VSUBS 0.251622f
C9153 VDDD.n2431 VSUBS 0.089116f
C9154 VDDD.n2432 VSUBS 0.08621f
C9155 VDDD.n2433 VSUBS 0.250175f
C9156 VDDD.n2434 VSUBS 0.251622f
C9157 VDDD.n2435 VSUBS 0.251622f
C9158 VDDD.n2436 VSUBS 0.251622f
C9159 VDDD.n2437 VSUBS 0.074102f
C9160 VDDD.n2438 VSUBS 0.305072f
C9161 VDDD.n2439 VSUBS 0.062962f
C9162 VDDD.n2440 VSUBS 0.149059f
C9163 VDDD.n2441 VSUBS 0.188716f
C9164 VDDD.n2442 VSUBS 0.251622f
C9165 VDDD.n2443 VSUBS 0.057151f
C9166 VDDD.n2444 VSUBS 0.521062f
C9167 VDDD.n2445 VSUBS 0.032934f
C9168 VDDD.n2446 VSUBS 0.251622f
C9169 VDDD.n2447 VSUBS 0.251622f
C9170 VDDD.n2448 VSUBS 0.05037f
C9171 VDDD.n2449 VSUBS 0.24113f
C9172 VDDD.n2450 VSUBS 0.070712f
C9173 VDDD.n2451 VSUBS 0.251622f
C9174 VDDD.n2452 VSUBS 0.251622f
C9175 VDDD.n2453 VSUBS 0.251622f
C9176 VDDD.n2454 VSUBS 0.085726f
C9177 VDDD.n2455 VSUBS 0.3381f
C9178 VDDD.n2456 VSUBS 0.056666f
C9179 VDDD.t182 VSUBS 0.032307f
C9180 VDDD.t509 VSUBS 0.047863f
C9181 VDDD.n2457 VSUBS 0.083298f
C9182 VDDD.n2458 VSUBS 0.235104f
C9183 VDDD.n2459 VSUBS 0.049401f
C9184 VDDD.n2460 VSUBS 0.251622f
C9185 VDDD.n2461 VSUBS 0.251622f
C9186 VDDD.n2462 VSUBS 0.251622f
C9187 VDDD.n2463 VSUBS 0.089116f
C9188 VDDD.n2464 VSUBS 0.089116f
C9189 VDDD.n2465 VSUBS 0.08621f
C9190 VDDD.n2466 VSUBS 0.251622f
C9191 VDDD.n2467 VSUBS 0.251622f
C9192 VDDD.n2468 VSUBS 0.251622f
C9193 VDDD.n2469 VSUBS 0.067806f
C9194 VDDD.n2470 VSUBS 0.074102f
C9195 VDDD.n2471 VSUBS 0.326891f
C9196 VDDD.n2472 VSUBS 0.242239f
C9197 VDDD.n2473 VSUBS 1.45366f
C9198 VDDD.n2474 VSUBS 19.216301f
C9199 VDDD.n2475 VSUBS 11.2767f
C9200 VDDD.n2476 VSUBS 11.9215f
C9201 VDDD.n2477 VSUBS 1.03982f
C9202 VDDD.n2478 VSUBS 14.1446f
C9203 VDDD.n2479 VSUBS 8.08255f
C9204 VDDD.n2480 VSUBS 6.56975f
C9205 VDDD.n2481 VSUBS 20.4689f
C9206 VDDD.n2482 VSUBS 1.72508f
C9207 VDDD.n2483 VSUBS 6.642951f
C9208 VDDD.n2484 VSUBS 10.5557f
C9209 VDDD.n2485 VSUBS 1.72675f
C9210 VDDD.n2486 VSUBS 10.4828f
C9211 VDDD.n2487 VSUBS 15.842402f
C9212 VDDD.n2488 VSUBS 6.54685f
C9213 VDDD.n2489 VSUBS 9.120879f
C9214 VDDD.n2490 VSUBS 15.842402f
C9215 VDDD.n2491 VSUBS 11.0095f
C9216 VDDD.n2492 VSUBS 1.92558f
C9217 VDDD.t1369 VSUBS 1.66443f
C9218 VDDD.t1371 VSUBS 1.3672f
C9219 VDDD.t1110 VSUBS 1.3672f
C9220 VDDD.t488 VSUBS 0.877942f
C9221 VDDD.t601 VSUBS 0.877942f
C9222 VDDD.t858 VSUBS 0.777344f
C9223 VDDD.t18 VSUBS 0.845919f
C9224 VDDD.t1235 VSUBS 1.35346f
C9225 VDDD.t1219 VSUBS 1.34432f
C9226 VDDD.t540 VSUBS 1.08369f
C9227 VDDD.t109 VSUBS 1.09284f
C9228 VDDD.t65 VSUBS 0.873355f
C9229 VDDD.t1450 VSUBS 1.64155f
C9230 VDDD.t19 VSUBS 1.60497f
C9231 VDDD.t284 VSUBS 0.681305f
C9232 VDDD.t1146 VSUBS 0.983097f
C9233 VDDD.t1144 VSUBS 1.3672f
C9234 VDDD.t931 VSUBS 1.3672f
C9235 VDDD.t311 VSUBS 0.877942f
C9236 VDDD.t897 VSUBS 0.877942f
C9237 VDDD.t934 VSUBS 0.777344f
C9238 VDDD.t1104 VSUBS 0.845919f
C9239 VDDD.t1081 VSUBS 1.35346f
C9240 VDDD.t615 VSUBS 1.34432f
C9241 VDDD.t611 VSUBS 1.08369f
C9242 VDDD.t1297 VSUBS 1.09284f
C9243 VDDD.t935 VSUBS 0.873355f
C9244 VDDD.t97 VSUBS 1.64155f
C9245 VDDD.t1102 VSUBS 1.60497f
C9246 VDDD.t644 VSUBS 0.681305f
C9247 VDDD.t754 VSUBS 0.983097f
C9248 VDDD.t699 VSUBS 1.3672f
C9249 VDDD.t255 VSUBS 1.3672f
C9250 VDDD.t1268 VSUBS 0.877942f
C9251 VDDD.t701 VSUBS 0.877942f
C9252 VDDD.t1182 VSUBS 0.777344f
C9253 VDDD.t916 VSUBS 0.845919f
C9254 VDDD.t1227 VSUBS 1.35346f
C9255 VDDD.t500 VSUBS 1.34432f
C9256 VDDD.t1298 VSUBS 1.08369f
C9257 VDDD.t151 VSUBS 1.09284f
C9258 VDDD.t233 VSUBS 0.873355f
C9259 VDDD.t662 VSUBS 1.64155f
C9260 VDDD.t152 VSUBS 1.60497f
C9261 VDDD.t983 VSUBS 0.681305f
C9262 VDDD.t1384 VSUBS 0.983097f
C9263 VDDD.t34 VSUBS 1.3672f
C9264 VDDD.t562 VSUBS 1.3672f
C9265 VDDD.t819 VSUBS 0.877942f
C9266 VDDD.t32 VSUBS 0.877942f
C9267 VDDD.t610 VSUBS 0.777344f
C9268 VDDD.t1079 VSUBS 0.845919f
C9269 VDDD.t259 VSUBS 1.35346f
C9270 VDDD.t823 VSUBS 1.34432f
C9271 VDDD.t835 VSUBS 1.08369f
C9272 VDDD.t1080 VSUBS 1.09284f
C9273 VDDD.t790 VSUBS 0.873355f
C9274 VDDD.t237 VSUBS 1.64155f
C9275 VDDD.t209 VSUBS 1.60497f
C9276 VDDD.t131 VSUBS 0.681305f
C9277 VDDD.t1423 VSUBS 0.983097f
C9278 VDDD.t1011 VSUBS 1.3672f
C9279 VDDD.t1159 VSUBS 1.3672f
C9280 VDDD.t1187 VSUBS 0.877942f
C9281 VDDD.t1013 VSUBS 0.877942f
C9282 VDDD.t740 VSUBS 0.777344f
C9283 VDDD.t1405 VSUBS 0.845919f
C9284 VDDD.t1066 VSUBS 1.35346f
C9285 VDDD.t465 VSUBS 1.34432f
C9286 VDDD.t1337 VSUBS 1.08369f
C9287 VDDD.t1402 VSUBS 1.09284f
C9288 VDDD.t96 VSUBS 0.873355f
C9289 VDDD.t416 VSUBS 1.64155f
C9290 VDDD.t1403 VSUBS 1.60497f
C9291 VDDD.t537 VSUBS 0.681305f
C9292 VDDD.t219 VSUBS 0.983097f
C9293 VDDD.t217 VSUBS 1.3672f
C9294 VDDD.t550 VSUBS 1.3672f
C9295 VDDD.t1217 VSUBS 0.877942f
C9296 VDDD.t909 VSUBS 0.877942f
C9297 VDDD.t738 VSUBS 0.777344f
C9298 VDDD.t1395 VSUBS 0.845919f
C9299 VDDD.t434 VSUBS 1.35346f
C9300 VDDD.t1215 VSUBS 1.34432f
C9301 VDDD.t889 VSUBS 1.08369f
C9302 VDDD.t1394 VSUBS 1.09284f
C9303 VDDD.t739 VSUBS 0.873355f
C9304 VDDD.t99 VSUBS 1.64155f
C9305 VDDD.t760 VSUBS 1.60497f
C9306 VDDD.t2 VSUBS 0.681305f
C9307 VDDD.t92 VSUBS 0.983097f
C9308 VDDD.t90 VSUBS 1.3672f
C9309 VDDD.t991 VSUBS 1.3672f
C9310 VDDD.t914 VSUBS 0.877942f
C9311 VDDD.t243 VSUBS 0.877942f
C9312 VDDD.t1225 VSUBS 0.777344f
C9313 VDDD.t436 VSUBS 0.845919f
C9314 VDDD.t61 VSUBS 1.35346f
C9315 VDDD.t1316 VSUBS 1.34432f
C9316 VDDD.t529 VSUBS 1.08369f
C9317 VDDD.t1277 VSUBS 1.09284f
C9318 VDDD.t1226 VSUBS 0.873355f
C9319 VDDD.t235 VSUBS 1.64155f
C9320 VDDD.t58 VSUBS 1.60497f
C9321 VDDD.t1291 VSUBS 0.681305f
C9322 VDDD.t1349 VSUBS 0.983097f
C9323 VDDD.t1335 VSUBS 1.3672f
C9324 VDDD.t1154 VSUBS 1.3672f
C9325 VDDD.t486 VSUBS 0.877942f
C9326 VDDD.t397 VSUBS 0.877942f
C9327 VDDD.t593 VSUBS 0.777344f
C9328 VDDD.t1157 VSUBS 0.845919f
C9329 VDDD.t1073 VSUBS 1.35346f
C9330 VDDD.t899 VSUBS 1.34432f
C9331 VDDD.t797 VSUBS 1.08369f
C9332 VDDD.t1158 VSUBS 1.09284f
C9333 VDDD.t767 VSUBS 0.873355f
C9334 VDDD.t36 VSUBS 1.64155f
C9335 VDDD.t833 VSUBS 1.60497f
C9336 VDDD.t667 VSUBS 0.681305f
C9337 VDDD.t748 VSUBS 0.983097f
C9338 VDDD.t861 VSUBS 1.3672f
C9339 VDDD.t1457 VSUBS 1.3672f
C9340 VDDD.t492 VSUBS 0.877942f
C9341 VDDD.t928 VSUBS 0.877942f
C9342 VDDD.t1128 VSUBS 0.777344f
C9343 VDDD.t805 VSUBS 0.845919f
C9344 VDDD.t458 VSUBS 1.35346f
C9345 VDDD.t903 VSUBS 1.34432f
C9346 VDDD.t1378 VSUBS 1.08369f
C9347 VDDD.t804 VSUBS 1.09284f
C9348 VDDD.t148 VSUBS 0.873355f
C9349 VDDD.t660 VSUBS 1.64155f
C9350 VDDD.t806 VSUBS 1.60497f
C9351 VDDD.t84 VSUBS 0.681305f
C9352 VDDD.t160 VSUBS 0.983097f
C9353 VDDD.t1247 VSUBS 1.3672f
C9354 VDDD.t288 VSUBS 1.3672f
C9355 VDDD.t784 VSUBS 0.877942f
C9356 VDDD.t1245 VSUBS 0.877942f
C9357 VDDD.t144 VSUBS 0.777344f
C9358 VDDD.t794 VSUBS 0.845919f
C9359 VDDD.t381 VSUBS 1.35346f
C9360 VDDD.t630 VSUBS 1.34432f
C9361 VDDD.t1237 VSUBS 1.08369f
C9362 VDDD.t793 VSUBS 1.09284f
C9363 VDDD.t145 VSUBS 0.873355f
C9364 VDDD.t1452 VSUBS 1.64155f
C9365 VDDD.t125 VSUBS 1.60497f
C9366 VDDD.t975 VSUBS 0.681305f
C9367 VDDD.t269 VSUBS 1.29403f
C9368 VDDD.t887 VSUBS 0.768199f
C9369 VDDD.t410 VSUBS 0.768199f
C9370 VDDD.t271 VSUBS 0.768199f
C9371 VDDD.t185 VSUBS 0.768199f
C9372 VDDD.t211 VSUBS 0.768199f
C9373 VDDD.t885 VSUBS 0.768199f
C9374 VDDD.t187 VSUBS 0.768199f
C9375 VDDD.t665 VSUBS 0.768199f
C9376 VDDD.t926 VSUBS 0.768199f
C9377 VDDD.t924 VSUBS 0.676747f
.ends

