magic
tech sky130A
magscale 1 2
timestamp 1727883862
<< error_s >>
rect 2240 -306 2298 -300
rect 2556 -306 2614 -300
rect 2872 -306 2930 -300
rect 2240 -340 2252 -306
rect 2556 -340 2568 -306
rect 2872 -340 2884 -306
rect 2240 -346 2298 -340
rect 2556 -346 2614 -340
rect 2872 -346 2930 -340
rect 2240 -616 2298 -610
rect 2556 -616 2614 -610
rect 2872 -616 2930 -610
rect 2240 -650 2252 -616
rect 2556 -650 2568 -616
rect 2872 -650 2884 -616
rect 2240 -656 2298 -650
rect 2556 -656 2614 -650
rect 2872 -656 2930 -650
rect 2240 -820 2298 -814
rect 2556 -820 2614 -814
rect 2872 -820 2930 -814
rect 2240 -854 2252 -820
rect 2556 -854 2568 -820
rect 2872 -854 2884 -820
rect 2240 -860 2298 -854
rect 2556 -860 2614 -854
rect 2872 -860 2930 -854
rect 2240 -1130 2298 -1124
rect 2556 -1130 2614 -1124
rect 2872 -1130 2930 -1124
rect 2240 -1164 2252 -1130
rect 2556 -1164 2568 -1130
rect 2872 -1164 2884 -1130
rect 2240 -1170 2298 -1164
rect 2556 -1170 2614 -1164
rect 2872 -1170 2930 -1164
<< viali >>
rect -186 36 -28 70
rect 710 -414 744 -114
rect 2822 -752 2980 -718
rect -186 -1266 -28 -1232
rect 2190 -1266 2348 -1232
rect 2506 -1266 2664 -1232
rect 2822 -1266 2980 -1232
<< metal1 >>
rect -318 70 3112 106
rect -318 36 -186 70
rect -28 36 3112 70
rect -318 6 3112 36
rect -140 -75 -74 -22
rect -86 -413 34 -113
rect -140 -860 -74 -454
rect -16 -632 34 -413
rect 428 -114 478 6
rect 536 -83 602 -27
rect 852 -83 918 -27
rect 704 -114 750 -102
rect 428 -414 548 -114
rect 590 -414 710 -114
rect 744 -414 864 -114
rect 906 -126 1026 -114
rect 906 -402 958 -126
rect 1018 -402 1028 -126
rect 906 -414 1026 -402
rect 704 -426 750 -414
rect 526 -511 536 -445
rect 602 -511 612 -445
rect 852 -632 918 -445
rect 2290 -578 2390 -378
rect 2606 -578 2880 -378
rect 2922 -578 3076 -378
rect -16 -682 918 -632
rect -16 -892 34 -682
rect 2340 -892 2390 -578
rect 2810 -718 2992 -712
rect 3042 -718 3076 -578
rect 2810 -752 2822 -718
rect 2980 -752 3076 -718
rect 2810 -758 2992 -752
rect -86 -1092 34 -892
rect 2290 -1092 2564 -892
rect 2606 -1092 2880 -892
rect -140 -1174 -74 -1121
rect -318 -1232 3112 -1202
rect -318 -1266 -186 -1232
rect -28 -1266 2190 -1232
rect 2348 -1266 2506 -1232
rect 2664 -1266 2822 -1232
rect 2980 -1266 3112 -1232
rect -318 -1302 3112 -1266
<< via1 >>
rect 958 -402 1018 -126
rect 536 -511 602 -445
<< metal2 >>
rect 958 -126 1018 -116
rect 958 -435 1018 -402
rect 536 -445 1018 -435
rect 602 -511 1018 -445
rect 536 -521 1018 -511
<< metal3 >>
rect 667 -402 677 -302
rect 777 -402 787 -302
<< via3 >>
rect 677 -402 777 -302
<< metal4 >>
rect 676 -302 1273 -301
rect 676 -402 677 -302
rect 777 -402 1273 -302
rect 676 -403 1273 -402
use sky130_fd_pr__cap_mim_m3_1_K22CKP  sky130_fd_pr__cap_mim_m3_1_K22CKP_0
timestamp 1727309470
transform 0 1 1417 -1 0 -608
box -386 -240 386 240
use sky130_fd_pr__pfet_01v8_J4PGPS  XM1
timestamp 1727882782
transform 1 0 -107 0 1 -263
box -211 -369 211 369
use sky130_fd_pr__pfet_01v8_J4PGPS  XM2
timestamp 1727882782
transform 1 0 569 0 1 -264
box -211 -369 211 369
use sky130_fd_pr__pfet_01v8_J4PGPS  XM3
timestamp 1727882782
transform 1 0 885 0 1 -264
box -211 -369 211 369
use sky130_fd_pr__nfet_01v8_TGNW9T  XM4
timestamp 1727882782
transform 1 0 -107 0 1 -992
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM5
timestamp 1727882782
transform 1 0 2269 0 1 -992
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM6
timestamp 1727882782
transform 1 0 2269 0 1 -478
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM7
timestamp 1727882782
transform -1 0 2585 0 1 -992
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM8
timestamp 1727882782
transform -1 0 2585 0 1 -478
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM9
timestamp 1727882782
transform -1 0 2901 0 1 -478
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM10
timestamp 1727882782
transform 1 0 2901 0 1 -992
box -211 -310 211 310
<< end >>
