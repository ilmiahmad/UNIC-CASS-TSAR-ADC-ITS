magic
tech sky130A
magscale 1 2
timestamp 1730816635
<< dnwell >>
rect -16839 -13632 17921 4899
<< nwell >>
rect -16919 4693 18001 4979
rect -16919 -13426 -16633 4693
rect 17715 -13426 18001 4693
rect -16919 -13712 18001 -13426
<< nsubdiff >>
rect -16882 4922 17964 4942
rect -16882 4888 -16802 4922
rect 17884 4888 17964 4922
rect -16882 4868 17964 4888
rect -16882 4862 -16808 4868
rect -16882 -13595 -16862 4862
rect -16828 -13595 -16808 4862
rect -16882 -13601 -16808 -13595
rect 17890 4862 17964 4868
rect 17890 -13595 17910 4862
rect 17944 -13595 17964 4862
rect 17890 -13601 17964 -13595
rect -16882 -13621 17964 -13601
rect -16882 -13655 -16802 -13621
rect 17884 -13655 17964 -13621
rect -16882 -13675 17964 -13655
<< nsubdiffcont >>
rect -16802 4888 17884 4922
rect -16862 -13595 -16828 4862
rect 17910 -13595 17944 4862
rect -16802 -13655 17884 -13621
<< locali >>
rect -16862 4888 -16802 4922
rect 17884 4888 17944 4922
rect -16862 4862 -16828 4888
rect 17910 4862 17944 4888
rect -16862 -13621 -16828 -13595
rect 17910 -13621 17944 -13595
rect -16862 -13655 -16802 -13621
rect 17884 -13655 17944 -13621
<< viali >>
rect -16556 4922 -16456 4956
rect -16156 4922 -16056 4956
rect -15756 4922 -15656 4956
rect -16556 4888 -16456 4922
rect -16156 4888 -16056 4922
rect -15756 4888 -15656 4922
rect -16556 4856 -16456 4888
rect -16156 4856 -16056 4888
rect -15756 4856 -15656 4888
rect -16556 -13621 -16456 -13588
rect -16156 -13621 -16056 -13588
rect -15756 -13621 -15656 -13588
rect -16556 -13655 -16456 -13621
rect -16156 -13655 -16056 -13621
rect -15756 -13655 -15656 -13621
rect -16556 -13688 -16456 -13655
rect -16156 -13688 -16056 -13655
rect -15756 -13688 -15656 -13655
<< metal1 >>
rect -16568 4956 -16444 4962
rect -16568 4856 -16556 4956
rect -16456 4856 -16444 4956
rect -16568 4850 -16444 4856
rect -16168 4956 -16044 4962
rect -16168 4856 -16156 4956
rect -16056 4856 -16044 4956
rect -16168 4850 -16044 4856
rect -15768 4956 -15644 4962
rect -15768 4856 -15756 4956
rect -15656 4856 -15644 4956
rect -15768 4850 -15644 4856
rect -16566 4006 -16556 4102
rect -16460 4006 -16155 4102
rect -16059 4006 -15754 4102
rect -15658 4006 -1879 4102
rect -14945 2947 -14935 2999
rect -14883 2947 -2204 2999
rect -2152 2947 -2142 2999
rect -15346 2811 -15334 2863
rect -15282 2811 -2206 2863
rect -2154 2811 -2144 2863
rect -16365 1782 -16355 1878
rect -16259 1782 -15954 1878
rect -15858 1782 -15556 1878
rect -15460 1782 -1976 1878
rect -14543 1568 -14533 1620
rect -14481 1568 2710 1620
rect 2762 1568 2772 1620
rect -14741 1420 -14731 1472
rect -14679 1420 2862 1472
rect 2914 1420 2924 1472
rect 2317 173 2327 225
rect 2379 173 11350 225
rect 11402 173 11412 225
rect 4247 54 4257 106
rect 4309 54 11548 106
rect 11600 54 11610 106
rect 6179 -77 6189 -25
rect 6241 -77 11755 -25
rect 11807 -77 11817 -25
rect 8111 -198 8121 -145
rect 8174 -198 11940 -145
rect 11993 -198 12003 -145
rect 9699 -301 9709 -248
rect 9761 -301 12156 -248
rect 12209 -301 12219 -248
rect -16552 -545 -16542 -484
rect -16481 -545 -16144 -484
rect -16083 -545 -15750 -484
rect -15689 -545 225 -484
rect -15358 -667 -15333 -601
rect -15267 -667 -1144 -601
rect -1078 -667 -1068 -601
rect -14947 -816 -14937 -755
rect -14876 -816 -1121 -755
rect -1060 -816 -1050 -755
rect -14541 -939 -14531 -878
rect -14470 -939 -1111 -878
rect -1050 -939 -1040 -878
rect -16367 -1124 -16357 -1028
rect -16261 -1124 -15956 -1028
rect -15860 -1124 -15556 -1028
rect -15460 -1124 -989 -1028
rect -15148 -1342 -15138 -1282
rect -15078 -1287 -15012 -1282
rect -15078 -1338 -938 -1287
rect -15078 -1342 -15012 -1338
rect -16565 -1668 -16555 -1572
rect -16459 -1668 -16155 -1572
rect -16059 -1668 -15756 -1572
rect -15660 -1668 -1028 -1572
rect 7599 -1940 7609 -1888
rect 7661 -1940 12346 -1888
rect 12398 -1940 12408 -1888
rect 5669 -2068 5679 -2016
rect 5731 -2068 12555 -2016
rect 12607 -2068 12617 -2016
rect 3737 -2191 3747 -2139
rect 3799 -2191 12755 -2139
rect 12807 -2191 12817 -2139
rect 1805 -2320 1815 -2268
rect 1867 -2320 12950 -2268
rect 13002 -2320 13012 -2268
rect 229 -2441 239 -2389
rect 291 -2441 13151 -2389
rect 13203 -2441 13213 -2389
rect -16366 -4631 -16356 -4535
rect -16260 -4631 -15955 -4535
rect -15859 -4631 -15553 -4535
rect -15457 -4631 -377 -4535
rect -15344 -4782 -15334 -4718
rect -15270 -4782 -670 -4718
rect -606 -4782 -596 -4718
rect -14937 -4902 -14927 -4843
rect -14868 -4902 -651 -4843
rect -592 -4902 -582 -4843
rect -16565 -5175 -16555 -5079
rect -16459 -5175 -16156 -5079
rect -16060 -5175 -15754 -5079
rect -15658 -5175 -373 -5079
rect -16368 -5719 -16358 -5623
rect -16262 -5719 -15952 -5623
rect -15856 -5719 -15553 -5623
rect -15457 -5719 -380 -5623
rect 17516 -7172 17526 -7138
rect -11115 -7206 17526 -7172
rect -11115 -9752 -11081 -7206
rect 17516 -7238 17526 -7206
rect 17626 -7238 17636 -7138
rect 17316 -7300 17326 -7272
rect -10791 -7334 17326 -7300
rect -10791 -9310 -10757 -7334
rect 17316 -7372 17326 -7334
rect 17426 -7372 17436 -7272
rect 1326 -7572 1336 -7568
rect -7562 -7630 -7552 -7572
rect -7494 -7628 1336 -7572
rect 1396 -7572 1406 -7568
rect 1396 -7628 15149 -7572
rect -7494 -7630 15149 -7628
rect 15207 -7630 15217 -7572
rect 8 -7696 18 -7692
rect -5630 -7754 -5620 -7696
rect -5562 -7752 18 -7696
rect 78 -7696 88 -7692
rect 78 -7752 14942 -7696
rect -5562 -7754 14942 -7752
rect 15000 -7754 15010 -7696
rect 3258 -7824 3268 -7821
rect -3698 -7882 -3688 -7824
rect -3630 -7881 3268 -7824
rect 3328 -7824 3338 -7821
rect 3328 -7881 14741 -7824
rect -3630 -7882 14741 -7881
rect 14799 -7882 14809 -7824
rect 1942 -7983 1952 -7981
rect -1766 -8041 -1756 -7983
rect -1698 -8041 1952 -7983
rect 2012 -7983 2022 -7981
rect 2012 -8041 14550 -7983
rect 14608 -8041 14618 -7983
rect 5190 -8142 5200 -8139
rect 166 -8200 176 -8142
rect 234 -8199 5200 -8142
rect 5260 -8142 5270 -8139
rect 5260 -8199 14349 -8142
rect 234 -8200 14349 -8199
rect 14407 -8200 14417 -8142
rect 3872 -8260 3882 -8257
rect 2098 -8318 2108 -8260
rect 2166 -8317 3882 -8260
rect 3942 -8260 3952 -8257
rect 3942 -8317 14154 -8260
rect 2166 -8318 14154 -8317
rect 14212 -8318 14222 -8260
rect 4030 -8482 4040 -8424
rect 4098 -8427 13947 -8424
rect 4098 -8482 7130 -8427
rect 7120 -8487 7130 -8482
rect 7190 -8482 13947 -8427
rect 14005 -8482 14015 -8424
rect 7190 -8487 7200 -8482
rect 5804 -8603 5814 -8545
rect 5872 -8603 5972 -8545
rect 6030 -8603 13742 -8545
rect 13800 -8603 13810 -8545
rect 9054 -8656 9064 -8653
rect 7894 -8714 7904 -8656
rect 7962 -8713 9064 -8656
rect 9124 -8656 9134 -8653
rect 9124 -8713 13549 -8656
rect 7962 -8714 13549 -8713
rect 13607 -8714 13617 -8656
rect 7736 -8829 7746 -8769
rect 7806 -8771 7816 -8769
rect 7806 -8829 9836 -8771
rect 9894 -8829 13349 -8771
rect 13407 -8829 13417 -8771
rect -10497 -9019 -10487 -8939
rect -10404 -9019 -10394 -8939
rect -10430 -9569 -10420 -9489
rect -10337 -9569 -10327 -9489
rect -11115 -9786 -10757 -9752
rect -16555 -10123 -16545 -10043
rect -16465 -10123 -16148 -10043
rect -16068 -10123 -15751 -10043
rect -15671 -10123 -10404 -10043
rect 9826 -10286 9836 -10228
rect 9894 -10286 15349 -10228
rect 15407 -10286 15417 -10228
rect 7894 -10398 7904 -10340
rect 7962 -10398 15547 -10340
rect 15605 -10398 15615 -10340
rect 5962 -10511 5972 -10453
rect 6030 -10511 15746 -10453
rect 15804 -10511 15814 -10453
rect 4030 -10625 4040 -10567
rect 4098 -10625 15947 -10567
rect 16005 -10625 16015 -10567
rect 2098 -10734 2108 -10676
rect 2166 -10734 16147 -10676
rect 16205 -10734 16215 -10676
rect 166 -10872 176 -10814
rect 234 -10872 16351 -10814
rect 16409 -10872 16419 -10814
rect -1766 -10994 -1756 -10936
rect -1698 -10994 16547 -10936
rect 16605 -10994 16615 -10936
rect -3698 -11127 -3688 -11069
rect -3630 -11127 16749 -11069
rect 16807 -11127 16817 -11069
rect -5630 -11274 -5620 -11216
rect -5562 -11274 16951 -11216
rect 17009 -11274 17019 -11216
rect -7562 -11384 -7552 -11326
rect -7494 -11384 17148 -11326
rect 17206 -11384 17216 -11326
rect 8036 -11535 8046 -11477
rect 8104 -11535 13153 -11477
rect 13211 -11535 13221 -11477
rect 6104 -11658 6114 -11600
rect 6172 -11658 12946 -11600
rect 13004 -11658 13014 -11600
rect 4172 -11783 4182 -11725
rect 4240 -11783 12740 -11725
rect 12798 -11783 12808 -11725
rect 2240 -11912 2250 -11854
rect 2308 -11912 12554 -11854
rect 12612 -11912 12622 -11854
rect 308 -12041 318 -11983
rect 376 -12041 12348 -11983
rect 12406 -12041 12416 -11983
rect -1624 -12169 -1614 -12111
rect -1556 -12169 12166 -12111
rect 12224 -12169 12234 -12111
rect -3556 -12294 -3546 -12236
rect -3488 -12294 11952 -12236
rect 12010 -12294 12020 -12236
rect -5488 -12431 -5478 -12373
rect -5420 -12431 11748 -12373
rect 11806 -12431 11816 -12373
rect -7420 -12559 -7410 -12501
rect -7352 -12559 11549 -12501
rect 11607 -12559 11617 -12501
rect -9352 -12698 -9342 -12640
rect -9284 -12698 11352 -12640
rect 11410 -12698 11420 -12640
rect -16568 -13588 -16444 -13582
rect -16568 -13688 -16556 -13588
rect -16456 -13688 -16444 -13588
rect -16568 -13694 -16444 -13688
rect -16168 -13588 -16044 -13582
rect -16168 -13688 -16156 -13588
rect -16056 -13688 -16044 -13588
rect -16168 -13694 -16044 -13688
rect -15768 -13588 -15644 -13582
rect -15768 -13688 -15756 -13588
rect -15656 -13688 -15644 -13588
rect -15768 -13694 -15644 -13688
<< via1 >>
rect -16556 4856 -16456 4956
rect -16156 4856 -16056 4956
rect -15756 4856 -15656 4956
rect -16556 4006 -16460 4102
rect -16155 4006 -16059 4102
rect -15754 4006 -15658 4102
rect -14935 2947 -14883 2999
rect -2204 2947 -2152 2999
rect -15334 2811 -15282 2863
rect -2206 2811 -2154 2863
rect -16355 1782 -16259 1878
rect -15954 1782 -15858 1878
rect -15556 1782 -15460 1878
rect -14533 1568 -14481 1620
rect 2710 1568 2762 1620
rect -14731 1420 -14679 1472
rect 2862 1420 2914 1472
rect 2327 173 2379 225
rect 11350 173 11402 225
rect 4257 54 4309 106
rect 11548 54 11600 106
rect 6189 -77 6241 -25
rect 11755 -77 11807 -25
rect 8121 -198 8174 -145
rect 11940 -198 11993 -145
rect 9709 -301 9761 -248
rect 12156 -301 12209 -248
rect -16542 -545 -16481 -484
rect -16144 -545 -16083 -484
rect -15750 -545 -15689 -484
rect -15333 -667 -15267 -601
rect -1144 -667 -1078 -601
rect -14937 -816 -14876 -755
rect -1121 -816 -1060 -755
rect -14531 -939 -14470 -878
rect -1111 -939 -1050 -878
rect -16357 -1124 -16261 -1028
rect -15956 -1124 -15860 -1028
rect -15556 -1124 -15460 -1028
rect -15138 -1342 -15078 -1282
rect -16555 -1668 -16459 -1572
rect -16155 -1668 -16059 -1572
rect -15756 -1668 -15660 -1572
rect 7609 -1940 7661 -1888
rect 12346 -1940 12398 -1888
rect 5679 -2068 5731 -2016
rect 12555 -2068 12607 -2016
rect 3747 -2191 3799 -2139
rect 12755 -2191 12807 -2139
rect 1815 -2320 1867 -2268
rect 12950 -2320 13002 -2268
rect 239 -2441 291 -2389
rect 13151 -2441 13203 -2389
rect -16356 -4631 -16260 -4535
rect -15955 -4631 -15859 -4535
rect -15553 -4631 -15457 -4535
rect -15334 -4782 -15270 -4718
rect -670 -4782 -606 -4718
rect -14927 -4902 -14868 -4843
rect -651 -4902 -592 -4843
rect -16555 -5175 -16459 -5079
rect -16156 -5175 -16060 -5079
rect -15754 -5175 -15658 -5079
rect -16358 -5719 -16262 -5623
rect -15952 -5719 -15856 -5623
rect -15553 -5719 -15457 -5623
rect 17526 -7238 17626 -7138
rect 17326 -7372 17426 -7272
rect -7552 -7630 -7494 -7572
rect 1336 -7628 1396 -7568
rect 15149 -7630 15207 -7572
rect -5620 -7754 -5562 -7696
rect 18 -7752 78 -7692
rect 14942 -7754 15000 -7696
rect -3688 -7882 -3630 -7824
rect 3268 -7881 3328 -7821
rect 14741 -7882 14799 -7824
rect -1756 -8041 -1698 -7983
rect 1952 -8041 2012 -7981
rect 14550 -8041 14608 -7983
rect 176 -8200 234 -8142
rect 5200 -8199 5260 -8139
rect 14349 -8200 14407 -8142
rect 2108 -8318 2166 -8260
rect 3882 -8317 3942 -8257
rect 14154 -8318 14212 -8260
rect 4040 -8482 4098 -8424
rect 7130 -8487 7190 -8427
rect 13947 -8482 14005 -8424
rect 5814 -8603 5872 -8545
rect 5972 -8603 6030 -8545
rect 13742 -8603 13800 -8545
rect 7904 -8714 7962 -8656
rect 9064 -8713 9124 -8653
rect 13549 -8714 13607 -8656
rect 7746 -8829 7806 -8769
rect 9836 -8829 9894 -8771
rect 13349 -8829 13407 -8771
rect -10487 -9019 -10404 -8939
rect -10420 -9569 -10337 -9489
rect -16545 -10123 -16465 -10043
rect -16148 -10123 -16068 -10043
rect -15751 -10123 -15671 -10043
rect 9836 -10286 9894 -10228
rect 15349 -10286 15407 -10228
rect 7904 -10398 7962 -10340
rect 15547 -10398 15605 -10340
rect 5972 -10511 6030 -10453
rect 15746 -10511 15804 -10453
rect 4040 -10625 4098 -10567
rect 15947 -10625 16005 -10567
rect 2108 -10734 2166 -10676
rect 16147 -10734 16205 -10676
rect 176 -10872 234 -10814
rect 16351 -10872 16409 -10814
rect -1756 -10994 -1698 -10936
rect 16547 -10994 16605 -10936
rect -3688 -11127 -3630 -11069
rect 16749 -11127 16807 -11069
rect -5620 -11274 -5562 -11216
rect 16951 -11274 17009 -11216
rect -7552 -11384 -7494 -11326
rect 17148 -11384 17206 -11326
rect 8046 -11535 8104 -11477
rect 13153 -11535 13211 -11477
rect 6114 -11658 6172 -11600
rect 12946 -11658 13004 -11600
rect 4182 -11783 4240 -11725
rect 12740 -11783 12798 -11725
rect 2250 -11912 2308 -11854
rect 12554 -11912 12612 -11854
rect 318 -12041 376 -11983
rect 12348 -12041 12406 -11983
rect -1614 -12169 -1556 -12111
rect 12166 -12169 12224 -12111
rect -3546 -12294 -3488 -12236
rect 11952 -12294 12010 -12236
rect -5478 -12431 -5420 -12373
rect 11748 -12431 11806 -12373
rect -7410 -12559 -7352 -12501
rect 11549 -12559 11607 -12501
rect -9342 -12698 -9284 -12640
rect 11352 -12698 11410 -12640
rect -16556 -13688 -16456 -13588
rect -16156 -13688 -16056 -13588
rect -15756 -13688 -15656 -13588
<< metal2 >>
rect -16556 4956 -16456 4966
rect -16556 4102 -16456 4856
rect -16156 4956 -16056 4966
rect -16460 4006 -16456 4102
rect -16556 -484 -16456 4006
rect -16556 -545 -16542 -484
rect -16481 -545 -16456 -484
rect -16556 -1572 -16456 -545
rect -16356 1878 -16256 4637
rect -16356 1782 -16355 1878
rect -16259 1782 -16256 1878
rect -16356 -1018 -16256 1782
rect -16357 -1028 -16256 -1018
rect -16261 -1124 -16256 -1028
rect -16357 -1134 -16256 -1124
rect -16556 -1668 -16555 -1572
rect -16459 -1668 -16456 -1572
rect -16556 -5079 -16456 -1668
rect -16556 -5175 -16555 -5079
rect -16459 -5175 -16456 -5079
rect -16556 -8939 -16456 -5175
rect -16356 -4535 -16256 -1134
rect -16260 -4631 -16256 -4535
rect -16356 -5613 -16256 -4631
rect -16358 -5623 -16256 -5613
rect -16262 -5719 -16256 -5623
rect -16358 -5729 -16256 -5719
rect -16556 -9019 -16548 -8939
rect -16468 -9019 -16456 -8939
rect -16556 -10043 -16456 -9019
rect -16556 -10123 -16545 -10043
rect -16465 -10123 -16456 -10043
rect -16556 -13588 -16456 -10123
rect -16356 -9573 -16256 -5729
rect -16356 -9653 -16345 -9573
rect -16265 -9653 -16256 -9573
rect -16356 -13385 -16256 -9653
rect -16156 4102 -16056 4856
rect -15756 4956 -15656 4966
rect -16156 4006 -16155 4102
rect -16059 4006 -16056 4102
rect -16156 -484 -16056 4006
rect -16156 -545 -16144 -484
rect -16083 -545 -16056 -484
rect -16156 -1572 -16056 -545
rect -16156 -1668 -16155 -1572
rect -16059 -1668 -16056 -1572
rect -16156 -5079 -16056 -1668
rect -16060 -5175 -16056 -5079
rect -16156 -8939 -16056 -5175
rect -16156 -9019 -16154 -8939
rect -16074 -9019 -16056 -8939
rect -16156 -10043 -16056 -9019
rect -16156 -10123 -16148 -10043
rect -16068 -10123 -16056 -10043
rect -16556 -13698 -16456 -13688
rect -16156 -13588 -16056 -10123
rect -15956 1878 -15856 4637
rect -15956 1782 -15954 1878
rect -15858 1782 -15856 1878
rect -15956 -1028 -15856 1782
rect -15860 -1124 -15856 -1028
rect -15956 -4535 -15856 -1124
rect -15956 -4631 -15955 -4535
rect -15859 -4631 -15856 -4535
rect -15956 -5623 -15856 -4631
rect -15956 -5719 -15952 -5623
rect -15956 -9573 -15856 -5719
rect -15956 -9653 -15946 -9573
rect -15866 -9653 -15856 -9573
rect -15956 -13385 -15856 -9653
rect -15756 4102 -15656 4856
rect -15756 4006 -15754 4102
rect -15658 4006 -15656 4102
rect -15756 -484 -15656 4006
rect -15756 -545 -15750 -484
rect -15689 -545 -15656 -484
rect -15756 -1572 -15656 -545
rect -15660 -1668 -15656 -1572
rect -15756 -5079 -15656 -1668
rect -15756 -5175 -15754 -5079
rect -15658 -5175 -15656 -5079
rect -15756 -8939 -15656 -5175
rect -15676 -9019 -15656 -8939
rect -15756 -10043 -15656 -9019
rect -15756 -10123 -15751 -10043
rect -15671 -10123 -15656 -10043
rect -16156 -13698 -16056 -13688
rect -15756 -13588 -15656 -10123
rect -15556 1878 -15456 4637
rect -15460 1782 -15456 1878
rect -15556 -1028 -15456 1782
rect -15460 -1124 -15456 -1028
rect -15556 -4535 -15456 -1124
rect -15556 -4631 -15553 -4535
rect -15457 -4631 -15456 -4535
rect -15556 -5623 -15456 -4631
rect -15556 -5719 -15553 -5623
rect -15457 -5719 -15456 -5623
rect -15556 -9573 -15456 -5719
rect -15556 -9653 -15536 -9573
rect -15556 -13385 -15456 -9653
rect -15356 2863 -15256 4637
rect -15356 2811 -15334 2863
rect -15282 2811 -15256 2863
rect -15356 -601 -15256 2811
rect -15356 -667 -15333 -601
rect -15267 -667 -15256 -601
rect -15356 -4718 -15256 -667
rect -15356 -4782 -15334 -4718
rect -15270 -4782 -15256 -4718
rect -15356 -13385 -15256 -4782
rect -15156 -1282 -15056 4637
rect -15156 -1342 -15138 -1282
rect -15078 -1342 -15056 -1282
rect -15156 -13385 -15056 -1342
rect -14956 2999 -14856 4637
rect -14956 2947 -14935 2999
rect -14883 2947 -14856 2999
rect -14956 -755 -14856 2947
rect -14956 -816 -14937 -755
rect -14876 -816 -14856 -755
rect -14956 -4843 -14856 -816
rect -14956 -4902 -14927 -4843
rect -14868 -4902 -14856 -4843
rect -14956 -13385 -14856 -4902
rect -14756 1472 -14656 4637
rect -14756 1420 -14731 1472
rect -14679 1420 -14656 1472
rect -14756 -13385 -14656 1420
rect -14556 1620 -14456 4637
rect -14556 1568 -14533 1620
rect -14481 1568 -14456 1620
rect -14556 -878 -14456 1568
rect -14556 -939 -14531 -878
rect -14470 -939 -14456 -878
rect -14556 -9365 -14456 -939
rect -14356 -2810 -14256 4637
rect -14356 -2870 -14340 -2810
rect -14280 -2870 -14256 -2810
rect -14556 -9375 -14452 -9365
rect -14556 -9455 -14532 -9375
rect -14556 -9465 -14452 -9455
rect -14556 -13385 -14456 -9465
rect -14356 -13385 -14256 -2870
rect -14156 -2949 -14056 4637
rect -14156 -3009 -14132 -2949
rect -14072 -3009 -14056 -2949
rect -14156 -13385 -14056 -3009
rect -13956 -3088 -13856 4637
rect -13956 -3148 -13942 -3088
rect -13882 -3148 -13856 -3088
rect -13956 -13385 -13856 -3148
rect -13756 -3217 -13656 4637
rect -13756 -3277 -13734 -3217
rect -13674 -3277 -13656 -3217
rect -13756 -13385 -13656 -3277
rect -13556 -3356 -13456 4637
rect -13556 -3416 -13540 -3356
rect -13480 -3416 -13456 -3356
rect -13556 -13385 -13456 -3416
rect -13356 -3551 -13256 4637
rect -13356 -3611 -13331 -3551
rect -13271 -3611 -13256 -3551
rect -13356 -13385 -13256 -3611
rect -13156 -3726 -13056 4637
rect -13156 -3786 -13137 -3726
rect -13077 -3786 -13056 -3726
rect -13156 -13385 -13056 -3786
rect -12956 -3893 -12856 4637
rect -12956 -3953 -12938 -3893
rect -12878 -3953 -12856 -3893
rect -12956 -13385 -12856 -3953
rect -12756 -4046 -12656 4637
rect -12756 -4106 -12730 -4046
rect -12670 -4106 -12656 -4046
rect -12756 -13385 -12656 -4106
rect -12556 -4219 -12456 4637
rect -2204 2999 -2152 3009
rect -2204 2937 -2152 2947
rect -2206 2863 -2154 2873
rect -2206 2801 -2154 2811
rect 2695 2107 2914 2159
rect 2710 1620 2762 2039
rect 2710 1558 2762 1568
rect 2862 1472 2914 2107
rect 2862 1410 2914 1420
rect 2327 225 2379 235
rect 2327 -306 2379 173
rect 11326 225 11426 4637
rect 11326 173 11350 225
rect 11402 173 11426 225
rect 4257 106 4309 116
rect 4257 -326 4309 54
rect 6189 -25 6241 -15
rect 6189 -309 6241 -77
rect 8121 -145 8174 -135
rect 8121 -208 8174 -198
rect 8121 -272 8173 -208
rect 9709 -248 9761 -238
rect 9709 -311 9761 -301
rect -1144 -601 -1078 -591
rect -1078 -667 -1027 -601
rect -1144 -677 -1078 -667
rect -1121 -755 -1060 -745
rect -1060 -816 -1018 -755
rect -1121 -826 -1060 -816
rect -1111 -878 -1050 -868
rect -1050 -939 -1014 -878
rect -1111 -949 -1050 -939
rect 239 -2389 291 -1880
rect 1815 -2268 1867 -1880
rect 3747 -2139 3799 -1881
rect 7609 -1888 7661 -1878
rect 5679 -2016 5731 -1888
rect 7609 -1950 7661 -1940
rect 5679 -2078 5731 -2068
rect 3747 -2201 3799 -2191
rect 1815 -2330 1867 -2320
rect 239 -2451 291 -2441
rect -12556 -4279 -12540 -4219
rect -12480 -4279 -12456 -4219
rect -12556 -13385 -12456 -4279
rect -670 -4718 -606 -4708
rect -606 -4782 -558 -4718
rect -670 -4792 -606 -4782
rect -651 -4843 -592 -4833
rect -592 -4902 -558 -4843
rect -651 -4912 -592 -4902
rect 18 -5988 78 -5978
rect -7552 -7572 -7494 -7562
rect -7552 -8883 -7494 -7630
rect -5620 -7696 -5562 -7686
rect -5620 -8893 -5562 -7754
rect 18 -7692 78 -6048
rect 1336 -5988 1396 -5978
rect 1336 -7568 1396 -6048
rect 1336 -7638 1396 -7628
rect 1952 -5988 2012 -5978
rect 18 -7762 78 -7752
rect -3688 -7824 -3630 -7814
rect -3688 -8885 -3630 -7882
rect -1756 -7983 -1698 -7973
rect -1756 -8896 -1698 -8041
rect 1952 -7981 2012 -6048
rect 3268 -5988 3328 -5978
rect 3268 -7821 3328 -6048
rect 3268 -7891 3328 -7881
rect 3882 -5988 3942 -5978
rect 1952 -8051 2012 -8041
rect 176 -8142 234 -8132
rect 176 -8883 234 -8200
rect 2108 -8260 2166 -8250
rect 2108 -8904 2166 -8318
rect 3882 -8257 3942 -6048
rect 5200 -5988 5260 -5978
rect 5200 -8139 5260 -6048
rect 5200 -8209 5260 -8199
rect 5814 -5984 5874 -5974
rect 3882 -8327 3942 -8317
rect 4040 -8424 4098 -8414
rect 4040 -8874 4098 -8482
rect 5814 -8545 5874 -6044
rect 7130 -5988 7190 -5978
rect 7130 -8427 7190 -6048
rect 7130 -8497 7190 -8487
rect 7746 -5988 7806 -5978
rect 5872 -8591 5874 -8545
rect 5972 -8545 6030 -8535
rect 5814 -8613 5872 -8603
rect 5972 -8871 6030 -8603
rect 7746 -8769 7806 -6048
rect 9064 -5987 9124 -5977
rect 7746 -8839 7806 -8829
rect 7904 -8656 7962 -8646
rect 7904 -8874 7962 -8714
rect 9064 -8653 9124 -6047
rect 9064 -8723 9124 -8713
rect 9836 -8771 9894 -8761
rect 9836 -8871 9894 -8829
rect -10487 -8939 -10404 -8929
rect -10487 -9029 -10404 -9019
rect -10420 -9489 -10337 -9479
rect -10420 -9573 -10337 -9569
rect -10420 -9663 -10337 -9653
rect -9342 -12640 -9284 -10129
rect -7552 -11326 -7494 -10197
rect -7552 -11394 -7494 -11384
rect -7410 -12501 -7352 -10119
rect -5620 -11216 -5562 -10189
rect -5620 -11284 -5562 -11274
rect -5478 -12373 -5420 -10129
rect -3688 -11069 -3630 -10197
rect -3688 -11137 -3630 -11127
rect -3546 -12236 -3488 -10129
rect -1756 -10936 -1698 -10190
rect -1756 -11004 -1698 -10994
rect -1614 -12111 -1556 -10129
rect 176 -10814 234 -10195
rect 176 -10882 234 -10872
rect 318 -11983 376 -10129
rect 2108 -10676 2166 -10192
rect 2108 -10744 2166 -10734
rect 2250 -11854 2308 -10119
rect 4040 -10567 4098 -10193
rect 4040 -10635 4098 -10625
rect 4182 -11725 4240 -10129
rect 5972 -10453 6030 -10197
rect 5972 -10521 6030 -10511
rect 6114 -11600 6172 -10129
rect 7904 -10340 7962 -10191
rect 7904 -10408 7962 -10398
rect 8046 -11477 8104 -10116
rect 9836 -10228 9894 -10197
rect 9836 -10296 9894 -10286
rect 8046 -11545 8104 -11535
rect 6114 -11668 6172 -11658
rect 4182 -11793 4240 -11783
rect 2250 -11922 2308 -11912
rect 318 -12051 376 -12041
rect -1614 -12179 -1556 -12169
rect -3546 -12304 -3488 -12294
rect -5478 -12441 -5420 -12431
rect -7410 -12569 -7352 -12559
rect -9342 -12708 -9284 -12698
rect 11326 -12640 11426 173
rect 11326 -12698 11352 -12640
rect 11410 -12698 11426 -12640
rect 11326 -13385 11426 -12698
rect 11526 106 11626 4637
rect 11526 54 11548 106
rect 11600 54 11626 106
rect 11526 -12501 11626 54
rect 11526 -12559 11549 -12501
rect 11607 -12559 11626 -12501
rect 11526 -13385 11626 -12559
rect 11726 -25 11826 4637
rect 11726 -77 11755 -25
rect 11807 -77 11826 -25
rect 11726 -12373 11826 -77
rect 11726 -12431 11748 -12373
rect 11806 -12431 11826 -12373
rect 11726 -13385 11826 -12431
rect 11926 -145 12026 4637
rect 11926 -198 11940 -145
rect 11993 -198 12026 -145
rect 11926 -12236 12026 -198
rect 11926 -12294 11952 -12236
rect 12010 -12294 12026 -12236
rect 11926 -13385 12026 -12294
rect 12126 -248 12226 4637
rect 12126 -301 12156 -248
rect 12209 -301 12226 -248
rect 12126 -12111 12226 -301
rect 12126 -12169 12166 -12111
rect 12224 -12169 12226 -12111
rect 12126 -13385 12226 -12169
rect 12326 -1888 12426 4637
rect 12326 -1940 12346 -1888
rect 12398 -1940 12426 -1888
rect 12326 -11983 12426 -1940
rect 12326 -12041 12348 -11983
rect 12406 -12041 12426 -11983
rect 12326 -13385 12426 -12041
rect 12526 -2016 12626 4637
rect 12526 -2068 12555 -2016
rect 12607 -2068 12626 -2016
rect 12526 -11854 12626 -2068
rect 12526 -11912 12554 -11854
rect 12612 -11912 12626 -11854
rect 12526 -13385 12626 -11912
rect 12726 -2139 12826 4637
rect 12726 -2191 12755 -2139
rect 12807 -2191 12826 -2139
rect 12726 -11725 12826 -2191
rect 12726 -11783 12740 -11725
rect 12798 -11783 12826 -11725
rect 12726 -13385 12826 -11783
rect 12926 -2268 13026 4637
rect 12926 -2320 12950 -2268
rect 13002 -2320 13026 -2268
rect 12926 -11600 13026 -2320
rect 12926 -11658 12946 -11600
rect 13004 -11658 13026 -11600
rect 12926 -13385 13026 -11658
rect 13126 -2389 13226 4637
rect 13126 -2441 13151 -2389
rect 13203 -2441 13226 -2389
rect 13126 -11477 13226 -2441
rect 13126 -11535 13153 -11477
rect 13211 -11535 13226 -11477
rect 13126 -13385 13226 -11535
rect 13326 -8771 13426 4637
rect 13326 -8829 13349 -8771
rect 13407 -8829 13426 -8771
rect 13326 -13385 13426 -8829
rect 13526 -8656 13626 4637
rect 13526 -8714 13549 -8656
rect 13607 -8714 13626 -8656
rect 13526 -13385 13626 -8714
rect 13726 -8545 13826 4637
rect 13726 -8603 13742 -8545
rect 13800 -8603 13826 -8545
rect 13726 -13385 13826 -8603
rect 13926 -8424 14026 4637
rect 13926 -8482 13947 -8424
rect 14005 -8482 14026 -8424
rect 13926 -13385 14026 -8482
rect 14126 -8260 14226 4637
rect 14126 -8318 14154 -8260
rect 14212 -8318 14226 -8260
rect 14126 -13385 14226 -8318
rect 14326 -8142 14426 4637
rect 14326 -8200 14349 -8142
rect 14407 -8200 14426 -8142
rect 14326 -13385 14426 -8200
rect 14526 -7983 14626 4637
rect 14526 -8041 14550 -7983
rect 14608 -8041 14626 -7983
rect 14526 -13385 14626 -8041
rect 14726 -7824 14826 4637
rect 14726 -7882 14741 -7824
rect 14799 -7882 14826 -7824
rect 14726 -13385 14826 -7882
rect 14926 -7696 15026 4637
rect 14926 -7754 14942 -7696
rect 15000 -7754 15026 -7696
rect 14926 -13385 15026 -7754
rect 15126 -7572 15226 4637
rect 15126 -7630 15149 -7572
rect 15207 -7630 15226 -7572
rect 15126 -13385 15226 -7630
rect 15326 -10228 15426 4637
rect 15326 -10286 15349 -10228
rect 15407 -10286 15426 -10228
rect 15326 -13385 15426 -10286
rect 15526 -10340 15626 4637
rect 15526 -10398 15547 -10340
rect 15605 -10398 15626 -10340
rect 15526 -13385 15626 -10398
rect 15726 -10453 15826 4637
rect 15726 -10511 15746 -10453
rect 15804 -10511 15826 -10453
rect 15726 -13385 15826 -10511
rect 15926 -10567 16026 4637
rect 15926 -10625 15947 -10567
rect 16005 -10625 16026 -10567
rect 15926 -13385 16026 -10625
rect 16126 -10676 16226 4637
rect 16126 -10734 16147 -10676
rect 16205 -10734 16226 -10676
rect 16126 -13385 16226 -10734
rect 16326 -10814 16426 4637
rect 16326 -10872 16351 -10814
rect 16409 -10872 16426 -10814
rect 16326 -13385 16426 -10872
rect 16526 -10936 16626 4637
rect 16526 -10994 16547 -10936
rect 16605 -10994 16626 -10936
rect 16526 -13385 16626 -10994
rect 16726 -11069 16826 4637
rect 16726 -11127 16749 -11069
rect 16807 -11127 16826 -11069
rect 16726 -13385 16826 -11127
rect 16926 -11216 17026 4637
rect 16926 -11274 16951 -11216
rect 17009 -11274 17026 -11216
rect 16926 -13385 17026 -11274
rect 17126 -11326 17226 4637
rect 17126 -11384 17148 -11326
rect 17206 -11384 17226 -11326
rect 17126 -13385 17226 -11384
rect 17326 -7272 17426 4637
rect 17326 -13385 17426 -7372
rect 17526 -7138 17626 4637
rect 17526 -13385 17626 -7238
rect -15756 -13698 -15656 -13688
<< via2 >>
rect -16548 -9019 -16468 -8939
rect -16345 -9653 -16265 -9573
rect -16154 -9019 -16074 -8939
rect -15946 -9653 -15866 -9573
rect -15756 -9019 -15676 -8939
rect -15536 -9653 -15456 -9573
rect -14340 -2870 -14280 -2810
rect -14532 -9455 -14452 -9375
rect -14132 -3009 -14072 -2949
rect -13942 -3148 -13882 -3088
rect -13734 -3277 -13674 -3217
rect -13540 -3416 -13480 -3356
rect -13331 -3611 -13271 -3551
rect -13137 -3786 -13077 -3726
rect -12938 -3953 -12878 -3893
rect -12730 -4106 -12670 -4046
rect -12540 -4279 -12480 -4219
rect 18 -6048 78 -5988
rect 1336 -6048 1396 -5988
rect 1952 -6048 2012 -5988
rect 3268 -6048 3328 -5988
rect 3882 -6048 3942 -5988
rect 5200 -6048 5260 -5988
rect 5814 -6044 5874 -5984
rect 7130 -6048 7190 -5988
rect 7746 -6048 7806 -5988
rect 9064 -6047 9124 -5987
rect -10487 -9019 -10404 -8939
rect -10420 -9653 -10337 -9573
<< metal3 >>
rect -14350 -2810 -14270 -2805
rect -14350 -2870 -14340 -2810
rect -14280 -2870 9296 -2810
rect -14350 -2875 -14270 -2870
rect -14142 -2949 -14062 -2944
rect -14142 -3009 -14132 -2949
rect -14072 -3009 7640 -2949
rect -14142 -3014 -14062 -3009
rect -13952 -3088 -13872 -3083
rect -13952 -3148 -13942 -3088
rect -13882 -3148 7364 -3088
rect -13952 -3153 -13872 -3148
rect -13744 -3217 -13664 -3212
rect -13744 -3277 -13734 -3217
rect -13674 -3277 5702 -3217
rect -13744 -3282 -13664 -3277
rect -13550 -3356 -13470 -3351
rect -13550 -3416 -13540 -3356
rect -13480 -3416 5432 -3356
rect -13550 -3421 -13470 -3416
rect -13341 -3551 -13261 -3546
rect -13341 -3611 -13331 -3551
rect -13271 -3611 3771 -3551
rect -13341 -3616 -13261 -3611
rect -13147 -3726 -13067 -3721
rect -13147 -3786 -13137 -3726
rect -13077 -3786 3500 -3726
rect -13147 -3791 -13067 -3786
rect -12948 -3893 -12868 -3888
rect -12948 -3953 -12938 -3893
rect -12878 -3953 1839 -3893
rect -12948 -3958 -12868 -3953
rect -12740 -4046 -12660 -4041
rect -12740 -4106 -12730 -4046
rect -12670 -4106 1562 -4046
rect -12740 -4111 -12660 -4106
rect -12550 -4219 -12470 -4214
rect -12550 -4279 -12540 -4219
rect -12480 -4279 -93 -4219
rect -12550 -4284 -12470 -4279
rect 1502 -4291 1562 -4106
rect 1779 -4305 1839 -3953
rect 3440 -4310 3500 -3786
rect 3711 -4282 3771 -3611
rect 5372 -4388 5432 -3416
rect 5642 -4296 5702 -3277
rect 7304 -4356 7364 -3148
rect 7580 -4347 7640 -3009
rect 9236 -4310 9296 -2870
rect 8 -5988 88 -5983
rect 8 -6048 18 -5988
rect 78 -6048 88 -5988
rect 8 -6053 88 -6048
rect 1326 -5988 1406 -5983
rect 1326 -6048 1336 -5988
rect 1396 -6048 1406 -5988
rect 1326 -6053 1406 -6048
rect 1942 -5988 2022 -5983
rect 1942 -6048 1952 -5988
rect 2012 -6048 2022 -5988
rect 1942 -6053 2022 -6048
rect 3258 -5988 3338 -5983
rect 3258 -6048 3268 -5988
rect 3328 -6048 3338 -5988
rect 3258 -6053 3338 -6048
rect 3872 -5988 3952 -5983
rect 3872 -6048 3882 -5988
rect 3942 -6048 3952 -5988
rect 3872 -6053 3952 -6048
rect 5190 -5988 5270 -5983
rect 5190 -6048 5200 -5988
rect 5260 -6048 5270 -5988
rect 5190 -6053 5270 -6048
rect 5804 -5984 5884 -5979
rect 5804 -6044 5814 -5984
rect 5874 -6044 5884 -5984
rect 5804 -6049 5884 -6044
rect 7120 -5988 7200 -5983
rect 7120 -6048 7130 -5988
rect 7190 -6048 7200 -5988
rect 7120 -6053 7200 -6048
rect 7736 -5988 7816 -5983
rect 7736 -6048 7746 -5988
rect 7806 -6048 7816 -5988
rect 7736 -6053 7816 -6048
rect 9054 -5987 9134 -5982
rect 9054 -6047 9064 -5987
rect 9124 -6047 9134 -5987
rect 9054 -6052 9134 -6047
rect -16558 -8939 -16458 -8934
rect -16164 -8939 -16064 -8934
rect -15766 -8939 -15666 -8934
rect -10497 -8939 -10394 -8934
rect -16558 -9019 -16548 -8939
rect -16468 -9019 -16154 -8939
rect -16074 -9019 -15756 -8939
rect -15676 -9019 -10487 -8939
rect -10404 -9019 -10394 -8939
rect -16558 -9024 -16458 -9019
rect -16164 -9024 -16064 -9019
rect -15766 -9024 -15666 -9019
rect -10497 -9024 -10394 -9019
rect -14542 -9375 -14442 -9370
rect -14542 -9455 -14532 -9375
rect -14452 -9455 -10606 -9375
rect -14542 -9460 -14442 -9455
rect -16355 -9573 -16255 -9568
rect -15956 -9573 -15856 -9568
rect -15546 -9573 -15446 -9568
rect -10430 -9573 -10327 -9568
rect -16355 -9653 -16345 -9573
rect -16265 -9653 -15946 -9573
rect -15866 -9653 -15536 -9573
rect -15456 -9653 -10420 -9573
rect -10337 -9653 -10327 -9573
rect -16355 -9658 -16255 -9653
rect -15956 -9658 -15856 -9653
rect -15546 -9658 -15446 -9653
rect -10430 -9658 -10327 -9653
use auto_sampling  auto_sampling_0
timestamp 1730797079
transform 1 0 -1322 0 1 5806
box -884 -4024 11778 -1704
use cdac_ctrl  cdac_ctrl_0
timestamp 1730797079
transform 1 0 -9316 0 1 -9531
box -1485 -724 19472 718
use cyclic_flag  cyclic_flag_0
timestamp 1730797164
transform 1 0 -987 0 1 -2850
box -169 910 11075 2602
use out_latch  out_latch_0
timestamp 1730797079
transform 1 0 -434 0 1 -5175
box -182 -873 10574 956
<< end >>
