magic
tech sky130A
magscale 1 2
timestamp 1731350402
<< metal1 >>
rect -4084864 -1944623 -4084854 -1942623
rect -4082854 -1944615 -3985360 -1942623
rect -4082854 -1944623 -4082844 -1944615
rect -3985370 -1944623 -3985360 -1944615
rect -3983360 -1944623 -3983350 -1942623
rect -4084854 -2087258 -4082854 -1944623
rect -4076864 -1952426 -4076854 -1950426
rect -4074854 -1950427 -4036211 -1950426
rect -4074854 -1952426 -4038014 -1950427
rect -4037885 -1952426 -4036211 -1950427
rect -4032109 -1952426 -4030396 -1950426
rect -4030267 -1952426 -3993360 -1950426
rect -3991360 -1952426 -3991350 -1950426
rect -4080871 -2039463 -4080861 -2039277
rect -4078853 -2039463 -4078843 -2039277
rect -4084864 -2087356 -4084854 -2087258
rect -4082854 -2087259 -4077909 -2087258
rect -4082854 -2087356 -4077910 -2087259
rect -4084854 -2087659 -4082854 -2087356
rect -4078008 -2087357 -4077910 -2087356
rect -4077920 -2087358 -4077910 -2087357
rect -4077811 -2087358 -4077801 -2087259
rect -4081936 -2087559 -4081930 -2087459
rect -4081830 -2087559 -4077908 -2087459
rect -4077808 -2087559 -4077802 -2087459
rect -4084864 -2087758 -4084854 -2087659
rect -4082854 -2087758 -4077907 -2087659
rect -4077808 -2087758 -4077798 -2087659
rect -4084854 -2088059 -4082854 -2087758
rect -4081938 -2087959 -4081928 -2087859
rect -4081828 -2087959 -4077906 -2087859
rect -4077806 -2087959 -4077796 -2087859
rect -4084864 -2088159 -4084854 -2088059
rect -4082854 -2088159 -4077905 -2088059
rect -4077805 -2088159 -4077795 -2088059
rect -4084854 -2111976 -4082854 -2088159
rect -4081937 -2088359 -4081927 -2088259
rect -4081827 -2088359 -4077905 -2088259
rect -4077805 -2088359 -4077795 -2088259
rect -4076854 -2103911 -4074854 -1952426
rect -4038014 -1956629 -4037885 -1952426
rect -4037066 -1953467 -4037056 -1953363
rect -4036952 -1953467 -4036942 -1953363
rect -4038024 -1956758 -4038014 -1956629
rect -4037885 -1956758 -4037875 -1956629
rect -4037056 -1956701 -4036952 -1953467
rect -4031380 -1953473 -4031370 -1953369
rect -4031266 -1953473 -4031256 -1953369
rect -4031370 -1956697 -4031266 -1953473
rect -4030396 -1956630 -4030267 -1952426
rect -3997370 -1956224 -3997360 -1954224
rect -3995360 -1956224 -3995350 -1954224
rect -4037066 -1956805 -4037056 -1956701
rect -4036952 -1956805 -4036942 -1956701
rect -4031380 -1956801 -4031370 -1956697
rect -4031266 -1956801 -4031256 -1956697
rect -4030406 -1956759 -4030396 -1956630
rect -4030267 -1956759 -4030257 -1956630
rect -4068864 -1960237 -4068854 -1958237
rect -4066854 -1960237 -4036211 -1958237
rect -4032109 -1960237 -4001360 -1958237
rect -3999360 -1960237 -3999350 -1958237
rect -4068854 -1971240 -4066854 -1960237
rect -4037066 -1963360 -4037056 -1963256
rect -4036952 -1963360 -4036942 -1963256
rect -4031380 -1963366 -4031370 -1963262
rect -4031266 -1963366 -4031256 -1963262
rect -4001360 -1971240 -3999360 -1960237
rect -4068864 -1971424 -4068854 -1971240
rect -4066854 -1971424 -4066844 -1971240
rect -4001370 -1971424 -4001360 -1971240
rect -3999360 -1971424 -3999350 -1971240
rect -4068854 -2004048 -4066854 -1971424
rect -4068864 -2004232 -4068854 -2004048
rect -4066854 -2004232 -4066844 -2004048
rect -4068854 -2004834 -4066854 -2004232
rect -4068864 -2005018 -4068854 -2004834
rect -4066854 -2005018 -4066844 -2004834
rect -4068854 -2037641 -4066854 -2005018
rect -4068864 -2037826 -4068854 -2037641
rect -4066854 -2037826 -4066844 -2037641
rect -4001360 -2037642 -3999360 -1971424
rect -4001370 -2037826 -4001360 -2037642
rect -3999363 -2037826 -3999353 -2037642
rect -4074063 -2039463 -4074053 -2039277
rect -4073867 -2039278 -4070460 -2039277
rect -4073867 -2039462 -4070554 -2039278
rect -4070370 -2039462 -4070360 -2039278
rect -4073867 -2039463 -4070460 -2039462
rect -4073889 -2087359 -4073879 -2087259
rect -4073779 -2087359 -4070551 -2087259
rect -4070451 -2087359 -4070441 -2087259
rect -4073886 -2087559 -4073880 -2087459
rect -4073780 -2087559 -4070552 -2087459
rect -4070452 -2087559 -4070442 -2087459
rect -4073888 -2087759 -4073878 -2087659
rect -4073778 -2087759 -4070557 -2087659
rect -4070457 -2087759 -4070447 -2087659
rect -4073889 -2087959 -4073879 -2087859
rect -4073779 -2087959 -4070548 -2087859
rect -4070448 -2087959 -4070438 -2087859
rect -4073891 -2088159 -4073881 -2088059
rect -4073781 -2088159 -4070546 -2088059
rect -4070446 -2088159 -4070436 -2088059
rect -4073889 -2088359 -4073879 -2088259
rect -4073779 -2088359 -4070544 -2088259
rect -4070444 -2088359 -4070434 -2088259
rect -4068854 -2094421 -4066854 -2037826
rect -4064664 -2038968 -4064654 -2038784
rect -4064470 -2038968 -4064460 -2038784
rect -4064654 -2039151 -4064470 -2038968
rect -4065347 -2086259 -4065295 -2048733
rect -4065357 -2086359 -4065347 -2086259
rect -4065295 -2086359 -4065285 -2086259
rect -4065347 -2086369 -4065295 -2086359
rect -4065205 -2086459 -4065153 -2048645
rect -4065214 -2086559 -4065205 -2086459
rect -4065153 -2086559 -4065143 -2086459
rect -4065205 -2086568 -4065153 -2086559
rect -4064654 -2086659 -4064471 -2039151
rect -4064665 -2086760 -4064655 -2086659
rect -4064470 -2086760 -4064460 -2086659
rect -4064654 -2086763 -4064471 -2086760
rect -4001360 -2094421 -3999360 -2037826
rect -3993360 -2039278 -3991360 -1952426
rect -3997791 -2039462 -3997781 -2039278
rect -3997597 -2039462 -3993360 -2039278
rect -3991360 -2039462 -3991350 -2039278
rect -4068864 -2096421 -4068854 -2094421
rect -4066854 -2096421 -4045578 -2094421
rect -4043578 -2096421 -4032760 -2094421
rect -4032359 -2096421 -4032222 -2094421
rect -4031821 -2096421 -4024807 -2094421
rect -4022807 -2096421 -4001360 -2094421
rect -3999360 -2096421 -3999350 -2094421
rect -3993360 -2103837 -3991360 -2039462
rect -4076864 -2105911 -4076854 -2103911
rect -4074854 -2103913 -4074844 -2103911
rect -3993370 -2103913 -3993360 -2103837
rect -4074854 -2105911 -4045578 -2103913
rect -4074494 -2105913 -4045578 -2105911
rect -4043578 -2105913 -4032760 -2103913
rect -4032359 -2105913 -4032222 -2103913
rect -4031821 -2105913 -4024754 -2103913
rect -4022754 -2105837 -3993360 -2103913
rect -3991360 -2105837 -3991350 -2103837
rect -4022754 -2105913 -3991360 -2105837
rect -3993360 -2105914 -3991360 -2105913
rect -3985360 -2111758 -3983360 -1944623
rect -3985370 -2111976 -3985360 -2111758
rect -4084864 -2113976 -4084854 -2111976
rect -4082854 -2113976 -4045578 -2111976
rect -4043578 -2113976 -4032760 -2111976
rect -4032359 -2113976 -4032222 -2111976
rect -4031821 -2113976 -4024754 -2111976
rect -4022754 -2113758 -3985360 -2111976
rect -3983360 -2113758 -3983350 -2111758
rect -4022754 -2113975 -3983360 -2113758
rect -4022754 -2113976 -3985379 -2113975
<< via1 >>
rect -4084854 -1944623 -4082854 -1942623
rect -3985360 -1944623 -3983360 -1942623
rect -4076854 -1952426 -4074854 -1950426
rect -4038014 -1952426 -4037885 -1950427
rect -4030396 -1952426 -4030267 -1950426
rect -3993360 -1952426 -3991360 -1950426
rect -4080861 -2039463 -4078853 -2039277
rect -4084854 -2087356 -4082854 -2087258
rect -4077910 -2087358 -4077811 -2087259
rect -4081930 -2087559 -4081830 -2087459
rect -4077908 -2087559 -4077808 -2087459
rect -4084854 -2087758 -4082854 -2087659
rect -4077907 -2087758 -4077808 -2087659
rect -4081928 -2087959 -4081828 -2087859
rect -4077906 -2087959 -4077806 -2087859
rect -4084854 -2088159 -4082854 -2088059
rect -4077905 -2088159 -4077805 -2088059
rect -4081927 -2088359 -4081827 -2088259
rect -4077905 -2088359 -4077805 -2088259
rect -4037056 -1953467 -4036952 -1953363
rect -4038014 -1956758 -4037885 -1956629
rect -4031370 -1953473 -4031266 -1953369
rect -3997360 -1956224 -3995360 -1954224
rect -4037056 -1956805 -4036952 -1956701
rect -4031370 -1956801 -4031266 -1956697
rect -4030396 -1956759 -4030267 -1956630
rect -4068854 -1960237 -4066854 -1958237
rect -4001360 -1960237 -3999360 -1958237
rect -4037056 -1963360 -4036952 -1963256
rect -4031370 -1963366 -4031266 -1963262
rect -4068854 -1971424 -4066854 -1971240
rect -4001360 -1971424 -3999360 -1971240
rect -4068854 -2004232 -4066854 -2004048
rect -4068854 -2005018 -4066854 -2004834
rect -4068854 -2037826 -4066854 -2037641
rect -4001360 -2037826 -3999363 -2037642
rect -4074053 -2039463 -4073867 -2039277
rect -4070554 -2039462 -4070370 -2039278
rect -4073879 -2087359 -4073779 -2087259
rect -4070551 -2087359 -4070451 -2087259
rect -4073880 -2087559 -4073780 -2087459
rect -4070552 -2087559 -4070452 -2087459
rect -4073878 -2087759 -4073778 -2087659
rect -4070557 -2087759 -4070457 -2087659
rect -4073879 -2087959 -4073779 -2087859
rect -4070548 -2087959 -4070448 -2087859
rect -4073881 -2088159 -4073781 -2088059
rect -4070546 -2088159 -4070446 -2088059
rect -4073879 -2088359 -4073779 -2088259
rect -4070544 -2088359 -4070444 -2088259
rect -4064654 -2038968 -4064470 -2038784
rect -4065347 -2086359 -4065295 -2086259
rect -4065205 -2086559 -4065153 -2086459
rect -4064655 -2086760 -4064470 -2086659
rect -3997781 -2039462 -3997597 -2039278
rect -3993360 -2039462 -3991360 -2039278
rect -4068854 -2096421 -4066854 -2094421
rect -4045578 -2096421 -4043578 -2094421
rect -4024807 -2096421 -4022807 -2094421
rect -4001360 -2096421 -3999360 -2094421
rect -4076854 -2105911 -4074854 -2103911
rect -4045578 -2105913 -4043578 -2103913
rect -4024754 -2105913 -4022754 -2103913
rect -3993360 -2105837 -3991360 -2103837
rect -4084854 -2113976 -4082854 -2111976
rect -4045578 -2113976 -4043578 -2111976
rect -4024754 -2113976 -4022754 -2111976
rect -3985360 -2113758 -3983360 -2111758
<< metal2 >>
rect -4034774 -1936461 -4034574 -1936460
rect -4088854 -1938117 -4086850 -1938107
rect -4086850 -1940119 -4036211 -1938117
rect -4086850 -1940121 -4080854 -1940119
rect -4088854 -1940131 -4086850 -1940121
rect -4088854 -2087449 -4086854 -1940131
rect -4084854 -1942623 -4082854 -1942613
rect -4084854 -1944633 -4082854 -1944623
rect -4080854 -1946414 -4078854 -1946404
rect -4037056 -1946414 -4036952 -1946404
rect -4078854 -1948414 -4037056 -1946414
rect -4036952 -1948414 -4036211 -1946414
rect -4080854 -2039267 -4078854 -1948414
rect -4076854 -1950426 -4074854 -1950416
rect -4076854 -1952436 -4074854 -1952426
rect -4038014 -1950427 -4037885 -1950417
rect -4038014 -1952436 -4037885 -1952426
rect -4037056 -1953363 -4036952 -1948414
rect -4037056 -1953477 -4036952 -1953467
rect -4072854 -1954224 -4070854 -1954214
rect -4070854 -1956224 -4036211 -1954224
rect -4072854 -1971635 -4070854 -1956224
rect -4038014 -1956629 -4037885 -1956619
rect -4068854 -1958237 -4066854 -1958227
rect -4068854 -1960247 -4066854 -1960237
rect -4038014 -1969734 -4037885 -1956758
rect -4037056 -1956701 -4036952 -1956691
rect -4037056 -1963256 -4036952 -1956805
rect -4037056 -1963370 -4036952 -1963360
rect -4034774 -1963311 -4034374 -1936461
rect -4034774 -1963447 -4034574 -1963311
rect -4033948 -1963313 -4033548 -1936460
rect -3981362 -1938117 -3979360 -1938107
rect -4032109 -1940119 -3981362 -1938117
rect -3981362 -1940129 -3979360 -1940119
rect -3985360 -1942623 -3983360 -1942613
rect -3985360 -1944633 -3983360 -1944623
rect -4031370 -1946414 -4031266 -1946404
rect -3989360 -1946414 -3987360 -1946406
rect -4032109 -1948414 -4031370 -1946414
rect -4031266 -1946416 -3987360 -1946414
rect -4031266 -1948414 -3989360 -1946416
rect -4031370 -1953369 -4031266 -1948414
rect -4030396 -1950426 -4030267 -1950416
rect -4030396 -1952436 -4030267 -1952426
rect -3993360 -1950426 -3991360 -1950416
rect -3993360 -1952436 -3991360 -1952426
rect -4031370 -1953483 -4031266 -1953473
rect -3997360 -1954224 -3995360 -1954214
rect -4032109 -1956224 -3997360 -1954224
rect -4030396 -1956630 -4030267 -1956620
rect -4033748 -1963447 -4033548 -1963313
rect -4031370 -1956697 -4031266 -1956687
rect -4031370 -1963262 -4031266 -1956801
rect -4031370 -1963376 -4031266 -1963366
rect -4030396 -1969734 -4030267 -1956759
rect -4001360 -1958237 -3999360 -1958227
rect -4001360 -1960247 -3999360 -1960237
rect -4070124 -1970838 -4069524 -1970828
rect -3998674 -1970836 -3998076 -1970826
rect -4069524 -1971022 -4065614 -1970838
rect -4070124 -1971032 -4069524 -1971022
rect -4065798 -1971028 -4065614 -1971022
rect -4002879 -1971020 -3998674 -1970836
rect -4002879 -1971028 -4002695 -1971020
rect -4065798 -1971212 -4064210 -1971028
rect -4004150 -1971212 -4002695 -1971028
rect -3998674 -1971031 -3998076 -1971021
rect -4068854 -1971240 -4066854 -1971230
rect -4001360 -1971240 -3999360 -1971230
rect -4066854 -1971424 -4064050 -1971240
rect -4004075 -1971424 -4001360 -1971240
rect -4068854 -1971434 -4066854 -1971424
rect -4001360 -1971434 -3999360 -1971424
rect -4065797 -1971635 -4064278 -1971452
rect -4070854 -1971636 -4064278 -1971635
rect -4004077 -1971635 -4002713 -1971452
rect -3997360 -1971625 -3995360 -1956224
rect -3997360 -1971635 -3995357 -1971625
rect -4004077 -1971636 -3997360 -1971635
rect -4070854 -1971819 -4065613 -1971636
rect -4002897 -1971819 -3997360 -1971636
rect -4072854 -2003655 -4070854 -1971819
rect -3997360 -1971829 -3995357 -1971819
rect -3997360 -2003642 -3995360 -1971829
rect -4070854 -2003836 -4065611 -2003656
rect -4002889 -2003826 -3997360 -2003642
rect -3995360 -2003826 -3995359 -2003642
rect -4002889 -2003836 -4002705 -2003826
rect -4070854 -2003840 -4064227 -2003836
rect -4072854 -2005222 -4070854 -2003840
rect -4065795 -2004020 -4064227 -2003840
rect -4004217 -2004020 -4002705 -2003836
rect -4068854 -2004048 -4066854 -2004038
rect -4001360 -2004048 -3999360 -2004038
rect -4068858 -2004232 -4068854 -2004048
rect -4066854 -2004232 -4064083 -2004048
rect -4004262 -2004232 -4001360 -2004048
rect -3999360 -2004232 -3999357 -2004048
rect -4068854 -2004242 -4066854 -2004232
rect -4001360 -2004242 -3999360 -2004232
rect -4070124 -2004441 -4069524 -2004431
rect -4064550 -2004441 -4064366 -2004276
rect -4069524 -2004625 -4064366 -2004441
rect -4070124 -2004635 -4069524 -2004625
rect -4064550 -2004806 -4064366 -2004625
rect -4003955 -2004438 -4003771 -2004273
rect -3998675 -2004438 -3998074 -2004428
rect -4003955 -2004622 -3998675 -2004438
rect -4003955 -2004806 -4003771 -2004622
rect -3998675 -2004632 -3998074 -2004622
rect -4068854 -2004834 -4066854 -2004824
rect -4001360 -2004834 -3999360 -2004824
rect -4068855 -2005018 -4068854 -2004834
rect -4066854 -2005018 -4064108 -2004834
rect -4004257 -2005018 -4001360 -2004834
rect -3999360 -2005018 -3999357 -2004834
rect -4068854 -2005028 -4066854 -2005018
rect -4001360 -2005028 -3999360 -2005018
rect -4072856 -2005232 -4070854 -2005222
rect -4065797 -2005230 -4064283 -2005046
rect -4004192 -2005230 -4002705 -2005046
rect -3997360 -2005230 -3995360 -2003826
rect -4065797 -2005232 -4065613 -2005230
rect -4070854 -2005416 -4065613 -2005232
rect -4002889 -2005414 -3997360 -2005230
rect -4072856 -2005426 -4070854 -2005416
rect -4072854 -2037243 -4070854 -2005426
rect -3997360 -2037232 -3995360 -2005414
rect -3997361 -2037242 -3995360 -2037232
rect -4070854 -2037427 -4065611 -2037243
rect -4080861 -2039277 -4078853 -2039267
rect -4074053 -2039277 -4073867 -2039267
rect -4078853 -2039463 -4074053 -2039277
rect -4080861 -2039473 -4078853 -2039463
rect -4074053 -2039473 -4073867 -2039463
rect -4084854 -2087258 -4082854 -2087248
rect -4084854 -2087366 -4082854 -2087356
rect -4088858 -2087459 -4086854 -2087449
rect -4081930 -2087459 -4081830 -2087449
rect -4086854 -2087559 -4081930 -2087459
rect -4088858 -2087569 -4086854 -2087559
rect -4081930 -2087569 -4081830 -2087559
rect -4088854 -2087859 -4086854 -2087569
rect -4084854 -2087659 -4082854 -2087649
rect -4084854 -2087768 -4082854 -2087758
rect -4081928 -2087859 -4081828 -2087849
rect -4086854 -2087959 -4081928 -2087859
rect -4088854 -2088259 -4086854 -2087959
rect -4081928 -2087969 -4081828 -2087959
rect -4084854 -2088059 -4082854 -2088049
rect -4084854 -2088169 -4082854 -2088159
rect -4081927 -2088259 -4081827 -2088249
rect -4086854 -2088359 -4081927 -2088259
rect -4088854 -2116206 -4086854 -2088359
rect -4081927 -2088369 -4081827 -2088359
rect -4080854 -2107845 -4078854 -2039473
rect -4077910 -2087259 -4077811 -2087249
rect -4073879 -2087259 -4073779 -2087249
rect -4077811 -2087358 -4073879 -2087259
rect -4077910 -2087368 -4077811 -2087358
rect -4073978 -2087359 -4073879 -2087358
rect -4073879 -2087369 -4073779 -2087359
rect -4077908 -2087459 -4077808 -2087449
rect -4073880 -2087459 -4073780 -2087449
rect -4077808 -2087559 -4073880 -2087459
rect -4077908 -2087569 -4077808 -2087559
rect -4073880 -2087569 -4073780 -2087559
rect -4077907 -2087659 -4077808 -2087649
rect -4073878 -2087659 -4073778 -2087649
rect -4077808 -2087758 -4073878 -2087659
rect -4077907 -2087768 -4077808 -2087758
rect -4073977 -2087759 -4073878 -2087758
rect -4073878 -2087769 -4073778 -2087759
rect -4077906 -2087859 -4077806 -2087849
rect -4073879 -2087859 -4073779 -2087849
rect -4077806 -2087959 -4073879 -2087859
rect -4077906 -2087969 -4077806 -2087959
rect -4073879 -2087969 -4073779 -2087959
rect -4077905 -2088059 -4077805 -2088049
rect -4073881 -2088059 -4073781 -2088049
rect -4077805 -2088159 -4073881 -2088059
rect -4077905 -2088169 -4077805 -2088159
rect -4073881 -2088169 -4073781 -2088159
rect -4077905 -2088259 -4077805 -2088249
rect -4073879 -2088259 -4073779 -2088249
rect -4077805 -2088359 -4073879 -2088259
rect -4077905 -2088369 -4077805 -2088359
rect -4073879 -2088369 -4073779 -2088359
rect -4072854 -2099361 -4070854 -2037427
rect -4065795 -2037430 -4065611 -2037427
rect -4002891 -2037426 -3997361 -2037242
rect -4002891 -2037430 -4002707 -2037426
rect -4065795 -2037614 -4064586 -2037430
rect -4004155 -2037614 -4002707 -2037430
rect -3997361 -2037436 -3995360 -2037426
rect -4068854 -2037641 -4066854 -2037631
rect -4001360 -2037642 -3999363 -2037632
rect -4066854 -2037826 -4064305 -2037642
rect -4004148 -2037826 -4001360 -2037642
rect -4068854 -2037836 -4066854 -2037826
rect -4001360 -2037836 -3999363 -2037826
rect -4065790 -2038038 -4064584 -2037854
rect -4004157 -2038038 -4002705 -2037854
rect -4070123 -2038052 -4069524 -2038042
rect -4065790 -2038052 -4065606 -2038038
rect -4069524 -2038236 -4065606 -2038052
rect -4002889 -2038071 -4002705 -2038038
rect -3998675 -2038071 -3998074 -2038061
rect -4070123 -2038246 -4069524 -2038236
rect -4002889 -2038255 -3998675 -2038071
rect -3998675 -2038265 -3998074 -2038255
rect -4064654 -2038784 -4064470 -2038774
rect -4064470 -2038968 -4063944 -2038784
rect -4064654 -2038978 -4064470 -2038968
rect -4070554 -2039278 -4070370 -2039268
rect -3997781 -2039278 -3997597 -2039268
rect -4070370 -2039462 -4063041 -2039278
rect -4003288 -2039462 -3997781 -2039278
rect -4070554 -2039472 -4070370 -2039462
rect -3997781 -2039472 -3997597 -2039462
rect -4027621 -2044907 -4027437 -2044897
rect -4040961 -2044978 -4040777 -2044968
rect -4027621 -2045101 -4027437 -2045091
rect -4040961 -2045172 -4040777 -2045162
rect -4027252 -2045407 -4027068 -2045397
rect -4041324 -2045480 -4041140 -2045470
rect -4027252 -2045601 -4027068 -2045591
rect -4041324 -2045674 -4041140 -2045664
rect -4026884 -2045907 -4026700 -2045897
rect -4041690 -2045976 -4041506 -2045966
rect -4026884 -2046101 -4026700 -2046091
rect -4041690 -2046170 -4041506 -2046160
rect -4026516 -2046407 -4026332 -2046397
rect -4042057 -2046478 -4041873 -2046468
rect -4026516 -2046601 -4026332 -2046591
rect -4042057 -2046672 -4041873 -2046662
rect -4026148 -2046907 -4025964 -2046897
rect -4042424 -2046978 -4042240 -2046968
rect -4026148 -2047101 -4025964 -2047091
rect -4042424 -2047172 -4042240 -2047162
rect -4034752 -2053558 -4034652 -2053548
rect -4034752 -2053668 -4034652 -2053658
rect -4033669 -2053603 -4033569 -2053593
rect -4033669 -2053713 -4033569 -2053703
rect -4033669 -2054177 -4033569 -2054167
rect -4033669 -2054287 -4033569 -2054277
rect -4034752 -2054377 -4034652 -2054367
rect -4034752 -2054487 -4034652 -2054477
rect -4027858 -2054589 -4027790 -2054579
rect -4027858 -2054672 -4027790 -2054662
rect -4028015 -2054788 -4027947 -2054778
rect -4028015 -2054871 -4027947 -2054861
rect -4028171 -2054987 -4028103 -2054977
rect -4028171 -2055070 -4028103 -2055060
rect -4028326 -2055188 -4028258 -2055178
rect -4028326 -2055271 -4028258 -2055261
rect -4028482 -2055388 -4028414 -2055378
rect -4028482 -2055471 -4028414 -2055461
rect -4028639 -2055590 -4028571 -2055580
rect -4028639 -2055673 -4028571 -2055663
rect -4028794 -2055790 -4028726 -2055780
rect -4028794 -2055873 -4028726 -2055863
rect -4028950 -2055988 -4028882 -2055978
rect -4028950 -2056071 -4028882 -2056061
rect -4029106 -2056190 -4029038 -2056180
rect -4029106 -2056273 -4029038 -2056263
rect -4029262 -2056390 -4029194 -2056380
rect -4029262 -2056473 -4029194 -2056463
rect -4040535 -2056589 -4040461 -2056579
rect -4040535 -2056677 -4040461 -2056667
rect -4040378 -2056787 -4040304 -2056777
rect -4040378 -2056875 -4040304 -2056865
rect -4040223 -2056987 -4040149 -2056977
rect -4040223 -2057075 -4040149 -2057065
rect -4040067 -2057188 -4039993 -2057178
rect -4040067 -2057276 -4039993 -2057266
rect -4039911 -2057388 -4039837 -2057378
rect -4039911 -2057476 -4039837 -2057466
rect -4039755 -2057587 -4039681 -2057577
rect -4039755 -2057675 -4039681 -2057665
rect -4039599 -2057787 -4039525 -2057777
rect -4039599 -2057875 -4039525 -2057865
rect -4039443 -2057987 -4039369 -2057977
rect -4039443 -2058075 -4039369 -2058065
rect -4039288 -2058188 -4039214 -2058178
rect -4039288 -2058276 -4039214 -2058266
rect -4039145 -2058387 -4038891 -2058377
rect -4039145 -2058465 -4039131 -2058387
rect -4039057 -2058465 -4038891 -2058387
rect -4039145 -2058477 -4038891 -2058465
rect -4040916 -2058577 -4040816 -2058567
rect -4040816 -2058677 -4039804 -2058577
rect -4040916 -2058687 -4040816 -2058677
rect -4041282 -2058777 -4041182 -2058767
rect -4042722 -2058877 -4041282 -2058777
rect -4041282 -2058887 -4041182 -2058877
rect -4041651 -2058977 -4041551 -2058967
rect -4042763 -2059077 -4041651 -2058977
rect -4041651 -2059087 -4041551 -2059077
rect -4042013 -2059177 -4041913 -2059167
rect -4042800 -2059277 -4042013 -2059177
rect -4042013 -2059287 -4041913 -2059277
rect -4042379 -2059377 -4042279 -2059367
rect -4042855 -2059477 -4042379 -2059377
rect -4042379 -2059487 -4042279 -2059477
rect -4026108 -2059577 -4026008 -2059567
rect -4027962 -2059677 -4026108 -2059577
rect -4026108 -2059687 -4026008 -2059677
rect -4026474 -2059777 -4026374 -2059767
rect -4027965 -2059877 -4026474 -2059777
rect -4026474 -2059887 -4026374 -2059877
rect -4026844 -2059977 -4026744 -2059967
rect -4027942 -2060077 -4026844 -2059977
rect -4026844 -2060087 -4026744 -2060077
rect -4027210 -2060177 -4027110 -2060167
rect -4027930 -2060277 -4027210 -2060177
rect -4027210 -2060287 -4027110 -2060277
rect -4027578 -2060377 -4027478 -2060367
rect -4027889 -2060477 -4027578 -2060377
rect -4027578 -2060487 -4027478 -2060477
rect -4038594 -2084022 -4038194 -2084012
rect -4038594 -2084153 -4038194 -2084143
rect -4034308 -2084153 -4034188 -2084013
rect -4038046 -2084258 -4037646 -2084248
rect -4038046 -2084369 -4037646 -2084359
rect -4037508 -2084458 -4037108 -2084448
rect -4037508 -2084569 -4037108 -2084559
rect -4036979 -2084658 -4036579 -2084648
rect -4036979 -2084769 -4036579 -2084759
rect -4036449 -2084858 -4036049 -2084848
rect -4036449 -2084969 -4036049 -2084959
rect -4035929 -2085058 -4035529 -2085048
rect -4035929 -2085169 -4035529 -2085159
rect -4035396 -2085259 -4034996 -2085249
rect -4035396 -2085370 -4034996 -2085360
rect -4034873 -2085458 -4034473 -2085448
rect -4034873 -2085569 -4034473 -2085559
rect -4034352 -2085658 -4033952 -2085648
rect -4034352 -2085769 -4033952 -2085759
rect -4033828 -2085858 -4033428 -2085848
rect -4033828 -2085969 -4033428 -2085959
rect -4033291 -2086058 -4032891 -2086048
rect -4033291 -2086169 -4032891 -2086159
rect -4065347 -2086259 -4065295 -2086249
rect -4065357 -2086359 -4065347 -2086259
rect -4065295 -2086359 -4032806 -2086259
rect -4031722 -2086359 -4025410 -2086259
rect -4065347 -2086369 -4065295 -2086359
rect -4065205 -2086459 -4065153 -2086449
rect -4065214 -2086559 -4065205 -2086459
rect -4065153 -2086559 -4032806 -2086459
rect -4031722 -2086559 -4025454 -2086459
rect -4065205 -2086568 -4065153 -2086559
rect -4064655 -2086659 -4064470 -2086649
rect -4032359 -2086659 -4032287 -2086649
rect -4031686 -2086659 -4031286 -2086649
rect -4064666 -2086759 -4064655 -2086659
rect -4064470 -2086759 -4032760 -2086659
rect -4032359 -2086759 -4032222 -2086659
rect -4031821 -2086759 -4031686 -2086659
rect -4064655 -2086770 -4064470 -2086760
rect -4032359 -2086769 -4032287 -2086759
rect -4031286 -2086759 -4025475 -2086659
rect -4031686 -2086770 -4031286 -2086760
rect -4031155 -2087059 -4030754 -2087049
rect -4031155 -2087169 -4030754 -2087159
rect -4070551 -2087259 -4070451 -2087249
rect -4070451 -2087359 -4043061 -2087259
rect -4070551 -2087369 -4070451 -2087359
rect -4070552 -2087459 -4070452 -2087449
rect -4070452 -2087559 -4043096 -2087459
rect -4070552 -2087569 -4070452 -2087559
rect -4070557 -2087659 -4070457 -2087649
rect -4070457 -2087759 -4043012 -2087659
rect -4070557 -2087769 -4070457 -2087759
rect -4070548 -2087859 -4070448 -2087849
rect -4070448 -2087959 -4043076 -2087859
rect -4070548 -2087969 -4070448 -2087959
rect -4070546 -2088059 -4070446 -2088049
rect -4070446 -2088159 -4043014 -2088059
rect -4070546 -2088169 -4070446 -2088159
rect -4070544 -2088259 -4070444 -2088249
rect -4070444 -2088359 -4043288 -2088259
rect -4070544 -2088369 -4070444 -2088359
rect -4068854 -2094421 -4066854 -2094411
rect -4068854 -2096431 -4066854 -2096421
rect -4045578 -2094421 -4043578 -2094411
rect -4045578 -2096431 -4043578 -2096421
rect -4024807 -2094421 -4022807 -2094411
rect -4024807 -2096431 -4022807 -2096421
rect -4001360 -2094421 -3999360 -2094411
rect -4001360 -2096431 -3999360 -2096421
rect -4045578 -2099361 -4043578 -2099351
rect -4024754 -2099361 -4022754 -2099351
rect -3997360 -2099361 -3995360 -2037436
rect -3993360 -2039278 -3991360 -2039268
rect -3993360 -2039472 -3991360 -2039462
rect -4070854 -2101361 -4045578 -2099361
rect -4043578 -2101361 -4032760 -2099361
rect -4032359 -2101361 -4032222 -2099361
rect -4031821 -2101361 -4024754 -2099361
rect -4022754 -2101361 -3997360 -2099361
rect -4072854 -2101371 -4070854 -2101361
rect -4045578 -2101371 -4043578 -2101361
rect -4024754 -2101371 -4022754 -2101361
rect -3997360 -2101371 -3995360 -2101361
rect -3993360 -2103837 -3991360 -2103827
rect -4076854 -2103911 -4074854 -2103901
rect -4076854 -2105921 -4074854 -2105911
rect -4045578 -2103913 -4043578 -2103903
rect -4045578 -2105923 -4043578 -2105913
rect -4024754 -2103913 -4022754 -2103903
rect -3993360 -2105847 -3991360 -2105837
rect -4024754 -2105923 -4022754 -2105913
rect -4045578 -2107845 -4043578 -2107835
rect -4024754 -2107845 -4022754 -2107835
rect -3989360 -2107845 -3987360 -1948416
rect -4080854 -2107846 -4045578 -2107845
rect -4078854 -2109845 -4045578 -2107846
rect -4043578 -2109845 -4032760 -2107845
rect -4032359 -2109845 -4032222 -2107845
rect -4031821 -2109845 -4024754 -2107845
rect -4022754 -2109845 -3989360 -2107845
rect -4080854 -2109856 -4078854 -2109846
rect -4045578 -2109855 -4043578 -2109845
rect -4024754 -2109855 -4022754 -2109845
rect -3989360 -2109855 -3987360 -2109845
rect -3985360 -2111758 -3983360 -2111748
rect -4084854 -2111976 -4082854 -2111966
rect -4084854 -2113986 -4082854 -2113976
rect -4045578 -2111976 -4043578 -2111966
rect -4045578 -2113986 -4043578 -2113976
rect -4024754 -2111976 -4022754 -2111966
rect -3985360 -2113768 -3983360 -2113758
rect -4024754 -2113986 -4022754 -2113976
rect -4045578 -2116206 -4043578 -2116196
rect -4024754 -2116206 -4022754 -2116196
rect -3981360 -2116206 -3979360 -1940129
rect -4086854 -2118206 -4045578 -2116206
rect -4043578 -2118206 -4032760 -2116206
rect -4032359 -2118206 -4032222 -2116206
rect -4031821 -2118206 -4024754 -2116206
rect -4022754 -2118206 -3981360 -2116206
rect -4088854 -2118216 -4086854 -2118206
rect -4045578 -2118216 -4043578 -2118206
rect -4024754 -2118216 -4022754 -2118206
rect -3981360 -2118216 -3979360 -2118206
<< via2 >>
rect -4088854 -1940121 -4086850 -1938117
rect -4084854 -1944623 -4082854 -1942623
rect -4080854 -1948414 -4078854 -1946414
rect -4037056 -1948414 -4036952 -1946414
rect -4076854 -1952426 -4074854 -1950426
rect -4038014 -1952426 -4037885 -1950427
rect -4072854 -1956224 -4070854 -1954224
rect -4068854 -1960237 -4066854 -1958237
rect -3981362 -1940119 -3979360 -1938117
rect -3985360 -1944623 -3983360 -1942623
rect -4031370 -1948414 -4031266 -1946414
rect -3989360 -1948416 -3987360 -1946416
rect -4030396 -1952426 -4030267 -1950426
rect -3993360 -1952426 -3991360 -1950426
rect -4001360 -1960237 -3999360 -1958237
rect -4070124 -1971022 -4069524 -1970838
rect -3998674 -1971021 -3998076 -1970836
rect -4068854 -1971424 -4066854 -1971240
rect -4001360 -1971424 -3999360 -1971240
rect -4072854 -1971819 -4070854 -1971635
rect -3997360 -1971819 -3995357 -1971635
rect -4072854 -2003840 -4070854 -2003655
rect -3997360 -2003826 -3995360 -2003642
rect -4068854 -2004232 -4066854 -2004048
rect -4001360 -2004232 -3999360 -2004048
rect -4070124 -2004625 -4069524 -2004441
rect -3998675 -2004622 -3998074 -2004438
rect -4068854 -2005018 -4066854 -2004834
rect -4001360 -2005018 -3999360 -2004834
rect -4072856 -2005416 -4070854 -2005232
rect -3997360 -2005414 -3995360 -2005230
rect -4072854 -2037427 -4070854 -2037243
rect -4080861 -2039463 -4078853 -2039277
rect -4084854 -2087356 -4082854 -2087258
rect -4088858 -2087559 -4086854 -2087459
rect -4084854 -2087758 -4082854 -2087659
rect -4088854 -2087959 -4086854 -2087859
rect -4084854 -2088159 -4082854 -2088059
rect -4088854 -2088359 -4086854 -2088259
rect -3997361 -2037426 -3995360 -2037242
rect -4068854 -2037826 -4066854 -2037641
rect -4001360 -2037826 -3999363 -2037642
rect -4070123 -2038236 -4069524 -2038052
rect -3998675 -2038255 -3998074 -2038071
rect -4040961 -2045162 -4040777 -2044978
rect -4027621 -2045091 -4027437 -2044907
rect -4041324 -2045664 -4041140 -2045480
rect -4027252 -2045591 -4027068 -2045407
rect -4041690 -2046160 -4041506 -2045976
rect -4026884 -2046091 -4026700 -2045907
rect -4042057 -2046662 -4041873 -2046478
rect -4026516 -2046591 -4026332 -2046407
rect -4042424 -2047162 -4042240 -2046978
rect -4026148 -2047091 -4025964 -2046907
rect -4034752 -2053658 -4034652 -2053558
rect -4033669 -2053703 -4033569 -2053603
rect -4033669 -2054277 -4033569 -2054177
rect -4034752 -2054477 -4034652 -2054377
rect -4027858 -2054662 -4027790 -2054589
rect -4028015 -2054861 -4027947 -2054788
rect -4028171 -2055060 -4028103 -2054987
rect -4028326 -2055261 -4028258 -2055188
rect -4028482 -2055461 -4028414 -2055388
rect -4028639 -2055663 -4028571 -2055590
rect -4028794 -2055863 -4028726 -2055790
rect -4028950 -2056061 -4028882 -2055988
rect -4029106 -2056263 -4029038 -2056190
rect -4029262 -2056463 -4029194 -2056390
rect -4040535 -2056667 -4040461 -2056589
rect -4040378 -2056865 -4040304 -2056787
rect -4040223 -2057065 -4040149 -2056987
rect -4040067 -2057266 -4039993 -2057188
rect -4039911 -2057466 -4039837 -2057388
rect -4039755 -2057665 -4039681 -2057587
rect -4039599 -2057865 -4039525 -2057787
rect -4039443 -2058065 -4039369 -2057987
rect -4039288 -2058266 -4039214 -2058188
rect -4039131 -2058465 -4039057 -2058387
rect -4040916 -2058677 -4040816 -2058577
rect -4041282 -2058877 -4041182 -2058777
rect -4041651 -2059077 -4041551 -2058977
rect -4042013 -2059277 -4041913 -2059177
rect -4042379 -2059477 -4042279 -2059377
rect -4026108 -2059677 -4026008 -2059577
rect -4026474 -2059877 -4026374 -2059777
rect -4026844 -2060077 -4026744 -2059977
rect -4027210 -2060277 -4027110 -2060177
rect -4027578 -2060477 -4027478 -2060377
rect -4038594 -2084143 -4038194 -2084022
rect -4038046 -2084359 -4037646 -2084258
rect -4037508 -2084559 -4037108 -2084458
rect -4036979 -2084759 -4036579 -2084658
rect -4036449 -2084959 -4036049 -2084858
rect -4035929 -2085159 -4035529 -2085058
rect -4035396 -2085360 -4034996 -2085259
rect -4034873 -2085559 -4034473 -2085458
rect -4034352 -2085759 -4033952 -2085658
rect -4033828 -2085959 -4033428 -2085858
rect -4033291 -2086159 -4032891 -2086058
rect -4031686 -2086760 -4031286 -2086659
rect -4031155 -2087159 -4030754 -2087059
rect -4068854 -2096421 -4066854 -2094421
rect -4045578 -2096421 -4043578 -2094421
rect -4024807 -2096421 -4022807 -2094421
rect -3993360 -2039462 -3991360 -2039278
rect -4072854 -2101361 -4070854 -2099361
rect -4045578 -2101361 -4043578 -2099361
rect -4024754 -2101361 -4022754 -2099361
rect -3997360 -2101361 -3995360 -2099361
rect -4076854 -2105911 -4074854 -2103911
rect -4045578 -2105913 -4043578 -2103913
rect -4024754 -2105913 -4022754 -2103913
rect -3993360 -2105837 -3991360 -2103837
rect -4080854 -2109846 -4078854 -2107846
rect -4045578 -2109845 -4043578 -2107845
rect -4024754 -2109845 -4022754 -2107845
rect -3989360 -2109845 -3987360 -2107845
rect -4084854 -2113976 -4082854 -2111976
rect -4045578 -2113976 -4043578 -2111976
rect -4024754 -2113976 -4022754 -2111976
rect -3985360 -2113758 -3983360 -2111758
rect -4088854 -2118206 -4086854 -2116206
rect -4045578 -2118206 -4043578 -2116206
rect -4024754 -2118206 -4022754 -2116206
rect -3981360 -2118206 -3979360 -2116206
<< metal3 >>
rect -4088864 -1938117 -4086840 -1938112
rect -4088864 -1940121 -4088854 -1938117
rect -4086850 -1940121 -4086840 -1938117
rect -4088864 -1940126 -4086840 -1940121
rect -3981372 -1938117 -3979350 -1938112
rect -3981372 -1940119 -3981362 -1938117
rect -3979360 -1940119 -3979350 -1938117
rect -3981372 -1940124 -3979350 -1940119
rect -4084864 -1942623 -4082844 -1942618
rect -3985370 -1942623 -3983350 -1942618
rect -4084864 -1944623 -4084854 -1942623
rect -4082854 -1944615 -4036211 -1942623
rect -4032109 -1944615 -3985360 -1942623
rect -4082854 -1944623 -4082844 -1944615
rect -4084864 -1944628 -4082844 -1944623
rect -3985370 -1944623 -3985360 -1944615
rect -3983360 -1944623 -3983350 -1942623
rect -3985370 -1944628 -3983350 -1944623
rect -4084854 -2087253 -4082854 -1944628
rect -4080864 -1946414 -4078844 -1946409
rect -4080864 -1948414 -4080854 -1946414
rect -4078854 -1948414 -4078844 -1946414
rect -4080864 -1948419 -4078844 -1948414
rect -4037066 -1946414 -4036942 -1946409
rect -4037066 -1948414 -4037056 -1946414
rect -4036952 -1948414 -4036942 -1946414
rect -4037066 -1948419 -4036942 -1948414
rect -4031380 -1946414 -4031256 -1946409
rect -4031380 -1948414 -4031370 -1946414
rect -4031266 -1948414 -4031256 -1946414
rect -4031380 -1948419 -4031256 -1948414
rect -3989370 -1946416 -3987350 -1946411
rect -3989370 -1948416 -3989360 -1946416
rect -3987360 -1948416 -3987350 -1946416
rect -3989370 -1948421 -3987350 -1948416
rect -4076864 -1950426 -4074844 -1950421
rect -4038024 -1950426 -4037875 -1950422
rect -4030406 -1950426 -4030257 -1950421
rect -3993370 -1950426 -3991350 -1950421
rect -4076864 -1952426 -4076854 -1950426
rect -4074854 -1950427 -4030396 -1950426
rect -4074854 -1952426 -4038014 -1950427
rect -4037885 -1952426 -4030396 -1950427
rect -4030267 -1952426 -3993360 -1950426
rect -3991360 -1952426 -3991350 -1950426
rect -4076864 -1952431 -4074844 -1952426
rect -4038024 -1952431 -4037875 -1952426
rect -4030406 -1952431 -4030257 -1952426
rect -3993370 -1952431 -3991350 -1952426
rect -4080871 -2039277 -4078843 -2039272
rect -4080871 -2039463 -4080861 -2039277
rect -4078853 -2039463 -4078843 -2039277
rect -4080871 -2039468 -4078843 -2039463
rect -4084864 -2087258 -4082844 -2087253
rect -4084864 -2087356 -4084854 -2087258
rect -4082854 -2087356 -4082844 -2087258
rect -4084864 -2087361 -4082844 -2087356
rect -4088868 -2087459 -4086844 -2087454
rect -4088868 -2087559 -4088858 -2087459
rect -4086854 -2087559 -4086844 -2087459
rect -4088868 -2087564 -4086844 -2087559
rect -4084854 -2087654 -4082854 -2087361
rect -4084864 -2087659 -4082844 -2087654
rect -4084864 -2087758 -4084854 -2087659
rect -4082854 -2087758 -4082844 -2087659
rect -4084864 -2087763 -4082844 -2087758
rect -4088864 -2087859 -4086844 -2087854
rect -4088864 -2087959 -4088854 -2087859
rect -4086854 -2087959 -4086844 -2087859
rect -4088864 -2087964 -4086844 -2087959
rect -4084854 -2088054 -4082854 -2087763
rect -4084864 -2088059 -4082844 -2088054
rect -4084864 -2088159 -4084854 -2088059
rect -4082854 -2088159 -4082844 -2088059
rect -4084864 -2088164 -4082844 -2088159
rect -4088864 -2088259 -4086844 -2088254
rect -4088864 -2088359 -4088854 -2088259
rect -4086854 -2088359 -4086844 -2088259
rect -4088864 -2088364 -4086844 -2088359
rect -4084854 -2111971 -4082854 -2088164
rect -4076854 -2103906 -4074854 -1952431
rect -4072864 -1954224 -4070844 -1954219
rect -4072864 -1956224 -4072854 -1954224
rect -4070854 -1956224 -4070844 -1954224
rect -3997370 -1956224 -3997360 -1954224
rect -3995360 -1956224 -3995350 -1954224
rect -4072864 -1956229 -4070844 -1956224
rect -4070124 -1956854 -4069524 -1956853
rect -4070124 -1957454 -4036211 -1956854
rect -4032109 -1957454 -3998075 -1956854
rect -4070124 -1970833 -4069524 -1957454
rect -4068864 -1958237 -4066844 -1958232
rect -4001370 -1958237 -3999350 -1958232
rect -4068864 -1960237 -4068854 -1958237
rect -4066854 -1960237 -4001360 -1958237
rect -3999360 -1960237 -3999350 -1958237
rect -4068864 -1960242 -4066844 -1960237
rect -4001370 -1960242 -3999350 -1960237
rect -4070134 -1970838 -4069514 -1970833
rect -4070134 -1971022 -4070124 -1970838
rect -4069524 -1971022 -4069514 -1970838
rect -4070134 -1971027 -4069514 -1971022
rect -4072864 -1971635 -4070844 -1971630
rect -4072864 -1971819 -4072854 -1971635
rect -4070854 -1971819 -4070844 -1971635
rect -4072864 -1971824 -4070844 -1971819
rect -4072864 -2003655 -4070844 -2003650
rect -4072864 -2003840 -4072854 -2003655
rect -4070854 -2003840 -4070844 -2003655
rect -4072864 -2003845 -4070844 -2003840
rect -4070124 -2004436 -4069524 -1971027
rect -4068854 -1971235 -4066854 -1960242
rect -4001360 -1971235 -3999360 -1960242
rect -3998675 -1970831 -3998075 -1957454
rect -3998684 -1970836 -3998066 -1970831
rect -3998684 -1971021 -3998674 -1970836
rect -3998076 -1971021 -3998066 -1970836
rect -3998684 -1971026 -3998066 -1971021
rect -4068864 -1971240 -4066844 -1971235
rect -4068864 -1971424 -4068854 -1971240
rect -4066854 -1971424 -4066844 -1971240
rect -4068864 -1971429 -4066844 -1971424
rect -4001370 -1971240 -3999350 -1971235
rect -4001370 -1971424 -4001360 -1971240
rect -3999360 -1971424 -3999350 -1971240
rect -4001370 -1971429 -3999350 -1971424
rect -4068854 -2004043 -4066854 -1971429
rect -4001360 -2004043 -3999360 -1971429
rect -4068864 -2004048 -4066844 -2004043
rect -4068864 -2004232 -4068854 -2004048
rect -4066854 -2004232 -4066844 -2004048
rect -4068864 -2004237 -4066844 -2004232
rect -4001370 -2004048 -3999350 -2004043
rect -4001370 -2004232 -4001360 -2004048
rect -3999360 -2004232 -3999350 -2004048
rect -4001370 -2004237 -3999350 -2004232
rect -4070134 -2004441 -4069514 -2004436
rect -4070134 -2004625 -4070124 -2004441
rect -4069524 -2004625 -4069514 -2004441
rect -4070134 -2004630 -4069514 -2004625
rect -4072866 -2005232 -4070844 -2005227
rect -4072866 -2005416 -4072856 -2005232
rect -4070854 -2005416 -4070844 -2005232
rect -4072866 -2005421 -4070844 -2005416
rect -4072864 -2037243 -4070844 -2037238
rect -4072864 -2037427 -4072854 -2037243
rect -4070854 -2037427 -4070844 -2037243
rect -4072864 -2037432 -4070844 -2037427
rect -4070124 -2038047 -4069524 -2004630
rect -4068854 -2004829 -4066854 -2004237
rect -4001360 -2004829 -3999360 -2004237
rect -3998675 -2004433 -3998075 -1971026
rect -3997370 -1971635 -3995347 -1971630
rect -3997370 -1971819 -3997360 -1971635
rect -3995357 -1971819 -3995347 -1971635
rect -3997370 -1971824 -3995347 -1971819
rect -3997370 -2003642 -3995350 -2003637
rect -3997370 -2003826 -3997360 -2003642
rect -3995360 -2003826 -3995350 -2003642
rect -3997370 -2003831 -3995350 -2003826
rect -3998685 -2004438 -3998064 -2004433
rect -3998685 -2004622 -3998675 -2004438
rect -3998074 -2004622 -3998064 -2004438
rect -3998685 -2004627 -3998064 -2004622
rect -4068864 -2004834 -4066844 -2004829
rect -4068864 -2005018 -4068854 -2004834
rect -4066854 -2005018 -4066844 -2004834
rect -4068864 -2005023 -4066844 -2005018
rect -4001370 -2004834 -3999350 -2004829
rect -4001370 -2005018 -4001360 -2004834
rect -3999360 -2005018 -3999350 -2004834
rect -4001370 -2005023 -3999350 -2005018
rect -4068854 -2037636 -4066854 -2005023
rect -4068864 -2037641 -4066844 -2037636
rect -4001360 -2037637 -3999360 -2005023
rect -4068864 -2037826 -4068854 -2037641
rect -4066854 -2037826 -4066844 -2037641
rect -4068864 -2037831 -4066844 -2037826
rect -4001370 -2037642 -3999353 -2037637
rect -4001370 -2037826 -4001360 -2037642
rect -3999363 -2037826 -3999353 -2037642
rect -4001370 -2037831 -3999353 -2037826
rect -4070133 -2038052 -4069514 -2038047
rect -4070133 -2038236 -4070123 -2038052
rect -4069524 -2038236 -4069514 -2038052
rect -4070133 -2038241 -4069514 -2038236
rect -4070124 -2097504 -4069524 -2038241
rect -4068854 -2094416 -4066854 -2037831
rect -4040971 -2044978 -4040767 -2044973
rect -4040971 -2045162 -4040961 -2044978
rect -4040777 -2045162 -4040767 -2044978
rect -4040971 -2045167 -4040767 -2045162
rect -4041334 -2045480 -4041130 -2045475
rect -4041334 -2045664 -4041324 -2045480
rect -4041140 -2045664 -4041130 -2045480
rect -4041334 -2045669 -4041130 -2045664
rect -4041700 -2045976 -4041496 -2045971
rect -4041700 -2046160 -4041690 -2045976
rect -4041506 -2046160 -4041496 -2045976
rect -4041700 -2046165 -4041496 -2046160
rect -4042067 -2046478 -4041863 -2046473
rect -4042067 -2046662 -4042057 -2046478
rect -4041873 -2046662 -4041863 -2046478
rect -4042067 -2046667 -4041863 -2046662
rect -4042434 -2046978 -4042230 -2046973
rect -4042434 -2047162 -4042424 -2046978
rect -4042240 -2047162 -4042230 -2046978
rect -4042434 -2047167 -4042230 -2047162
rect -4042424 -2059377 -4042240 -2047167
rect -4042057 -2059177 -4041873 -2046667
rect -4041690 -2058977 -4041506 -2046165
rect -4041324 -2058777 -4041140 -2045669
rect -4040961 -2058577 -4040777 -2045167
rect -4040546 -2056589 -4040450 -2039612
rect -4040546 -2056667 -4040535 -2056589
rect -4040461 -2056667 -4040450 -2056589
rect -4040546 -2056675 -4040450 -2056667
rect -4040390 -2056787 -4040294 -2040174
rect -4040390 -2056865 -4040378 -2056787
rect -4040304 -2056865 -4040294 -2056787
rect -4040390 -2056875 -4040294 -2056865
rect -4040234 -2056987 -4040138 -2040668
rect -4040234 -2057065 -4040223 -2056987
rect -4040149 -2057065 -4040138 -2056987
rect -4040234 -2057075 -4040138 -2057065
rect -4040078 -2057188 -4039982 -2041190
rect -4040078 -2057266 -4040067 -2057188
rect -4039993 -2057266 -4039982 -2057188
rect -4040078 -2057275 -4039982 -2057266
rect -4039922 -2057388 -4039826 -2041672
rect -4039922 -2057466 -4039911 -2057388
rect -4039837 -2057466 -4039826 -2057388
rect -4039922 -2057475 -4039826 -2057466
rect -4039766 -2057587 -4039670 -2042191
rect -4039766 -2057665 -4039755 -2057587
rect -4039681 -2057665 -4039670 -2057587
rect -4039766 -2057677 -4039670 -2057665
rect -4039610 -2057787 -4039514 -2042667
rect -4039610 -2057865 -4039599 -2057787
rect -4039525 -2057865 -4039514 -2057787
rect -4039610 -2057875 -4039514 -2057865
rect -4039454 -2057987 -4039358 -2043155
rect -4039454 -2058065 -4039443 -2057987
rect -4039369 -2058065 -4039358 -2057987
rect -4039454 -2058077 -4039358 -2058065
rect -4039298 -2058188 -4039202 -2043668
rect -4039298 -2058266 -4039288 -2058188
rect -4039214 -2058266 -4039202 -2058188
rect -4039298 -2058275 -4039202 -2058266
rect -4039142 -2058387 -4039046 -2044119
rect -4034762 -2053558 -4034642 -2053553
rect -4034762 -2053658 -4034752 -2053558
rect -4034652 -2053658 -4034642 -2053558
rect -4034762 -2053663 -4034642 -2053658
rect -4033679 -2053603 -4033559 -2053598
rect -4034752 -2054372 -4034652 -2053663
rect -4033679 -2053703 -4033669 -2053603
rect -4033569 -2053703 -4033559 -2053603
rect -4033679 -2053708 -4033559 -2053703
rect -4033669 -2054172 -4033569 -2053708
rect -4033679 -2054177 -4033559 -2054172
rect -4033679 -2054277 -4033669 -2054177
rect -4033569 -2054277 -4033559 -2054177
rect -4033679 -2054282 -4033559 -2054277
rect -4034762 -2054377 -4034642 -2054372
rect -4034762 -2054477 -4034752 -2054377
rect -4034652 -2054477 -4034642 -2054377
rect -4034762 -2054482 -4034642 -2054477
rect -4029276 -2056390 -4029180 -2043984
rect -4029120 -2056190 -4029024 -2043535
rect -4028964 -2055988 -4028868 -2043088
rect -4028808 -2055790 -4028712 -2042621
rect -4028652 -2055590 -4028556 -2042189
rect -4028496 -2055388 -4028400 -2041687
rect -4028340 -2055188 -4028244 -2041162
rect -4028184 -2054987 -4028088 -2040681
rect -4028028 -2054788 -4027932 -2040181
rect -4027872 -2054589 -4027776 -2039982
rect -4027631 -2044907 -4027427 -2044902
rect -4027631 -2045091 -4027621 -2044907
rect -4027437 -2045091 -4027427 -2044907
rect -4027631 -2045096 -4027427 -2045091
rect -4027872 -2054662 -4027858 -2054589
rect -4027790 -2054662 -4027776 -2054589
rect -4027872 -2054676 -4027776 -2054662
rect -4028028 -2054861 -4028015 -2054788
rect -4027947 -2054861 -4027932 -2054788
rect -4028028 -2054875 -4027932 -2054861
rect -4028184 -2055060 -4028171 -2054987
rect -4028103 -2055060 -4028088 -2054987
rect -4028184 -2055074 -4028088 -2055060
rect -4028340 -2055261 -4028326 -2055188
rect -4028258 -2055261 -4028244 -2055188
rect -4028340 -2055275 -4028244 -2055261
rect -4028496 -2055461 -4028482 -2055388
rect -4028414 -2055461 -4028400 -2055388
rect -4028496 -2055476 -4028400 -2055461
rect -4028652 -2055663 -4028639 -2055590
rect -4028571 -2055663 -4028556 -2055590
rect -4028652 -2055677 -4028556 -2055663
rect -4028808 -2055863 -4028794 -2055790
rect -4028726 -2055863 -4028712 -2055790
rect -4028808 -2055876 -4028712 -2055863
rect -4028964 -2056061 -4028950 -2055988
rect -4028882 -2056061 -4028868 -2055988
rect -4028964 -2056075 -4028868 -2056061
rect -4029120 -2056263 -4029106 -2056190
rect -4029038 -2056263 -4029024 -2056190
rect -4029120 -2056276 -4029024 -2056263
rect -4029276 -2056463 -4029262 -2056390
rect -4029194 -2056463 -4029180 -2056390
rect -4029276 -2056476 -4029180 -2056463
rect -4039142 -2058465 -4039131 -2058387
rect -4039057 -2058465 -4039046 -2058387
rect -4039142 -2058475 -4039046 -2058465
rect -4040961 -2058675 -4040916 -2058577
rect -4040926 -2058677 -4040916 -2058675
rect -4040816 -2058675 -4040777 -2058577
rect -4040816 -2058677 -4040806 -2058675
rect -4040926 -2058682 -4040806 -2058677
rect -4041324 -2058876 -4041282 -2058777
rect -4041292 -2058877 -4041282 -2058876
rect -4041182 -2058876 -4041140 -2058777
rect -4041182 -2058877 -4041172 -2058876
rect -4041292 -2058882 -4041172 -2058877
rect -4041690 -2059077 -4041651 -2058977
rect -4041551 -2059077 -4041506 -2058977
rect -4041661 -2059082 -4041541 -2059077
rect -4042057 -2059277 -4042013 -2059177
rect -4041913 -2059277 -4041873 -2059177
rect -4042057 -2059278 -4041873 -2059277
rect -4042023 -2059282 -4041903 -2059278
rect -4042424 -2059475 -4042379 -2059377
rect -4042389 -2059477 -4042379 -2059475
rect -4042279 -2059475 -4042240 -2059377
rect -4042279 -2059477 -4042269 -2059475
rect -4042389 -2059482 -4042269 -2059477
rect -4027621 -2060377 -4027437 -2045096
rect -4027262 -2045407 -4027058 -2045402
rect -4027262 -2045591 -4027252 -2045407
rect -4027068 -2045591 -4027058 -2045407
rect -4027262 -2045596 -4027058 -2045591
rect -4027252 -2060177 -4027068 -2045596
rect -4026894 -2045907 -4026690 -2045902
rect -4026894 -2046091 -4026884 -2045907
rect -4026700 -2046091 -4026690 -2045907
rect -4026894 -2046096 -4026690 -2046091
rect -4026883 -2059977 -4026699 -2046096
rect -4026526 -2046407 -4026322 -2046402
rect -4026526 -2046591 -4026516 -2046407
rect -4026332 -2046591 -4026322 -2046407
rect -4026526 -2046596 -4026322 -2046591
rect -4026516 -2059777 -4026332 -2046596
rect -4026158 -2046907 -4025954 -2046902
rect -4026158 -2047091 -4026148 -2046907
rect -4025964 -2047091 -4025954 -2046907
rect -4026158 -2047096 -4025954 -2047091
rect -4026148 -2059577 -4025964 -2047096
rect -4026148 -2059676 -4026108 -2059577
rect -4026118 -2059677 -4026108 -2059676
rect -4026008 -2059676 -4025964 -2059577
rect -4026008 -2059677 -4025998 -2059676
rect -4026118 -2059682 -4025998 -2059677
rect -4026516 -2059877 -4026474 -2059777
rect -4026374 -2059877 -4026332 -2059777
rect -4026484 -2059882 -4026364 -2059877
rect -4026883 -2060077 -4026844 -2059977
rect -4026744 -2060077 -4026699 -2059977
rect -4026854 -2060082 -4026734 -2060077
rect -4027252 -2060275 -4027210 -2060177
rect -4027220 -2060277 -4027210 -2060275
rect -4027110 -2060275 -4027068 -2060177
rect -4027110 -2060277 -4027100 -2060275
rect -4027220 -2060282 -4027100 -2060277
rect -4027621 -2060476 -4027578 -2060377
rect -4027588 -2060477 -4027578 -2060476
rect -4027478 -2060476 -4027437 -2060377
rect -4027478 -2060477 -4027468 -2060476
rect -4027588 -2060482 -4027468 -2060477
rect -4038604 -2084022 -4038184 -2084017
rect -4038604 -2084143 -4038594 -2084022
rect -4038194 -2084143 -4038184 -2084022
rect -4038604 -2084148 -4038184 -2084143
rect -4038056 -2084258 -4037636 -2084253
rect -4038056 -2084359 -4038046 -2084258
rect -4037646 -2084359 -4037636 -2084258
rect -4038056 -2084364 -4037636 -2084359
rect -4037518 -2084458 -4037098 -2084453
rect -4037518 -2084559 -4037508 -2084458
rect -4037108 -2084559 -4037098 -2084458
rect -4037518 -2084564 -4037098 -2084559
rect -4036989 -2084658 -4036569 -2084653
rect -4036989 -2084759 -4036979 -2084658
rect -4036579 -2084759 -4036569 -2084658
rect -4036989 -2084764 -4036569 -2084759
rect -4036459 -2084858 -4036039 -2084853
rect -4036459 -2084959 -4036449 -2084858
rect -4036049 -2084959 -4036039 -2084858
rect -4036459 -2084964 -4036039 -2084959
rect -4035939 -2085058 -4035519 -2085053
rect -4035939 -2085159 -4035929 -2085058
rect -4035529 -2085159 -4035519 -2085058
rect -4035939 -2085164 -4035519 -2085159
rect -4035406 -2085259 -4034986 -2085254
rect -4035406 -2085360 -4035396 -2085259
rect -4034996 -2085360 -4034986 -2085259
rect -4035406 -2085365 -4034986 -2085360
rect -4034883 -2085458 -4034463 -2085453
rect -4034883 -2085559 -4034873 -2085458
rect -4034473 -2085559 -4034463 -2085458
rect -4034883 -2085564 -4034463 -2085559
rect -4034362 -2085658 -4033942 -2085653
rect -4034362 -2085759 -4034352 -2085658
rect -4033952 -2085759 -4033942 -2085658
rect -4034362 -2085764 -4033942 -2085759
rect -4033838 -2085858 -4033418 -2085853
rect -4033838 -2085959 -4033828 -2085858
rect -4033428 -2085959 -4033418 -2085858
rect -4033838 -2085964 -4033418 -2085959
rect -4033301 -2086058 -4032881 -2086053
rect -4033301 -2086159 -4033291 -2086058
rect -4032891 -2086159 -4032881 -2086058
rect -4033301 -2086164 -4032881 -2086159
rect -4031696 -2086659 -4031276 -2086654
rect -4031696 -2086760 -4031686 -2086659
rect -4031286 -2086760 -4031276 -2086659
rect -4031696 -2086765 -4031276 -2086760
rect -4031165 -2087059 -4030744 -2087054
rect -4031165 -2087159 -4031155 -2087059
rect -4030754 -2087159 -4030744 -2087059
rect -4031165 -2087164 -4030744 -2087159
rect -4068864 -2094421 -4066844 -2094416
rect -4045588 -2094421 -4043568 -2094416
rect -4068864 -2096421 -4068854 -2094421
rect -4066854 -2096421 -4045578 -2094421
rect -4043578 -2096421 -4043568 -2094421
rect -4068864 -2096426 -4066844 -2096421
rect -4045588 -2096426 -4043568 -2096421
rect -4024817 -2094421 -4022797 -2094416
rect -4001360 -2094421 -3999360 -2037831
rect -3998675 -2038066 -3998075 -2004627
rect -3997370 -2005230 -3995350 -2005225
rect -3997370 -2005414 -3997360 -2005230
rect -3995360 -2005414 -3995350 -2005230
rect -3997370 -2005419 -3995350 -2005414
rect -3997371 -2037242 -3995350 -2037237
rect -3997371 -2037426 -3997361 -2037242
rect -3995360 -2037426 -3995350 -2037242
rect -3997371 -2037431 -3995350 -2037426
rect -3998685 -2038071 -3998064 -2038066
rect -3998685 -2038255 -3998675 -2038071
rect -3998074 -2038255 -3998064 -2038071
rect -3998685 -2038260 -3998064 -2038255
rect -4024817 -2096421 -4024807 -2094421
rect -4022807 -2096421 -3999360 -2094421
rect -4024817 -2096426 -4022797 -2096421
rect -3998675 -2097504 -3998075 -2038260
rect -3993360 -2039273 -3991360 -1952431
rect -3993370 -2039278 -3991350 -2039273
rect -3993370 -2039462 -3993360 -2039278
rect -3991360 -2039462 -3991350 -2039278
rect -3993370 -2039467 -3991350 -2039462
rect -4070124 -2098104 -4032760 -2097504
rect -4032359 -2098104 -4032222 -2097504
rect -4031821 -2098104 -3998075 -2097504
rect -4072864 -2099361 -4070844 -2099356
rect -4072864 -2101361 -4072854 -2099361
rect -4070854 -2101361 -4070844 -2099361
rect -4072864 -2101366 -4070844 -2101361
rect -4045588 -2099361 -4043568 -2099356
rect -4045588 -2101361 -4045578 -2099361
rect -4043578 -2101361 -4043568 -2099361
rect -4045588 -2101366 -4043568 -2101361
rect -4024764 -2099361 -4022744 -2099356
rect -4024764 -2101361 -4024754 -2099361
rect -4022754 -2101361 -4022744 -2099361
rect -4024764 -2101366 -4022744 -2101361
rect -3997370 -2099361 -3995350 -2099356
rect -3997370 -2101361 -3997360 -2099361
rect -3995360 -2101361 -3995350 -2099361
rect -3997370 -2101366 -3995350 -2101361
rect -3993360 -2103832 -3991360 -2039467
rect -3993370 -2103837 -3991350 -2103832
rect -4076864 -2103911 -4074844 -2103906
rect -4076864 -2105911 -4076854 -2103911
rect -4074854 -2103913 -4074844 -2103911
rect -4045588 -2103913 -4043568 -2103908
rect -4074854 -2105911 -4045578 -2103913
rect -4076864 -2105916 -4074844 -2105911
rect -4074494 -2105913 -4045578 -2105911
rect -4043578 -2105913 -4043568 -2103913
rect -4045588 -2105918 -4043568 -2105913
rect -4024764 -2103913 -4022744 -2103908
rect -3993370 -2103913 -3993360 -2103837
rect -4024764 -2105913 -4024754 -2103913
rect -4022754 -2105837 -3993360 -2103913
rect -3991360 -2105837 -3991350 -2103837
rect -4022754 -2105842 -3991350 -2105837
rect -4022754 -2105913 -3991360 -2105842
rect -4024764 -2105918 -4022744 -2105913
rect -3993360 -2105914 -3991360 -2105913
rect -4080864 -2107846 -4078844 -2107841
rect -4080864 -2109846 -4080854 -2107846
rect -4078854 -2109846 -4078844 -2107846
rect -4080864 -2109851 -4078844 -2109846
rect -4045588 -2107845 -4043568 -2107840
rect -4045588 -2109845 -4045578 -2107845
rect -4043578 -2109845 -4043568 -2107845
rect -4045588 -2109850 -4043568 -2109845
rect -4024764 -2107845 -4022744 -2107840
rect -4024764 -2109845 -4024754 -2107845
rect -4022754 -2109845 -4022744 -2107845
rect -4024764 -2109850 -4022744 -2109845
rect -3989370 -2107845 -3987350 -2107840
rect -3989370 -2109845 -3989360 -2107845
rect -3987360 -2109845 -3987350 -2107845
rect -3989370 -2109850 -3987350 -2109845
rect -3985360 -2111753 -3983360 -1944628
rect -3985370 -2111758 -3983350 -2111753
rect -4084864 -2111976 -4082844 -2111971
rect -4045588 -2111976 -4043568 -2111971
rect -4084864 -2113976 -4084854 -2111976
rect -4082854 -2113976 -4045578 -2111976
rect -4043578 -2113976 -4043568 -2111976
rect -4084864 -2113981 -4082844 -2113976
rect -4045588 -2113981 -4043568 -2113976
rect -4024764 -2111976 -4022744 -2111971
rect -3985370 -2111976 -3985360 -2111758
rect -4024764 -2113976 -4024754 -2111976
rect -4022754 -2113758 -3985360 -2111976
rect -3983360 -2113758 -3983350 -2111758
rect -4022754 -2113763 -3983350 -2113758
rect -4022754 -2113975 -3983360 -2113763
rect -4022754 -2113976 -3984002 -2113975
rect -4024764 -2113981 -4022744 -2113976
rect -4088864 -2116206 -4086844 -2116201
rect -4088864 -2118206 -4088854 -2116206
rect -4086854 -2118206 -4086844 -2116206
rect -4088864 -2118211 -4086844 -2118206
rect -4045588 -2116206 -4043568 -2116201
rect -4045588 -2118206 -4045578 -2116206
rect -4043578 -2118206 -4043568 -2116206
rect -4045588 -2118211 -4043568 -2118206
rect -4024764 -2116206 -4022744 -2116201
rect -4024764 -2118206 -4024754 -2116206
rect -4022754 -2118206 -4022744 -2116206
rect -4024764 -2118211 -4022744 -2118206
rect -3981370 -2116206 -3979350 -2116201
rect -3981370 -2118206 -3981360 -2116206
rect -3979360 -2118206 -3979350 -2116206
rect -3981370 -2118211 -3979350 -2118206
<< via3 >>
rect -4088854 -1940121 -4086850 -1938117
rect -3981362 -1940119 -3979360 -1938117
rect -4080854 -1948414 -4078854 -1946414
rect -4037056 -1948414 -4036952 -1946414
rect -4031370 -1948414 -4031266 -1946414
rect -3989360 -1948416 -3987360 -1946416
rect -4080861 -2039463 -4078853 -2039277
rect -4088858 -2087559 -4086854 -2087459
rect -4088854 -2087959 -4086854 -2087859
rect -4088854 -2088359 -4086854 -2088259
rect -4072854 -1956224 -4070854 -1954224
rect -3997360 -1956224 -3995360 -1954224
rect -4072854 -1971819 -4070854 -1971635
rect -4072854 -2003840 -4070854 -2003655
rect -4072856 -2005416 -4070854 -2005232
rect -4072854 -2037427 -4070854 -2037243
rect -3997360 -1971819 -3995357 -1971635
rect -3997360 -2003826 -3995360 -2003642
rect -4038594 -2084143 -4038194 -2084022
rect -4038046 -2084359 -4037646 -2084258
rect -4037508 -2084559 -4037108 -2084458
rect -4036979 -2084759 -4036579 -2084658
rect -4036449 -2084959 -4036049 -2084858
rect -4035929 -2085159 -4035529 -2085058
rect -4035396 -2085360 -4034996 -2085259
rect -4034873 -2085559 -4034473 -2085458
rect -4034352 -2085759 -4033952 -2085658
rect -4033828 -2085959 -4033428 -2085858
rect -4033291 -2086159 -4032891 -2086058
rect -4031686 -2086760 -4031286 -2086659
rect -4031155 -2087159 -4030754 -2087059
rect -3997360 -2005414 -3995360 -2005230
rect -3997361 -2037426 -3995360 -2037242
rect -3993360 -2039462 -3991360 -2039278
rect -4072854 -2101361 -4070854 -2099361
rect -4045578 -2101361 -4043578 -2099361
rect -4024754 -2101361 -4022754 -2099361
rect -3997360 -2101361 -3995360 -2099361
rect -4080854 -2109846 -4078854 -2107846
rect -4045578 -2109845 -4043578 -2107845
rect -4024754 -2109845 -4022754 -2107845
rect -3989360 -2109845 -3987360 -2107845
rect -4088854 -2118206 -4086854 -2116206
rect -4045578 -2118206 -4043578 -2116206
rect -4024754 -2118206 -4022754 -2116206
rect -3981360 -2118206 -3979360 -2116206
<< metal4 >>
rect -4088855 -1938117 -4086849 -1938116
rect -3981363 -1938117 -3979359 -1938116
rect -4088855 -1940121 -4088854 -1938117
rect -4086850 -1940119 -3981362 -1938117
rect -3979360 -1940119 -3979359 -1938117
rect -4086850 -1940121 -4086849 -1940119
rect -3981363 -1940120 -3979359 -1940119
rect -4088855 -1940122 -4086849 -1940121
rect -4088854 -2087458 -4086854 -1940122
rect -4080855 -1946414 -4078853 -1946413
rect -4037057 -1946414 -4036951 -1946413
rect -4031371 -1946414 -4031265 -1946413
rect -4080855 -1948414 -4080854 -1946414
rect -4078854 -1948414 -4037056 -1946414
rect -4036952 -1948414 -4031370 -1946414
rect -4031266 -1946415 -3988451 -1946414
rect -4031266 -1946416 -3987359 -1946415
rect -4031266 -1948414 -3989360 -1946416
rect -4080855 -1948415 -4078853 -1948414
rect -4037057 -1948415 -4036951 -1948414
rect -4031371 -1948415 -4031265 -1948414
rect -4080854 -2039276 -4078854 -1948415
rect -3989361 -1948416 -3989360 -1948414
rect -3987360 -1948416 -3987359 -1946416
rect -3989361 -1948417 -3987359 -1948416
rect -4072855 -1954224 -4070853 -1954223
rect -3997361 -1954224 -3995359 -1954223
rect -4072855 -1956224 -4072854 -1954224
rect -4070854 -1956224 -3997360 -1954224
rect -3995360 -1956224 -3995359 -1954224
rect -4072855 -1956225 -4070853 -1956224
rect -3997361 -1956225 -3995359 -1956224
rect -4072854 -1971634 -4070854 -1956225
rect -3997360 -1971634 -3995360 -1956225
rect -4072855 -1971635 -4070853 -1971634
rect -4072855 -1971819 -4072854 -1971635
rect -4070854 -1971819 -4070853 -1971635
rect -4072855 -1971820 -4070853 -1971819
rect -3997361 -1971635 -3995356 -1971634
rect -3997361 -1971819 -3997360 -1971635
rect -3995357 -1971819 -3995356 -1971635
rect -3997361 -1971820 -3995356 -1971819
rect -4072854 -2003654 -4070854 -1971820
rect -3997360 -2003641 -3995360 -1971820
rect -3997361 -2003642 -3995359 -2003641
rect -4072855 -2003655 -4070853 -2003654
rect -4072855 -2003840 -4072854 -2003655
rect -4070854 -2003840 -4070853 -2003655
rect -3997361 -2003826 -3997360 -2003642
rect -3995360 -2003826 -3995359 -2003642
rect -3997361 -2003827 -3995359 -2003826
rect -4072855 -2003841 -4070853 -2003840
rect -4072854 -2005231 -4070854 -2003841
rect -3997360 -2005229 -3995360 -2003827
rect -3997361 -2005230 -3995359 -2005229
rect -4072857 -2005232 -4070853 -2005231
rect -4072857 -2005416 -4072856 -2005232
rect -4070854 -2005416 -4070853 -2005232
rect -3997361 -2005414 -3997360 -2005230
rect -3995360 -2005414 -3995359 -2005230
rect -3997361 -2005415 -3995359 -2005414
rect -4072857 -2005417 -4070853 -2005416
rect -4072854 -2037242 -4070854 -2005417
rect -3997360 -2037241 -3995360 -2005415
rect -3997362 -2037242 -3995359 -2037241
rect -4072855 -2037243 -4070853 -2037242
rect -4072855 -2037427 -4072854 -2037243
rect -4070854 -2037427 -4070853 -2037243
rect -3997362 -2037426 -3997361 -2037242
rect -3995360 -2037426 -3995359 -2037242
rect -3997362 -2037427 -3995359 -2037426
rect -4072855 -2037428 -4070853 -2037427
rect -4080862 -2039277 -4078852 -2039276
rect -4080862 -2039463 -4080861 -2039277
rect -4078853 -2039463 -4078852 -2039277
rect -4080862 -2039464 -4078852 -2039463
rect -4088859 -2087459 -4086853 -2087458
rect -4088859 -2087559 -4088858 -2087459
rect -4086854 -2087559 -4086853 -2087459
rect -4088859 -2087560 -4086853 -2087559
rect -4088854 -2087858 -4086854 -2087560
rect -4088855 -2087859 -4086853 -2087858
rect -4088855 -2087959 -4088854 -2087859
rect -4086854 -2087959 -4086853 -2087859
rect -4088855 -2087960 -4086853 -2087959
rect -4088854 -2088258 -4086854 -2087960
rect -4088855 -2088259 -4086853 -2088258
rect -4088855 -2088359 -4088854 -2088259
rect -4086854 -2088359 -4086853 -2088259
rect -4088855 -2088360 -4086853 -2088359
rect -4088854 -2116205 -4086854 -2088360
rect -4080854 -2107845 -4078854 -2039464
rect -4072854 -2099360 -4070854 -2037428
rect -4038595 -2084022 -4038193 -2084021
rect -4038595 -2084143 -4038594 -2084022
rect -4038194 -2084143 -4038193 -2084022
rect -4038595 -2084144 -4038193 -2084143
rect -4072855 -2099361 -4070853 -2099360
rect -4045579 -2099361 -4043577 -2099360
rect -4072855 -2101361 -4072854 -2099361
rect -4070854 -2101361 -4045578 -2099361
rect -4043578 -2101361 -4043577 -2099361
rect -4072855 -2101362 -4070853 -2101361
rect -4045579 -2101362 -4043577 -2101361
rect -4045579 -2107845 -4043577 -2107844
rect -4080855 -2107846 -4045578 -2107845
rect -4080855 -2109846 -4080854 -2107846
rect -4078854 -2109845 -4045578 -2107846
rect -4043578 -2109845 -4043577 -2107845
rect -4078854 -2109846 -4078853 -2109845
rect -4045579 -2109846 -4043577 -2109845
rect -4080855 -2109847 -4078853 -2109846
rect -4088855 -2116206 -4086853 -2116205
rect -4045579 -2116206 -4043577 -2116205
rect -4088855 -2118206 -4088854 -2116206
rect -4086854 -2118206 -4045578 -2116206
rect -4043578 -2118206 -4043577 -2116206
rect -4088855 -2118207 -4086853 -2118206
rect -4045579 -2118207 -4043577 -2118206
rect -4038594 -2125168 -4038194 -2084144
rect -4038047 -2084258 -4037645 -2084257
rect -4038047 -2084359 -4038046 -2084258
rect -4037646 -2084359 -4037645 -2084258
rect -4038047 -2084360 -4037645 -2084359
rect -4064847 -2125568 -4038194 -2125168
rect -4064847 -2125988 -4064451 -2125568
rect -4064851 -2142525 -4064451 -2125988
rect -4038046 -2126005 -4037646 -2084360
rect -4037508 -2084457 -4037108 -2084455
rect -4037509 -2084458 -4037107 -2084457
rect -4037509 -2084559 -4037508 -2084458
rect -4037108 -2084559 -4037107 -2084458
rect -4037509 -2084560 -4037107 -2084559
rect -4060336 -2126405 -4037646 -2126005
rect -4060336 -2142525 -4059936 -2126405
rect -4037508 -2126951 -4037108 -2084560
rect -4036980 -2084658 -4036578 -2084657
rect -4036980 -2084759 -4036979 -2084658
rect -4036579 -2084759 -4036578 -2084658
rect -4036980 -2084760 -4036578 -2084759
rect -4055876 -2127351 -4037108 -2126951
rect -4055876 -2142525 -4055476 -2127351
rect -4036979 -2127754 -4036579 -2084760
rect -4036450 -2084858 -4036048 -2084857
rect -4036450 -2084959 -4036449 -2084858
rect -4036049 -2084959 -4036048 -2084858
rect -4036450 -2084960 -4036048 -2084959
rect -4051552 -2128154 -4036579 -2127754
rect -4051552 -2142525 -4051152 -2128154
rect -4036449 -2128673 -4036049 -2084960
rect -4035930 -2085058 -4035528 -2085057
rect -4035930 -2085159 -4035929 -2085058
rect -4035529 -2085159 -4035528 -2085058
rect -4035930 -2085160 -4035528 -2085159
rect -4047282 -2129073 -4036049 -2128673
rect -4047282 -2142525 -4046882 -2129073
rect -4035929 -2129537 -4035529 -2085160
rect -4035397 -2085259 -4034995 -2085258
rect -4035397 -2085360 -4035396 -2085259
rect -4034996 -2085360 -4034995 -2085259
rect -4035397 -2085361 -4034995 -2085360
rect -4043323 -2129937 -4035529 -2129537
rect -4043323 -2142525 -4042923 -2129937
rect -4035396 -2130346 -4034996 -2085361
rect -4034874 -2085458 -4034472 -2085457
rect -4034874 -2085559 -4034873 -2085458
rect -4034473 -2085559 -4034472 -2085458
rect -4034874 -2085560 -4034472 -2085559
rect -4038799 -2130746 -4034996 -2130346
rect -4038799 -2142525 -4038399 -2130746
rect -4034873 -2142525 -4034472 -2085560
rect -4034353 -2085658 -4033951 -2085657
rect -4034353 -2085759 -4034352 -2085658
rect -4033952 -2085759 -4033951 -2085658
rect -4034353 -2085760 -4033951 -2085759
rect -4034352 -2130349 -4033951 -2085760
rect -4033829 -2085858 -4033427 -2085857
rect -4033829 -2085959 -4033828 -2085858
rect -4033428 -2085959 -4033427 -2085858
rect -4033829 -2085960 -4033427 -2085959
rect -4033828 -2129568 -4033427 -2085960
rect -4033292 -2086058 -4032890 -2086057
rect -4033292 -2086159 -4033291 -2086058
rect -4032891 -2086159 -4032890 -2086058
rect -4033292 -2086160 -4032890 -2086159
rect -4033291 -2128678 -4032890 -2086160
rect -4031687 -2086659 -4031285 -2086658
rect -4031687 -2086760 -4031686 -2086659
rect -4031286 -2086760 -4031285 -2086659
rect -4031687 -2086761 -4031285 -2086760
rect -4031686 -2126021 -4031285 -2086761
rect -4031156 -2087059 -4030753 -2087058
rect -4031156 -2087159 -4031155 -2087059
rect -4030754 -2087159 -4030753 -2087059
rect -4031156 -2087160 -4030753 -2087159
rect -4031155 -2125186 -4030754 -2087160
rect -3997360 -2099360 -3995360 -2037427
rect -3993361 -2039278 -3991359 -2039277
rect -3993361 -2039462 -3993360 -2039278
rect -3991360 -2039462 -3991359 -2039278
rect -3993361 -2039463 -3991359 -2039462
rect -4024755 -2099361 -4022753 -2099360
rect -3997361 -2099361 -3995359 -2099360
rect -4024755 -2101361 -4024754 -2099361
rect -4022754 -2101361 -3997360 -2099361
rect -3995360 -2101361 -3995359 -2099361
rect -4024755 -2101362 -4022753 -2101361
rect -3997361 -2101362 -3995359 -2101361
rect -3989360 -2107844 -3987360 -1948417
rect -4024755 -2107845 -4022753 -2107844
rect -3989361 -2107845 -3987359 -2107844
rect -4024755 -2109845 -4024754 -2107845
rect -4022754 -2109845 -3989360 -2107845
rect -3987360 -2109845 -3987359 -2107845
rect -4024755 -2109846 -4022753 -2109845
rect -3989361 -2109846 -3987359 -2109845
rect -3981360 -2116205 -3979360 -1940120
rect -4024755 -2116206 -4022753 -2116205
rect -3981361 -2116206 -3979359 -2116205
rect -4024755 -2118206 -4024754 -2116206
rect -4022754 -2118206 -3981360 -2116206
rect -3979360 -2118206 -3979359 -2116206
rect -4024755 -2118207 -4022753 -2118206
rect -3981361 -2118207 -3979359 -2118206
rect -4031155 -2125587 -4005528 -2125186
rect -4031686 -2126422 -4010103 -2126021
rect -4033291 -2129079 -4022498 -2128678
rect -4033828 -2129969 -4026484 -2129568
rect -4034352 -2130750 -4030565 -2130349
rect -4030966 -2142525 -4030565 -2130750
rect -4026885 -2142525 -4026484 -2129969
rect -4022899 -2142525 -4022498 -2129079
rect -4010504 -2142525 -4010103 -2126422
rect -4005929 -2142525 -4005528 -2125587
use analog_block  analog_block_0
timestamp 1731349849
transform 0 -1 -4003743 1 0 -2038012
box -15790 -954 74799 61971
use sar  sar_0
timestamp 1731350402
transform 0 1 -4029800 1 0 -2071803
box -16648 -13778 17740 5046
<< labels >>
flabel metal2 -4034716 -1936685 -4034656 -1936511 0 FreeSans 320 0 0 0 VIP
port 28 nsew
flabel metal2 -4033670 -1936677 -4033610 -1936503 0 FreeSans 320 0 0 0 VIN
port 29 nsew
flabel metal3 -4055120 -2095857 -4054592 -2095482 0 FreeSans 4800 0 0 0 VSSR
port 30 nsew
flabel metal3 -4055075 -2097974 -4054547 -2097599 0 FreeSans 4800 0 0 0 VCM
port 31 nsew
flabel metal4 -4055075 -2100551 -4054547 -2100176 0 FreeSans 4800 0 0 0 VDDR
port 32 nsew
flabel metal3 -4055075 -2105261 -4054547 -2104886 0 FreeSans 4800 0 0 0 VSSA
port 33 nsew
flabel metal4 -4055075 -2108971 -4054547 -2108596 0 FreeSans 4800 0 0 0 VDDA
port 34 nsew
flabel metal3 -4055097 -2113192 -4054569 -2112817 0 FreeSans 4800 0 0 0 VSSD
port 35 nsew
flabel metal4 -4055053 -2117324 -4054525 -2116949 0 FreeSans 4800 0 0 0 VDDD
port 36 nsew
flabel metal4 -4064806 -2142428 -4064561 -2142228 0 FreeSans 3200 0 0 0 CKO
port 37 nsew
flabel metal4 -4060251 -2142450 -4060006 -2142250 0 FreeSans 3200 0 0 0 DOUT[0]
port 38 nsew
flabel metal4 -4055776 -2142415 -4055531 -2142215 0 FreeSans 3200 0 0 0 DOUT[1]
port 39 nsew
flabel metal4 -4051483 -2142392 -4051238 -2142192 0 FreeSans 3200 0 0 0 DOUT[2]
port 40 nsew
flabel metal4 -4047168 -2142392 -4046923 -2142192 0 FreeSans 3200 0 0 0 DOUT[3]
port 41 nsew
flabel metal4 -4043235 -2142370 -4042990 -2142170 0 FreeSans 3200 0 0 0 DOUT[4]
port 42 nsew
flabel metal4 -4038695 -2142392 -4038450 -2142192 0 FreeSans 3200 0 0 0 DOUT[5]
port 43 nsew
flabel metal4 -4034785 -2142370 -4034540 -2142170 0 FreeSans 3200 0 0 0 DOUT[6]
port 44 nsew
flabel metal4 -4030897 -2142370 -4030652 -2142170 0 FreeSans 3200 0 0 0 DOUT[7]
port 45 nsew
flabel metal4 -4026784 -2142370 -4026539 -2142170 0 FreeSans 3200 0 0 0 DOUT[8]
port 46 nsew
flabel metal4 -4022806 -2142370 -4022561 -2142170 0 FreeSans 3200 0 0 0 DOUT[9]
port 47 nsew
flabel metal4 -4010423 -2142378 -4010178 -2142178 0 FreeSans 3200 0 0 0 CLK
port 50 nsew
flabel metal4 -4005842 -2142401 -4005597 -2142201 0 FreeSans 3200 0 0 0 EN
port 51 nsew
<< end >>
