magic
tech sky130A
magscale 1 2
<<<<<<< HEAD
timestamp 1730798039
=======
timestamp 1730796434
<< error_s >>
rect 2334 -386 2502 -126
rect 1502 -526 1902 -386
rect 2334 -526 2734 -386
rect 1502 -834 1902 -694
rect 2334 -834 2734 -694
rect 2334 -1094 2502 -834
>>>>>>> 2788aa0 (update)
<< metal3 >>
rect 3186 -654 3246 -403
<< metal4 >>
rect 2553 -815 2613 -335
use sky130_fd_pr__cap_mim_m3_1_UCPR8Z  sky130_fd_pr__cap_mim_m3_1_UCPR8Z_0
timestamp 1730777901
transform 1 0 1848 0 1 -174
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_VCTT89  sky130_fd_pr__cap_mim_m3_1_VCTT89_0
<<<<<<< HEAD
timestamp 1730797230
transform 1 0 2860 0 1 -894
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_VCTT89  sky130_fd_pr__cap_mim_m3_1_VCTT89_1
timestamp 1730797230
transform 1 0 2860 0 1 -174
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_VCTT89  XC2
timestamp 1730797230
=======
timestamp 1730269323
transform 1 0 2680 0 1 -894
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_VCTT89  sky130_fd_pr__cap_mim_m3_1_VCTT89_1
timestamp 1730269323
transform 1 0 2680 0 1 -326
box -386 -240 386 240
use sky130_fd_pr__cap_mim_m3_1_VCTT89  XC2
timestamp 1730269323
>>>>>>> 2788aa0 (update)
transform 1 0 1848 0 1 -894
box -386 -240 386 240
<< labels >>
flabel metal4 s 1703 -174 1703 -174 0 FreeSans 320 0 0 0 VPBT1
port 1 nsew
flabel metal3 s 2043 -172 2043 -172 0 FreeSans 320 0 0 0 VNBT1
port 2 nsew
flabel metal4 s 1698 -895 1698 -895 0 FreeSans 320 0 0 0 VPBT2
port 3 nsew
flabel metal4 s 2713 -174 2713 -174 0 FreeSans 320 0 0 0 VPBT3
port 4 nsew
flabel metal3 s 3085 -174 3085 -174 0 FreeSans 320 0 0 0 VNBT3
port 5 nsew
flabel metal3 s 2050 -899 2050 -899 0 FreeSans 320 0 0 0 CLKS
port 6 nsew
<< end >>
