magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect 716 -3234 750 -3158
rect 716 -3324 750 -3318
rect 1102 -3234 1136 -3158
rect 1102 -3324 1136 -3318
rect 1488 -3234 1522 -3158
rect 1488 -3324 1522 -3318
rect 1594 -3358 1628 -3158
rect 1594 -3448 1628 -3442
rect 1980 -3358 2014 -3158
rect 1980 -3448 2014 -3442
rect 2366 -3358 2400 -3158
rect 2366 -3448 2400 -3442
<< viali >>
rect 716 -3318 750 -3234
rect 1102 -3318 1136 -3234
rect 1488 -3318 1522 -3234
rect 1594 -3442 1628 -3358
rect 1980 -3442 2014 -3358
rect 2366 -3442 2400 -3358
<< metal1 >>
rect 880 -2135 900 -2083
rect 952 -2135 972 -2083
rect 1265 -2135 1286 -2083
rect 1338 -2135 1357 -2083
rect 810 -2225 816 -2173
rect 868 -2225 874 -2173
rect 810 -2298 874 -2225
rect 810 -2350 816 -2298
rect 868 -2350 874 -2298
rect 810 -2421 874 -2350
rect 810 -2473 816 -2421
rect 868 -2473 874 -2421
rect 978 -2225 984 -2173
rect 1036 -2225 1202 -2173
rect 1254 -2225 1260 -2173
rect 978 -2298 1260 -2225
rect 978 -2350 984 -2298
rect 1036 -2350 1202 -2298
rect 1254 -2350 1260 -2298
rect 978 -2421 1260 -2350
rect 978 -2473 984 -2421
rect 1036 -2473 1202 -2421
rect 1254 -2473 1260 -2421
rect 1364 -2225 1370 -2173
rect 1422 -2225 1428 -2173
rect 1364 -2298 1428 -2225
rect 1364 -2350 1370 -2298
rect 1422 -2350 1428 -2298
rect 1364 -2421 1428 -2350
rect 1364 -2473 1370 -2421
rect 1422 -2473 1428 -2421
rect 880 -2563 900 -2511
rect 952 -2563 972 -2511
rect 1266 -2563 1286 -2511
rect 1338 -2563 1358 -2511
rect 1758 -2571 1778 -2519
rect 1830 -2571 1850 -2519
rect 2144 -2571 2164 -2519
rect 2216 -2571 2236 -2519
rect 880 -2671 900 -2619
rect 952 -2671 972 -2619
rect 1266 -2671 1286 -2619
rect 1338 -2671 1358 -2619
rect 1688 -2648 1752 -2600
rect 1688 -2700 1694 -2648
rect 1746 -2700 1752 -2648
rect 1856 -2648 2138 -2600
rect 1856 -2700 1862 -2648
rect 1914 -2700 2080 -2648
rect 2132 -2700 2138 -2648
rect 2242 -2648 2306 -2600
rect 2242 -2700 2248 -2648
rect 2300 -2700 2306 -2648
rect 810 -2761 816 -2709
rect 868 -2761 874 -2709
rect 810 -2833 874 -2761
rect 810 -2885 816 -2833
rect 868 -2885 874 -2833
rect 810 -2957 874 -2885
rect 810 -3009 816 -2957
rect 868 -3009 874 -2957
rect 978 -2761 984 -2709
rect 1036 -2761 1202 -2709
rect 1254 -2761 1260 -2709
rect 978 -2833 1260 -2761
rect 978 -2885 984 -2833
rect 1036 -2885 1202 -2833
rect 1254 -2885 1260 -2833
rect 978 -2957 1260 -2885
rect 978 -3009 984 -2957
rect 1036 -3009 1202 -2957
rect 1254 -3009 1260 -2957
rect 1364 -2761 1370 -2709
rect 1422 -2761 1428 -2709
rect 1364 -2833 1428 -2761
rect 1758 -2781 1778 -2729
rect 1830 -2781 1850 -2729
rect 2144 -2781 2164 -2729
rect 2216 -2781 2236 -2729
rect 1364 -2885 1370 -2833
rect 1422 -2885 1428 -2833
rect 1364 -2918 1428 -2885
rect 1758 -2889 1778 -2837
rect 1830 -2889 1850 -2837
rect 2144 -2889 2164 -2837
rect 2216 -2889 2236 -2837
rect 1364 -2957 1752 -2918
rect 1364 -3009 1370 -2957
rect 1422 -2966 1752 -2957
rect 1422 -3009 1694 -2966
rect 1364 -3018 1694 -3009
rect 1746 -3018 1752 -2966
rect 1856 -2966 2138 -2918
rect 1856 -3018 1862 -2966
rect 1914 -3018 2080 -2966
rect 2132 -3018 2138 -2966
rect 2242 -2966 2306 -2918
rect 2242 -3018 2248 -2966
rect 2300 -3018 2306 -2966
rect 880 -3099 900 -3047
rect 952 -3099 972 -3047
rect 1266 -3099 1286 -3047
rect 1338 -3099 1358 -3047
rect 1758 -3099 1778 -3047
rect 1830 -3099 1850 -3047
rect 2144 -3099 2164 -3047
rect 2216 -3099 2236 -3047
rect 894 -3185 900 -3133
rect 952 -3185 2164 -3133
rect 894 -3191 2164 -3185
rect 2216 -3191 2222 -3133
rect 680 -3234 816 -3228
rect 680 -3318 716 -3234
rect 750 -3318 816 -3234
rect 868 -3234 2436 -3228
rect 868 -3318 1102 -3234
rect 1136 -3318 1488 -3234
rect 1522 -3318 2436 -3234
rect 680 -3324 2436 -3318
rect 680 -3358 2248 -3352
rect 680 -3442 1594 -3358
rect 1628 -3442 1980 -3358
rect 2014 -3442 2248 -3358
rect 2300 -3358 2436 -3352
rect 2300 -3442 2366 -3358
rect 2400 -3442 2436 -3358
rect 680 -3448 2436 -3442
<< via1 >>
rect 900 -2135 952 -2083
rect 1286 -2135 1338 -2083
rect 816 -2225 868 -2173
rect 816 -2350 868 -2298
rect 816 -2473 868 -2421
rect 984 -2225 1036 -2173
rect 1202 -2225 1254 -2173
rect 984 -2350 1036 -2298
rect 1202 -2350 1254 -2298
rect 984 -2473 1036 -2421
rect 1202 -2473 1254 -2421
rect 1370 -2225 1422 -2173
rect 1370 -2350 1422 -2298
rect 1370 -2473 1422 -2421
rect 900 -2563 952 -2511
rect 1286 -2563 1338 -2511
rect 1778 -2571 1830 -2519
rect 2164 -2571 2216 -2519
rect 900 -2671 952 -2619
rect 1286 -2671 1338 -2619
rect 1694 -2700 1746 -2648
rect 1862 -2700 1914 -2648
rect 2080 -2700 2132 -2648
rect 2248 -2700 2300 -2648
rect 816 -2761 868 -2709
rect 816 -2885 868 -2833
rect 816 -3009 868 -2957
rect 984 -2761 1036 -2709
rect 1202 -2761 1254 -2709
rect 984 -2885 1036 -2833
rect 1202 -2885 1254 -2833
rect 984 -3009 1036 -2957
rect 1202 -3009 1254 -2957
rect 1370 -2761 1422 -2709
rect 1778 -2781 1830 -2729
rect 2164 -2781 2216 -2729
rect 1370 -2885 1422 -2833
rect 1778 -2889 1830 -2837
rect 2164 -2889 2216 -2837
rect 1370 -3009 1422 -2957
rect 1694 -3018 1746 -2966
rect 1862 -3018 1914 -2966
rect 2080 -3018 2132 -2966
rect 2248 -3018 2300 -2966
rect 900 -3099 952 -3047
rect 1286 -3099 1338 -3047
rect 1778 -3099 1830 -3047
rect 2164 -3099 2216 -3047
rect 900 -3185 952 -3133
rect 2164 -3191 2216 -3133
rect 816 -3318 868 -3228
rect 2248 -3442 2300 -3352
<< metal2 >>
rect 898 -2083 954 -2077
rect 898 -2135 900 -2083
rect 952 -2135 954 -2083
rect 814 -2173 870 -2167
rect 814 -2225 816 -2173
rect 868 -2225 870 -2173
rect 814 -2298 870 -2225
rect 814 -2350 816 -2298
rect 868 -2350 870 -2298
rect 814 -2421 870 -2350
rect 814 -2473 816 -2421
rect 868 -2473 870 -2421
rect 814 -2709 870 -2473
rect 814 -2761 816 -2709
rect 868 -2761 870 -2709
rect 814 -2833 870 -2761
rect 814 -2885 816 -2833
rect 868 -2885 870 -2833
rect 814 -2957 870 -2885
rect 814 -3009 816 -2957
rect 868 -3009 870 -2957
rect 814 -3228 870 -3009
rect 898 -2511 954 -2135
rect 1284 -2083 1340 -2077
rect 1284 -2135 1286 -2083
rect 1338 -2135 1340 -2083
rect 898 -2563 900 -2511
rect 952 -2563 954 -2511
rect 898 -2619 954 -2563
rect 898 -2671 900 -2619
rect 952 -2671 954 -2619
rect 898 -3047 954 -2671
rect 982 -2173 1038 -2167
rect 982 -2225 984 -2173
rect 1036 -2225 1038 -2173
rect 982 -2298 1038 -2225
rect 982 -2350 984 -2298
rect 1036 -2350 1038 -2298
rect 982 -2421 1038 -2350
rect 982 -2473 984 -2421
rect 1036 -2473 1038 -2421
rect 982 -2709 1038 -2473
rect 982 -2761 984 -2709
rect 1036 -2761 1038 -2709
rect 982 -2833 1038 -2761
rect 982 -2885 984 -2833
rect 1036 -2885 1038 -2833
rect 982 -2957 1038 -2885
rect 982 -3009 984 -2957
rect 1036 -3009 1038 -2957
rect 982 -3015 1038 -3009
rect 1200 -2173 1256 -2167
rect 1200 -2225 1202 -2173
rect 1254 -2225 1256 -2173
rect 1200 -2298 1256 -2225
rect 1200 -2350 1202 -2298
rect 1254 -2350 1256 -2298
rect 1200 -2421 1256 -2350
rect 1200 -2473 1202 -2421
rect 1254 -2473 1256 -2421
rect 1200 -2709 1256 -2473
rect 1200 -2761 1202 -2709
rect 1254 -2761 1256 -2709
rect 1200 -2833 1256 -2761
rect 1200 -2885 1202 -2833
rect 1254 -2885 1256 -2833
rect 1200 -2957 1256 -2885
rect 1200 -3009 1202 -2957
rect 1254 -3009 1256 -2957
rect 1200 -3015 1256 -3009
rect 1284 -2511 1340 -2135
rect 1284 -2563 1286 -2511
rect 1338 -2563 1340 -2511
rect 1284 -2619 1340 -2563
rect 1284 -2671 1286 -2619
rect 1338 -2671 1340 -2619
rect 898 -3099 900 -3047
rect 952 -3099 954 -3047
rect 898 -3133 954 -3099
rect 1284 -3047 1340 -2671
rect 1368 -2173 1424 -2167
rect 1368 -2225 1370 -2173
rect 1422 -2225 1424 -2173
rect 1368 -2298 1424 -2225
rect 1368 -2350 1370 -2298
rect 1422 -2350 1424 -2298
rect 1368 -2421 1424 -2350
rect 1368 -2473 1370 -2421
rect 1422 -2473 1424 -2421
rect 1368 -2709 1424 -2473
rect 1776 -2519 1832 -2513
rect 1776 -2571 1778 -2519
rect 1830 -2571 1832 -2519
rect 1368 -2761 1370 -2709
rect 1422 -2761 1424 -2709
rect 1368 -2833 1424 -2761
rect 1368 -2885 1370 -2833
rect 1422 -2885 1424 -2833
rect 1368 -2957 1424 -2885
rect 1368 -3009 1370 -2957
rect 1422 -3009 1424 -2957
rect 1368 -3015 1424 -3009
rect 1692 -2648 1748 -2642
rect 1692 -2700 1694 -2648
rect 1746 -2700 1748 -2648
rect 1692 -2966 1748 -2700
rect 1692 -3018 1694 -2966
rect 1746 -3018 1748 -2966
rect 1692 -3024 1748 -3018
rect 1776 -2729 1832 -2571
rect 2162 -2519 2218 -2513
rect 2162 -2571 2164 -2519
rect 2216 -2571 2218 -2519
rect 1776 -2781 1778 -2729
rect 1830 -2781 1832 -2729
rect 1776 -2837 1832 -2781
rect 1776 -2889 1778 -2837
rect 1830 -2889 1832 -2837
rect 1284 -3099 1286 -3047
rect 1338 -3099 1340 -3047
rect 1284 -3105 1340 -3099
rect 1776 -3047 1832 -2889
rect 1860 -2648 1916 -2642
rect 1860 -2700 1862 -2648
rect 1914 -2700 1916 -2648
rect 1860 -2966 1916 -2700
rect 1860 -3018 1862 -2966
rect 1914 -3018 1916 -2966
rect 1860 -3024 1916 -3018
rect 2078 -2648 2134 -2642
rect 2078 -2700 2080 -2648
rect 2132 -2700 2134 -2648
rect 2078 -2966 2134 -2700
rect 2078 -3018 2080 -2966
rect 2132 -3018 2134 -2966
rect 2078 -3024 2134 -3018
rect 2162 -2729 2218 -2571
rect 2162 -2781 2164 -2729
rect 2216 -2781 2218 -2729
rect 2162 -2837 2218 -2781
rect 2162 -2889 2164 -2837
rect 2216 -2889 2218 -2837
rect 1776 -3099 1778 -3047
rect 1830 -3099 1832 -3047
rect 1776 -3105 1832 -3099
rect 2162 -3047 2218 -2889
rect 2162 -3099 2164 -3047
rect 2216 -3099 2218 -3047
rect 898 -3185 900 -3133
rect 952 -3185 954 -3133
rect 898 -3191 954 -3185
rect 2162 -3133 2218 -3099
rect 2162 -3191 2164 -3133
rect 2216 -3191 2218 -3133
rect 2162 -3197 2218 -3191
rect 2246 -2648 2302 -2642
rect 2246 -2700 2248 -2648
rect 2300 -2700 2302 -2648
rect 2246 -2966 2302 -2700
rect 2246 -3018 2248 -2966
rect 2300 -3018 2302 -2966
rect 814 -3318 816 -3228
rect 868 -3318 870 -3228
rect 814 -3324 870 -3318
rect 2246 -3352 2302 -3018
rect 2246 -3442 2248 -3352
rect 2300 -3442 2302 -3352
rect 2246 -3448 2302 -3442
use sky130_fd_pr__pfet_01v8_TMYQY6  XM1
timestamp 1730624594
transform 1 0 926 0 1 -2591
box -246 -637 246 637
use sky130_fd_pr__pfet_01v8_TMYQY6  XM2
timestamp 1730624594
transform 1 0 1312 0 1 -2591
box -246 -637 246 637
use sky130_fd_pr__nfet_01v8_DJGLWN  XM3
timestamp 1730624594
transform 1 0 1804 0 1 -2809
box -246 -419 246 419
use sky130_fd_pr__nfet_01v8_DJGLWN  XM4
timestamp 1730624594
transform 1 0 2190 0 1 -2809
box -246 -419 246 419
<< labels >>
flabel via1 1286 -3099 1338 -3047 0 FreeSans 320 0 0 0 ckb
port 4 nsew
flabel via1 1778 -3099 1830 -3047 0 FreeSans 320 0 0 0 ck
port 3 nsew
flabel metal1 680 -3324 776 -3228 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel metal1 680 -3448 776 -3352 0 FreeSans 320 0 0 0 vssa
port 5 nsew
flabel via1 1370 -2225 1422 -2173 0 FreeSans 320 0 0 0 out
port 6 nsew
flabel via1 2164 -2571 2216 -2519 0 FreeSans 320 0 0 0 in
port 2 nsew
<< end >>
