magic
tech sky130A
magscale 1 2
timestamp 1727309470
<< error_s >>
rect 1921 509 1979 515
rect 1921 475 1933 509
rect 1921 469 1979 475
rect 1921 81 1979 87
rect 1921 47 1933 81
rect 1921 41 1979 47
rect 2374 -88 2415 650
rect 2556 512 2614 518
rect 2872 512 2930 518
rect 2556 478 2568 512
rect 2872 478 2884 512
rect 2556 472 2614 478
rect 2872 472 2930 478
rect 2556 84 2614 90
rect 2872 84 2930 90
rect 2556 50 2568 84
rect 2872 50 2884 84
rect 2556 44 2614 50
rect 2872 44 2930 50
rect 2240 -306 2298 -300
rect 2556 -306 2614 -300
rect 2872 -306 2930 -300
rect 2240 -340 2252 -306
rect 2556 -340 2568 -306
rect 2872 -340 2884 -306
rect 2240 -346 2298 -340
rect 2556 -346 2614 -340
rect 2872 -346 2930 -340
rect 2240 -616 2298 -610
rect 2556 -616 2614 -610
rect 2872 -616 2930 -610
rect 2240 -650 2252 -616
rect 2556 -650 2568 -616
rect 2872 -650 2884 -616
rect 2240 -656 2298 -650
rect 2556 -656 2614 -650
rect 2872 -656 2930 -650
rect 1924 -820 1982 -814
rect 2240 -820 2298 -814
rect 2556 -820 2614 -814
rect 2872 -820 2930 -814
rect 1924 -854 1936 -820
rect 2240 -854 2252 -820
rect 2556 -854 2568 -820
rect 2872 -854 2884 -820
rect 1924 -860 1982 -854
rect 2240 -860 2298 -854
rect 2556 -860 2614 -854
rect 2872 -860 2930 -854
rect 1924 -1130 1982 -1124
rect 2240 -1130 2298 -1124
rect 2556 -1130 2614 -1124
rect 2872 -1130 2930 -1124
rect 1924 -1164 1936 -1130
rect 2240 -1164 2252 -1130
rect 2556 -1164 2568 -1130
rect 2872 -1164 2884 -1130
rect 1924 -1170 1982 -1164
rect 2240 -1170 2298 -1164
rect 2556 -1170 2614 -1164
rect 2872 -1170 2930 -1164
<< viali >>
rect 3042 -656 3076 -300
<< metal1 >>
rect 3036 -300 3082 -288
rect 3036 -378 3042 -300
rect 2290 -578 2390 -378
rect 2606 -578 2880 -378
rect 2922 -578 3042 -378
rect 2340 -892 2390 -578
rect 3036 -656 3042 -578
rect 3076 -656 3082 -300
rect 3036 -668 3082 -656
rect 2290 -1092 2564 -892
rect 2606 -1092 2880 -892
use sky130_fd_pr__cap_mim_m3_1_K22CKP  sky130_fd_pr__cap_mim_m3_1_K22CKP_0
timestamp 1727309470
transform 0 1 618 -1 0 -269
box -386 -240 386 240
use sky130_fd_pr__pfet_01v8_J4PGPS  XM1
timestamp 1727309470
transform 1 0 1950 0 1 278
box -211 -369 211 369
use sky130_fd_pr__pfet_01v8_J4PGPS  XM2
timestamp 1727309470
transform 1 0 2585 0 1 281
box -211 -369 211 369
use sky130_fd_pr__pfet_01v8_J4PGPS  XM3
timestamp 1727309470
transform 1 0 2901 0 1 281
box -211 -369 211 369
use sky130_fd_pr__nfet_01v8_TGNW9T  XM4
timestamp 1727309470
transform 1 0 1953 0 1 -992
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM5
timestamp 1727309470
transform 1 0 2269 0 1 -992
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM6
timestamp 1727309470
transform 1 0 2269 0 1 -478
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM7
timestamp 1727309470
transform -1 0 2585 0 1 -992
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM8
timestamp 1727309470
transform -1 0 2585 0 1 -478
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM9
timestamp 1727309470
transform -1 0 2901 0 1 -478
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_TGNW9T  XM10
timestamp 1727309470
transform 1 0 2901 0 1 -992
box -211 -310 211 310
<< end >>
