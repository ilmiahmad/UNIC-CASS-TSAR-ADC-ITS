magic
tech sky130A
magscale 1 2
timestamp 1730745419
<< nwell >>
rect -1201 496 -1138 582
rect -1201 293 -1111 496
rect -1201 261 -1138 293
rect -1201 -582 -1132 -261
<< pwell >>
rect -1201 48 -1100 203
rect -1201 -48 19311 48
rect -1201 -203 -1100 -48
<< psubdiff >>
rect -1165 48 -1131 129
rect -1165 -129 -1131 -48
<< nsubdiff >>
rect -1165 445 -1131 479
rect -1165 309 -1131 343
rect -1165 -343 -1131 -309
rect -1165 -479 -1131 -445
<< psubdiffcont >>
rect -1165 -48 -1131 48
<< nsubdiffcont >>
rect -1165 343 -1131 445
rect -1165 -445 -1131 -343
<< locali >>
rect -1165 445 -1131 479
rect -1165 309 -1131 343
rect -1165 48 -1131 129
rect -1131 -17 -1075 17
rect -1165 -129 -1131 -48
rect -1165 -343 -1131 -309
rect -1165 -479 -1131 -445
<< viali >>
rect -1165 343 -1131 445
rect -229 427 -195 461
rect 302 427 336 461
rect 2234 427 2268 461
rect 4166 427 4200 461
rect 6098 427 6132 461
rect 8030 427 8064 461
rect 9962 427 9996 461
rect 11894 428 11928 462
rect 13826 428 13860 462
rect 15758 427 15792 461
rect 17690 427 17724 461
rect 1776 289 1810 323
rect 3708 289 3742 323
rect 5640 289 5674 323
rect 7572 289 7606 323
rect 9504 289 9538 323
rect 11436 289 11470 323
rect 13368 289 13402 323
rect 15300 289 15334 323
rect 17232 289 17266 323
rect 19164 289 19198 323
rect 30 221 64 255
rect 1962 221 1996 255
rect 3894 221 3928 255
rect 5826 221 5860 255
rect 7758 221 7792 255
rect 9690 221 9724 255
rect 11622 221 11656 255
rect 13554 221 13588 255
rect 15486 221 15520 255
rect 17418 221 17452 255
rect -1165 -48 -1131 48
rect 30 -255 64 -221
rect 1962 -255 1996 -221
rect 3894 -255 3928 -221
rect 5826 -255 5860 -221
rect 7758 -255 7792 -221
rect 9690 -255 9724 -221
rect 11622 -255 11656 -221
rect 13554 -255 13588 -221
rect 15486 -255 15520 -221
rect 17418 -255 17452 -221
rect 1776 -323 1810 -289
rect 3708 -323 3742 -289
rect 5640 -323 5674 -289
rect 7572 -323 7606 -289
rect 9504 -323 9538 -289
rect 11436 -323 11470 -289
rect 13368 -323 13402 -289
rect 15300 -323 15334 -289
rect 17232 -323 17266 -289
rect 19164 -323 19198 -289
rect -1165 -445 -1131 -343
rect -229 -461 -195 -427
rect 302 -461 336 -427
rect 2234 -461 2268 -427
rect 4166 -461 4200 -427
rect 6098 -461 6132 -427
rect 8030 -461 8064 -427
rect 9962 -461 9996 -427
rect 11894 -461 11928 -427
rect 13826 -461 13860 -427
rect 15758 -461 15792 -427
rect 17690 -461 17724 -427
<< metal1 >>
rect -1171 496 -1074 592
rect 19291 496 19472 592
rect -1171 445 -1125 496
rect -1171 343 -1165 445
rect -1131 343 -1125 445
rect -241 461 -183 467
rect 290 461 348 467
rect 2222 461 2280 467
rect 4154 461 4212 467
rect 6086 461 6144 467
rect 8018 461 8076 467
rect 9950 461 10008 467
rect 11882 462 11940 468
rect 11882 461 11894 462
rect -241 427 -229 461
rect -195 427 302 461
rect 336 427 2234 461
rect 2268 427 4166 461
rect 4200 427 6098 461
rect 6132 427 8030 461
rect 8064 427 9962 461
rect 9996 428 11894 461
rect 11928 461 11940 462
rect 13814 462 13872 468
rect 13814 461 13826 462
rect 11928 428 13826 461
rect 13860 461 13872 462
rect 15746 461 15804 467
rect 17678 461 17736 467
rect 13860 428 15758 461
rect 9996 427 15758 428
rect 15792 427 17690 461
rect 17724 427 17736 461
rect -241 421 -183 427
rect 290 421 348 427
rect 2222 421 2280 427
rect 4154 421 4212 427
rect 6086 421 6144 427
rect 8018 421 8076 427
rect 9950 421 10008 427
rect 11882 422 11940 427
rect 13814 422 13872 427
rect 15746 421 15804 427
rect 17678 421 17736 427
rect -1171 331 -1125 343
rect 1754 277 1764 329
rect 1822 277 1832 329
rect 3686 277 3696 329
rect 3754 277 3764 329
rect 5618 277 5628 329
rect 5686 277 5696 329
rect 7550 277 7560 329
rect 7618 277 7628 329
rect 9482 277 9492 329
rect 9550 277 9560 329
rect 11414 277 11424 329
rect 11482 277 11492 329
rect 13346 277 13356 329
rect 13414 277 13424 329
rect 15278 277 15288 329
rect 15346 277 15356 329
rect 17210 277 17220 329
rect 17278 277 17288 329
rect 19142 277 19152 329
rect 19210 277 19220 329
rect -36 209 -26 261
rect 32 255 76 261
rect 64 221 76 255
rect 32 209 76 221
rect 1896 209 1906 261
rect 1964 255 2008 261
rect 1996 221 2008 255
rect 1964 209 2008 221
rect 3828 209 3838 261
rect 3896 255 3940 261
rect 3928 221 3940 255
rect 3896 209 3940 221
rect 5760 209 5770 261
rect 5828 255 5872 261
rect 5860 221 5872 255
rect 5828 209 5872 221
rect 7692 209 7702 261
rect 7760 255 7804 261
rect 7792 221 7804 255
rect 7760 209 7804 221
rect 9624 209 9634 261
rect 9692 255 9736 261
rect 9724 221 9736 255
rect 9692 209 9736 221
rect 11556 209 11566 261
rect 11624 255 11668 261
rect 11656 221 11668 255
rect 11624 209 11668 221
rect 13488 209 13498 261
rect 13556 255 13600 261
rect 13588 221 13600 255
rect 13556 209 13600 221
rect 15420 209 15430 261
rect 15488 255 15532 261
rect 15520 221 15532 255
rect 15488 209 15532 221
rect 17352 209 17362 261
rect 17420 255 17464 261
rect 17452 221 17464 255
rect 17420 209 17464 221
rect -1171 48 -1125 60
rect -1177 -48 -1165 48
rect -1131 -48 -1089 48
rect -1171 -60 -1125 -48
rect -36 -267 -26 -215
rect 32 -221 76 -215
rect 64 -255 76 -221
rect 32 -267 76 -255
rect 1896 -267 1906 -215
rect 1964 -221 2008 -215
rect 1996 -255 2008 -221
rect 1964 -267 2008 -255
rect 3828 -267 3838 -215
rect 3896 -221 3940 -215
rect 3928 -255 3940 -221
rect 3896 -267 3940 -255
rect 5760 -267 5770 -215
rect 5828 -221 5872 -215
rect 5860 -255 5872 -221
rect 5828 -267 5872 -255
rect 7692 -267 7702 -215
rect 7760 -221 7804 -215
rect 7792 -255 7804 -221
rect 7760 -267 7804 -255
rect 9624 -267 9634 -215
rect 9692 -221 9736 -215
rect 9724 -255 9736 -221
rect 9692 -267 9736 -255
rect 11556 -267 11566 -215
rect 11624 -221 11668 -215
rect 11656 -255 11668 -221
rect 11624 -267 11668 -255
rect 13488 -267 13498 -215
rect 13556 -221 13600 -215
rect 13588 -255 13600 -221
rect 13556 -267 13600 -255
rect 15420 -267 15430 -215
rect 15488 -221 15532 -215
rect 15520 -255 15532 -221
rect 15488 -267 15532 -255
rect 17352 -267 17362 -215
rect 17420 -221 17464 -215
rect 17452 -255 17464 -221
rect 17420 -267 17464 -255
rect -1171 -343 -1125 -331
rect 1754 -335 1764 -283
rect 1822 -335 1832 -283
rect 3686 -335 3696 -283
rect 3754 -335 3764 -283
rect 5618 -335 5628 -283
rect 5686 -335 5696 -283
rect 7550 -335 7560 -283
rect 7618 -335 7628 -283
rect 9482 -335 9492 -283
rect 9550 -335 9560 -283
rect 11414 -335 11424 -283
rect 11482 -335 11492 -283
rect 13346 -335 13356 -283
rect 13414 -335 13424 -283
rect 15278 -335 15288 -283
rect 15346 -335 15356 -283
rect 17210 -335 17220 -283
rect 17278 -335 17288 -283
rect 19142 -335 19152 -283
rect 19210 -335 19220 -283
rect -1171 -445 -1165 -343
rect -1131 -445 -1125 -343
rect -1171 -496 -1125 -445
rect -241 -427 -183 -421
rect 290 -427 348 -421
rect 2222 -427 2280 -421
rect 4154 -427 4212 -421
rect 6086 -427 6144 -421
rect 8018 -427 8076 -421
rect 9950 -427 10008 -421
rect 11882 -427 11940 -421
rect 13814 -427 13872 -421
rect 15746 -427 15804 -421
rect 17678 -427 17736 -421
rect -241 -461 -229 -427
rect -195 -461 302 -427
rect 336 -461 2234 -427
rect 2268 -461 4166 -427
rect 4200 -461 6098 -427
rect 6132 -461 8030 -427
rect 8064 -461 9962 -427
rect 9996 -461 11894 -427
rect 11928 -461 13826 -427
rect 13860 -461 15758 -427
rect 15792 -461 17690 -427
rect 17724 -461 17736 -427
rect -241 -467 -183 -461
rect 290 -467 348 -461
rect 2222 -467 2280 -461
rect 4154 -467 4212 -461
rect 6086 -467 6144 -461
rect 8018 -467 8076 -461
rect 9950 -467 10008 -461
rect 11882 -467 11940 -461
rect 13814 -467 13872 -461
rect 15746 -467 15804 -461
rect 17678 -467 17736 -461
rect 19376 -496 19472 496
rect -1171 -592 -1097 -496
rect 19291 -592 19472 -496
<< via1 >>
rect 1764 323 1822 329
rect 1764 289 1776 323
rect 1776 289 1810 323
rect 1810 289 1822 323
rect 1764 277 1822 289
rect 3696 323 3754 329
rect 3696 289 3708 323
rect 3708 289 3742 323
rect 3742 289 3754 323
rect 3696 277 3754 289
rect 5628 323 5686 329
rect 5628 289 5640 323
rect 5640 289 5674 323
rect 5674 289 5686 323
rect 5628 277 5686 289
rect 7560 323 7618 329
rect 7560 289 7572 323
rect 7572 289 7606 323
rect 7606 289 7618 323
rect 7560 277 7618 289
rect 9492 323 9550 329
rect 9492 289 9504 323
rect 9504 289 9538 323
rect 9538 289 9550 323
rect 9492 277 9550 289
rect 11424 323 11482 329
rect 11424 289 11436 323
rect 11436 289 11470 323
rect 11470 289 11482 323
rect 11424 277 11482 289
rect 13356 323 13414 329
rect 13356 289 13368 323
rect 13368 289 13402 323
rect 13402 289 13414 323
rect 13356 277 13414 289
rect 15288 323 15346 329
rect 15288 289 15300 323
rect 15300 289 15334 323
rect 15334 289 15346 323
rect 15288 277 15346 289
rect 17220 323 17278 329
rect 17220 289 17232 323
rect 17232 289 17266 323
rect 17266 289 17278 323
rect 17220 277 17278 289
rect 19152 323 19210 329
rect 19152 289 19164 323
rect 19164 289 19198 323
rect 19198 289 19210 323
rect 19152 277 19210 289
rect -26 255 32 261
rect -26 221 30 255
rect 30 221 32 255
rect -26 209 32 221
rect 1906 255 1964 261
rect 1906 221 1962 255
rect 1962 221 1964 255
rect 1906 209 1964 221
rect 3838 255 3896 261
rect 3838 221 3894 255
rect 3894 221 3896 255
rect 3838 209 3896 221
rect 5770 255 5828 261
rect 5770 221 5826 255
rect 5826 221 5828 255
rect 5770 209 5828 221
rect 7702 255 7760 261
rect 7702 221 7758 255
rect 7758 221 7760 255
rect 7702 209 7760 221
rect 9634 255 9692 261
rect 9634 221 9690 255
rect 9690 221 9692 255
rect 9634 209 9692 221
rect 11566 255 11624 261
rect 11566 221 11622 255
rect 11622 221 11624 255
rect 11566 209 11624 221
rect 13498 255 13556 261
rect 13498 221 13554 255
rect 13554 221 13556 255
rect 13498 209 13556 221
rect 15430 255 15488 261
rect 15430 221 15486 255
rect 15486 221 15488 255
rect 15430 209 15488 221
rect 17362 255 17420 261
rect 17362 221 17418 255
rect 17418 221 17420 255
rect 17362 209 17420 221
rect -26 -221 32 -215
rect -26 -255 30 -221
rect 30 -255 32 -221
rect -26 -267 32 -255
rect 1906 -221 1964 -215
rect 1906 -255 1962 -221
rect 1962 -255 1964 -221
rect 1906 -267 1964 -255
rect 3838 -221 3896 -215
rect 3838 -255 3894 -221
rect 3894 -255 3896 -221
rect 3838 -267 3896 -255
rect 5770 -221 5828 -215
rect 5770 -255 5826 -221
rect 5826 -255 5828 -221
rect 5770 -267 5828 -255
rect 7702 -221 7760 -215
rect 7702 -255 7758 -221
rect 7758 -255 7760 -221
rect 7702 -267 7760 -255
rect 9634 -221 9692 -215
rect 9634 -255 9690 -221
rect 9690 -255 9692 -221
rect 9634 -267 9692 -255
rect 11566 -221 11624 -215
rect 11566 -255 11622 -221
rect 11622 -255 11624 -221
rect 11566 -267 11624 -255
rect 13498 -221 13556 -215
rect 13498 -255 13554 -221
rect 13554 -255 13556 -221
rect 13498 -267 13556 -255
rect 15430 -221 15488 -215
rect 15430 -255 15486 -221
rect 15486 -255 15488 -221
rect 15430 -267 15488 -255
rect 17362 -221 17420 -215
rect 17362 -255 17418 -221
rect 17418 -255 17420 -221
rect 17362 -267 17420 -255
rect 1764 -289 1822 -283
rect 1764 -323 1776 -289
rect 1776 -323 1810 -289
rect 1810 -323 1822 -289
rect 1764 -335 1822 -323
rect 3696 -289 3754 -283
rect 3696 -323 3708 -289
rect 3708 -323 3742 -289
rect 3742 -323 3754 -289
rect 3696 -335 3754 -323
rect 5628 -289 5686 -283
rect 5628 -323 5640 -289
rect 5640 -323 5674 -289
rect 5674 -323 5686 -289
rect 5628 -335 5686 -323
rect 7560 -289 7618 -283
rect 7560 -323 7572 -289
rect 7572 -323 7606 -289
rect 7606 -323 7618 -289
rect 7560 -335 7618 -323
rect 9492 -289 9550 -283
rect 9492 -323 9504 -289
rect 9504 -323 9538 -289
rect 9538 -323 9550 -289
rect 9492 -335 9550 -323
rect 11424 -289 11482 -283
rect 11424 -323 11436 -289
rect 11436 -323 11470 -289
rect 11470 -323 11482 -289
rect 11424 -335 11482 -323
rect 13356 -289 13414 -283
rect 13356 -323 13368 -289
rect 13368 -323 13402 -289
rect 13402 -323 13414 -289
rect 13356 -335 13414 -323
rect 15288 -289 15346 -283
rect 15288 -323 15300 -289
rect 15300 -323 15334 -289
rect 15334 -323 15346 -289
rect 15288 -335 15346 -323
rect 17220 -289 17278 -283
rect 17220 -323 17232 -289
rect 17232 -323 17266 -289
rect 17266 -323 17278 -289
rect 17220 -335 17278 -323
rect 19152 -289 19210 -283
rect 19152 -323 19164 -289
rect 19164 -323 19198 -289
rect 19198 -323 19210 -289
rect 19152 -335 19210 -323
<< metal2 >>
rect 1764 329 1822 718
rect -26 261 32 271
rect 1764 267 1822 277
rect 3696 329 3754 718
rect -26 -215 32 209
rect -26 -656 32 -267
rect 1906 261 1964 271
rect 3696 267 3754 277
rect 5628 329 5686 718
rect 1906 -215 1964 209
rect 1764 -283 1822 -273
rect 1764 -724 1822 -335
rect 1906 -656 1964 -267
rect 3838 261 3896 271
rect 5628 267 5686 277
rect 7560 329 7618 718
rect 3838 -215 3896 209
rect 3696 -283 3754 -273
rect 3696 -724 3754 -335
rect 3838 -656 3896 -267
rect 5770 261 5828 271
rect 7560 267 7618 277
rect 9492 329 9550 718
rect 5770 -215 5828 209
rect 5628 -283 5686 -273
rect 5628 -724 5686 -335
rect 5770 -656 5828 -267
rect 7702 261 7760 271
rect 9492 267 9550 277
rect 11424 329 11482 718
rect 7702 -215 7760 209
rect 7560 -283 7618 -273
rect 7560 -724 7618 -335
rect 7702 -656 7760 -267
rect 9634 261 9692 271
rect 11424 267 11482 277
rect 13356 329 13414 718
rect 9634 -215 9692 209
rect 9492 -283 9550 -273
rect 9492 -724 9550 -335
rect 9634 -656 9692 -267
rect 11566 261 11624 271
rect 13356 267 13414 277
rect 15288 329 15346 718
rect 11566 -215 11624 209
rect 11424 -283 11482 -273
rect 11424 -724 11482 -335
rect 11566 -656 11624 -267
rect 13498 261 13556 271
rect 15288 267 15346 277
rect 17220 329 17278 718
rect 13498 -215 13556 209
rect 13356 -283 13414 -273
rect 13356 -724 13414 -335
rect 13498 -656 13556 -267
rect 15430 261 15488 271
rect 17220 267 17278 277
rect 19152 329 19210 718
rect 15430 -215 15488 209
rect 15288 -283 15346 -273
rect 15288 -724 15346 -335
rect 15430 -656 15488 -267
rect 17362 261 17420 271
rect 19152 267 19210 277
rect 17362 -215 17420 209
rect 17220 -283 17278 -273
rect 17220 -723 17278 -335
rect 17362 -656 17420 -267
rect 19152 -283 19210 -273
rect 19152 -724 19210 -335
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform 1 0 1932 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_1
timestamp 1730246015
transform 1 0 0 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_2
timestamp 1730246015
transform 1 0 5796 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_3
timestamp 1730246015
transform 1 0 3864 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_4
timestamp 1730246015
transform 1 0 9660 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_5
timestamp 1730246015
transform 1 0 7728 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_6
timestamp 1730246015
transform 1 0 13524 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_7
timestamp 1730246015
transform 1 0 11592 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_8
timestamp 1730246015
transform 1 0 17388 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sky130_fd_sc_hd__dfrtp_2_9
timestamp 1730246015
transform 1 0 15456 0 -1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1[1]
timestamp 1730246015
transform 1 0 1932 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1[2]
timestamp 1730246015
transform 1 0 3864 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1[3]
timestamp 1730246015
transform 1 0 5796 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1[4]
timestamp 1730246015
transform 1 0 7728 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1[5]
timestamp 1730246015
transform 1 0 9660 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1[6]
timestamp 1730246015
transform 1 0 11592 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1[7]
timestamp 1730246015
transform 1 0 13524 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1[8]
timestamp 1730246015
transform 1 0 15456 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1[9]
timestamp 1730246015
transform 1 0 17388 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_8  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform 1 0 -1104 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  x1[0]
timestamp 1730246015
transform 1 0 0 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_8  x2
timestamp 1730246015
transform 1 0 -1104 0 -1 0
box -38 -48 1142 592
<< end >>
