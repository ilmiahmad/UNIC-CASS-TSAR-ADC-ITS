magic
tech sky130A
magscale 1 2
timestamp 1730995243
<< dnwell >>
rect -8 -2 67002 60777
<< metal1 >>
rect 32790 40494 32800 40975
rect 32984 40974 32994 40975
rect 34000 40974 34010 40976
rect 32984 40495 34010 40974
rect 34194 40495 34204 40976
rect 32984 40494 34194 40495
rect 33002 39775 33012 40256
rect 33196 39775 33798 40256
rect 33982 39775 33992 40256
rect 33214 39054 33224 39535
rect 33408 39054 33586 39535
rect 33770 39054 33780 39535
rect 33215 21241 33225 21722
rect 33409 21721 33419 21722
rect 33409 21241 33586 21721
rect 33576 21240 33586 21241
rect 33770 21240 33780 21721
rect 33002 20521 33012 21002
rect 33196 21001 33206 21002
rect 33196 20521 33798 21001
rect 33788 20520 33798 20521
rect 33982 20520 33992 21001
rect 32790 19801 32800 20282
rect 32984 20281 32994 20282
rect 32984 19801 34010 20281
rect 34000 19800 34010 19801
rect 34194 19800 34204 20281
<< via1 >>
rect 32800 40494 32984 40975
rect 34010 40495 34194 40976
rect 33012 39775 33196 40256
rect 33798 39775 33982 40256
rect 33224 39054 33408 39535
rect 33586 39054 33770 39535
rect 33225 21241 33409 21722
rect 33586 21240 33770 21721
rect 33012 20521 33196 21002
rect 33798 20520 33982 21001
rect 32800 19801 32984 20282
rect 34010 19800 34194 20281
<< metal2 >>
rect 32800 40975 32984 40985
rect 32800 40484 32984 40494
rect 34010 40976 34194 40986
rect 34010 40485 34194 40495
rect 33012 40256 33196 40266
rect 33012 39765 33196 39775
rect 33798 40256 33982 40266
rect 33798 39765 33982 39775
rect 33224 39535 33408 39545
rect 33224 39044 33408 39054
rect 33586 39535 33770 39545
rect 33586 39044 33770 39054
rect -8 37251 176 37663
rect 204 37228 388 37656
rect 416 37208 600 37637
rect 33225 21722 33409 21732
rect 33225 21231 33409 21241
rect 33586 21721 33770 21731
rect 33586 21230 33770 21240
rect 33012 21002 33196 21012
rect 33012 20511 33196 20521
rect 33798 21001 33982 21011
rect 33798 20510 33982 20520
rect 32800 20282 32984 20292
rect 32800 19791 32984 19801
rect 34010 20281 34194 20291
rect 34010 19790 34194 19800
<< metal3 >>
rect -2 36677 180 36773
rect 33312 36677 33738 36773
rect 5 36521 199 36617
rect 33312 36521 33692 36617
rect -5 36365 190 36461
rect 33306 36365 33684 36461
rect -8 36209 195 36305
rect 33262 36209 33698 36305
rect -8 36053 195 36149
rect 33281 36053 33685 36149
rect 3 35897 187 35993
rect 33293 35897 33692 35993
rect -8 35741 195 35837
rect 33305 35741 33693 35837
rect 11 35585 214 35681
rect 33256 35585 33713 35681
rect -8 35429 212 35525
rect 33267 35429 33726 35525
rect -8 35273 243 35369
rect 33279 35273 33696 35369
rect -8 31042 198 31138
rect 33311 31042 33728 31138
rect -8 30886 222 30982
rect 33277 30886 33755 30982
rect -7 30730 225 30826
rect 33271 30730 33752 30826
rect -8 30574 228 30670
rect 33259 30574 33728 30670
rect -8 30418 228 30514
rect 33269 30418 33753 30514
rect -8 30262 230 30358
rect 33261 30262 33742 30358
rect -8 30106 230 30202
rect 33244 30106 33732 30202
rect -3 29950 228 30046
rect 33250 29950 33735 30046
rect -8 29794 230 29890
rect 33246 29794 33739 29890
rect -7 29638 244 29734
rect 33265 29638 33719 29734
rect -8 25407 223 25503
rect 33298 25407 33690 25503
rect -8 25251 247 25347
rect 33312 25251 33705 25347
rect -8 25095 271 25191
rect 33269 25095 33698 25191
rect 0 24939 262 25035
rect 33277 24939 33703 25035
rect -8 24783 268 24879
rect 33255 24783 33705 24879
rect -7 24627 262 24723
rect 33285 24627 33701 24723
rect -5 24471 249 24567
rect 33259 24471 33698 24567
rect -8 24315 271 24411
rect 33285 24315 33707 24411
rect -8 24159 270 24255
rect 33267 24159 33705 24255
rect 8 24003 279 24099
rect 33245 24003 33711 24099
<< metal4 >>
rect 980 60673 65652 60777
rect 1094 -1 66098 103
use single_10b_cdac  single_10b_cdac_0
timestamp 1730971434
transform 1 0 -69036 0 1 40901
box 102622 -40903 136038 19876
use single_10b_cdac  single_10b_cdac_1
timestamp 1730971434
transform 1 0 -102630 0 1 40901
box 102622 -40903 136038 19876
<< labels >>
flabel metal2 44 37567 104 37632 0 FreeSans 800 0 0 0 VCM
port 0 nsew
flabel metal2 257 37436 317 37501 0 FreeSans 800 0 0 0 VSREF
port 1 nsew
flabel metal2 467 37279 527 37344 0 FreeSans 800 0 0 0 VDREF
port 2 nsew
flabel metal3 34 36705 59 36749 0 FreeSans 800 0 0 0 SWP_IN[0]
port 3 nsew
flabel metal3 33 36549 58 36593 0 FreeSans 800 0 0 0 SWP_IN[1]
port 4 nsew
flabel metal3 40 36387 65 36431 0 FreeSans 800 0 0 0 SWP_IN[2]
port 5 nsew
flabel metal3 35 36242 60 36286 0 FreeSans 800 0 0 0 SWP_IN[3]
port 6 nsew
flabel metal3 37 36085 62 36129 0 FreeSans 800 0 0 0 SWP_IN[4]
port 7 nsew
flabel metal3 47 35916 72 35960 0 FreeSans 800 0 0 0 SWP_IN[5]
port 8 nsew
flabel metal3 37 35770 62 35814 0 FreeSans 800 0 0 0 SWP_IN[6]
port 9 nsew
flabel metal3 45 35619 70 35663 0 FreeSans 800 0 0 0 SWP_IN[7]
port 10 nsew
flabel metal3 36 35450 61 35494 0 FreeSans 800 0 0 0 SWP_IN[8]
port 11 nsew
flabel metal3 35 35303 60 35347 0 FreeSans 800 0 0 0 SWP_IN[9]
port 12 nsew
flabel metal3 26 31073 51 31117 0 FreeSans 800 0 0 0 CF[9]
port 13 nsew
flabel metal3 31 30911 56 30955 0 FreeSans 800 0 0 0 CF[8]
port 14 nsew
flabel metal3 52 30759 77 30803 0 FreeSans 800 0 0 0 CF[7]
port 15 nsew
flabel metal3 47 30610 72 30654 0 FreeSans 800 0 0 0 CF[6]
port 16 nsew
flabel metal3 42 30455 67 30499 0 FreeSans 800 0 0 0 CF[5]
port 17 nsew
flabel metal3 54 30293 79 30337 0 FreeSans 800 0 0 0 CF[4]
port 18 nsew
flabel metal3 51 30136 76 30180 0 FreeSans 800 0 0 0 CF[3]
port 19 nsew
flabel metal3 46 29981 71 30025 0 FreeSans 800 0 0 0 CF[2]
port 20 nsew
flabel metal3 52 29828 77 29872 0 FreeSans 800 0 0 0 CF[1]
port 21 nsew
flabel metal3 47 29672 72 29716 0 FreeSans 800 0 0 0 CF[0]
port 22 nsew
flabel metal3 24 25430 49 25474 0 FreeSans 800 0 0 0 SWN_IN[9]
port 23 nsew
flabel metal3 34 25293 59 25337 0 FreeSans 800 0 0 0 SWN_IN[8]
port 24 nsew
flabel metal3 25 25114 50 25158 0 FreeSans 800 0 0 0 SWN_IN[7]
port 25 nsew
flabel metal3 20 24974 45 25018 0 FreeSans 800 0 0 0 SWN_IN[6]
port 26 nsew
flabel metal3 30 24805 55 24849 0 FreeSans 800 0 0 0 SWN_IN[5]
port 27 nsew
flabel metal3 29 24652 54 24696 0 FreeSans 800 0 0 0 SWN_IN[4]
port 28 nsew
flabel metal3 30 24500 55 24544 0 FreeSans 800 0 0 0 SWN_IN[3]
port 29 nsew
flabel metal3 22 24340 47 24384 0 FreeSans 800 0 0 0 SWN_IN[2]
port 30 nsew
flabel metal3 30 24182 55 24226 0 FreeSans 800 0 0 0 SWN_IN[1]
port 31 nsew
flabel metal3 37 24027 62 24071 0 FreeSans 800 0 0 0 SWN_IN[0]
port 32 nsew
flabel metal4 32479 60688 32581 60751 0 FreeSans 800 0 0 0 VCP
port 33 nsew
flabel metal4 34363 27 34437 71 0 FreeSans 800 0 0 0 VCN
port 34 nsew
<< end >>
