magic
tech sky130A
magscale 1 2
timestamp 1730868737
use cdac_10b  cdac_10b_0
timestamp 1730868527
transform 1 0 -18 0 1 30
box -8 -2 67002 60777
use sh_bsw4  sh_bsw4_0
timestamp 1730800698
transform 1 0 67227 0 1 26250
box -23 -164 5575 3264
use tdc  tdc_0
timestamp 1730868527
transform 1 0 -31840 0 1 13821
box -4836 -3709 9311 2246
<< end >>
