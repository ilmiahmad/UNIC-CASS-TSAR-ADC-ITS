magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect 278 -2147 312 -2071
rect 278 -2237 312 -2231
rect 664 -2147 698 -2071
rect 664 -2237 698 -2231
rect 1050 -2147 1084 -2071
rect 1050 -2237 1084 -2231
rect 1156 -2271 1190 -2071
rect 1156 -2361 1190 -2355
rect 1542 -2271 1576 -2071
rect 1542 -2361 1576 -2355
rect 1928 -2271 1962 -2071
rect 1928 -2361 1962 -2355
<< viali >>
rect 278 -2231 312 -2147
rect 664 -2231 698 -2147
rect 1050 -2231 1084 -2147
rect 1156 -2355 1190 -2271
rect 1542 -2355 1576 -2271
rect 1928 -2355 1962 -2271
<< metal1 >>
rect 442 2168 462 2220
rect 514 2168 534 2220
rect 828 2168 848 2220
rect 900 2168 920 2220
rect 372 2078 378 2130
rect 430 2078 436 2130
rect 372 2006 436 2078
rect 372 1954 378 2006
rect 430 1954 436 2006
rect 372 1882 436 1954
rect 372 1830 378 1882
rect 430 1830 436 1882
rect 540 2078 546 2130
rect 598 2078 764 2130
rect 816 2078 822 2130
rect 540 2006 822 2078
rect 540 1954 546 2006
rect 598 1954 764 2006
rect 816 1954 822 2006
rect 540 1882 822 1954
rect 540 1830 546 1882
rect 598 1830 764 1882
rect 816 1830 822 1882
rect 926 2078 932 2130
rect 984 2078 990 2130
rect 926 2006 990 2078
rect 926 1954 932 2006
rect 984 1954 990 2006
rect 926 1882 990 1954
rect 926 1830 932 1882
rect 984 1830 990 1882
rect 442 1740 462 1792
rect 514 1740 534 1792
rect 828 1740 848 1792
rect 900 1740 920 1792
rect 442 1632 462 1684
rect 514 1632 534 1684
rect 828 1632 848 1684
rect 900 1632 920 1684
rect 372 1542 378 1594
rect 430 1542 436 1594
rect 372 1470 436 1542
rect 372 1418 378 1470
rect 430 1418 436 1470
rect 372 1346 436 1418
rect 372 1294 378 1346
rect 430 1294 436 1346
rect 540 1542 546 1594
rect 598 1542 764 1594
rect 816 1542 822 1594
rect 540 1470 822 1542
rect 540 1418 546 1470
rect 598 1418 764 1470
rect 816 1418 822 1470
rect 540 1346 822 1418
rect 540 1294 546 1346
rect 598 1294 764 1346
rect 816 1294 822 1346
rect 926 1542 932 1594
rect 984 1542 990 1594
rect 926 1470 990 1542
rect 926 1418 932 1470
rect 984 1418 990 1470
rect 926 1346 990 1418
rect 926 1294 932 1346
rect 984 1294 990 1346
rect 442 1204 462 1256
rect 514 1204 534 1256
rect 828 1204 848 1256
rect 900 1204 920 1256
rect 442 1096 462 1148
rect 514 1096 534 1148
rect 828 1096 848 1148
rect 900 1096 920 1148
rect 372 1006 378 1058
rect 430 1006 436 1058
rect 372 934 436 1006
rect 372 882 378 934
rect 430 882 436 934
rect 372 810 436 882
rect 372 758 378 810
rect 430 758 436 810
rect 540 1006 546 1058
rect 598 1006 764 1058
rect 816 1006 822 1058
rect 540 934 822 1006
rect 540 882 546 934
rect 598 882 764 934
rect 816 882 822 934
rect 540 810 822 882
rect 540 758 546 810
rect 598 758 764 810
rect 816 758 822 810
rect 926 1006 932 1058
rect 984 1006 990 1058
rect 926 934 990 1006
rect 926 882 932 934
rect 984 882 990 934
rect 926 810 990 882
rect 926 758 932 810
rect 984 758 990 810
rect 442 668 462 720
rect 514 668 534 720
rect 828 668 848 720
rect 900 668 920 720
rect 442 560 462 612
rect 514 560 534 612
rect 828 560 848 612
rect 900 560 920 612
rect 372 470 378 522
rect 430 470 436 522
rect 372 398 436 470
rect 372 346 378 398
rect 430 346 436 398
rect 372 274 436 346
rect 372 222 378 274
rect 430 222 436 274
rect 540 470 546 522
rect 598 470 764 522
rect 816 470 822 522
rect 540 398 822 470
rect 540 346 546 398
rect 598 346 764 398
rect 816 346 822 398
rect 540 274 822 346
rect 540 222 546 274
rect 598 222 764 274
rect 816 222 822 274
rect 926 470 932 522
rect 984 470 990 522
rect 926 398 990 470
rect 1320 424 1340 476
rect 1392 424 1412 476
rect 1706 424 1726 476
rect 1778 424 1798 476
rect 926 346 932 398
rect 984 395 990 398
rect 984 347 1314 395
rect 984 346 1256 347
rect 926 295 1256 346
rect 1308 295 1314 347
rect 1418 347 1700 395
rect 1418 295 1424 347
rect 1476 295 1642 347
rect 1694 295 1700 347
rect 1804 347 1868 395
rect 1804 295 1810 347
rect 1862 295 1868 347
rect 926 274 990 295
rect 926 222 932 274
rect 984 222 990 274
rect 1320 214 1340 266
rect 1392 214 1412 266
rect 1706 214 1726 266
rect 1778 214 1798 266
rect 442 132 462 184
rect 514 132 534 184
rect 828 132 848 184
rect 900 132 920 184
rect 1320 106 1340 158
rect 1392 106 1412 158
rect 1706 106 1726 158
rect 1778 106 1798 158
rect 442 24 462 76
rect 514 24 534 76
rect 828 24 848 76
rect 900 24 920 76
rect 1250 29 1314 77
rect 372 -66 378 -14
rect 430 -66 436 -14
rect 372 -138 436 -66
rect 372 -190 378 -138
rect 430 -190 436 -138
rect 372 -262 436 -190
rect 372 -314 378 -262
rect 430 -314 436 -262
rect 540 -66 546 -14
rect 598 -66 764 -14
rect 816 -66 822 -14
rect 540 -138 822 -66
rect 540 -190 546 -138
rect 598 -190 764 -138
rect 816 -190 822 -138
rect 540 -262 822 -190
rect 540 -314 546 -262
rect 598 -314 764 -262
rect 816 -314 822 -262
rect 926 -66 932 -14
rect 984 -66 990 -14
rect 1250 -23 1256 29
rect 1308 -23 1314 29
rect 1418 29 1700 77
rect 1418 -23 1424 29
rect 1476 -23 1642 29
rect 1694 -23 1700 29
rect 1804 29 1868 77
rect 1804 -23 1810 29
rect 1862 -23 1868 29
rect 926 -138 990 -66
rect 1320 -104 1340 -52
rect 1392 -104 1412 -52
rect 1706 -104 1726 -52
rect 1778 -104 1798 -52
rect 926 -190 932 -138
rect 984 -190 990 -138
rect 926 -262 990 -190
rect 1321 -212 1340 -160
rect 1392 -212 1413 -160
rect 1706 -212 1726 -160
rect 1778 -212 1798 -160
rect 926 -314 932 -262
rect 984 -314 990 -262
rect 1250 -289 1314 -241
rect 1250 -341 1256 -289
rect 1308 -341 1314 -289
rect 1418 -289 1700 -241
rect 1418 -341 1424 -289
rect 1476 -341 1642 -289
rect 1694 -341 1700 -289
rect 1804 -289 1868 -241
rect 1804 -341 1810 -289
rect 1862 -341 1868 -289
rect 442 -404 462 -352
rect 514 -404 534 -352
rect 828 -404 848 -352
rect 900 -404 920 -352
rect 1320 -422 1340 -370
rect 1392 -422 1412 -370
rect 1706 -422 1726 -370
rect 1778 -422 1798 -370
rect 442 -512 462 -460
rect 514 -512 534 -460
rect 828 -512 848 -460
rect 900 -512 920 -460
rect 1320 -530 1340 -478
rect 1392 -530 1412 -478
rect 1705 -530 1726 -478
rect 1778 -530 1797 -478
rect 372 -602 378 -550
rect 430 -602 436 -550
rect 372 -674 436 -602
rect 372 -726 378 -674
rect 430 -726 436 -674
rect 372 -798 436 -726
rect 372 -850 378 -798
rect 430 -850 436 -798
rect 540 -602 546 -550
rect 598 -602 764 -550
rect 816 -602 822 -550
rect 540 -674 822 -602
rect 540 -726 546 -674
rect 598 -726 764 -674
rect 816 -726 822 -674
rect 540 -798 822 -726
rect 540 -850 546 -798
rect 598 -850 764 -798
rect 816 -850 822 -798
rect 926 -602 932 -550
rect 984 -559 990 -550
rect 984 -602 1314 -559
rect 926 -607 1314 -602
rect 926 -659 1256 -607
rect 1308 -659 1314 -607
rect 1418 -607 1700 -559
rect 1418 -659 1424 -607
rect 1476 -659 1642 -607
rect 1694 -659 1700 -607
rect 1804 -607 1868 -559
rect 1804 -659 1810 -607
rect 1862 -659 1868 -607
rect 926 -674 990 -659
rect 926 -726 932 -674
rect 984 -726 990 -674
rect 926 -798 990 -726
rect 1320 -740 1340 -688
rect 1392 -740 1412 -688
rect 1706 -740 1726 -688
rect 1778 -740 1798 -688
rect 926 -850 932 -798
rect 984 -850 990 -798
rect 1320 -848 1340 -796
rect 1392 -848 1412 -796
rect 1706 -848 1726 -796
rect 1778 -848 1798 -796
rect 442 -940 462 -888
rect 514 -940 534 -888
rect 828 -940 848 -888
rect 900 -940 920 -888
rect 1250 -925 1314 -877
rect 1250 -977 1256 -925
rect 1308 -977 1314 -925
rect 1418 -925 1700 -877
rect 1418 -977 1424 -925
rect 1476 -977 1642 -925
rect 1694 -977 1700 -925
rect 1804 -925 1868 -877
rect 1804 -977 1810 -925
rect 1862 -977 1868 -925
rect 442 -1048 462 -996
rect 514 -1048 534 -996
rect 828 -1048 848 -996
rect 900 -1048 920 -996
rect 1320 -1058 1340 -1006
rect 1392 -1058 1412 -1006
rect 1706 -1058 1726 -1006
rect 1778 -1058 1798 -1006
rect 372 -1138 378 -1086
rect 430 -1138 436 -1086
rect 372 -1210 436 -1138
rect 372 -1262 378 -1210
rect 430 -1262 436 -1210
rect 372 -1334 436 -1262
rect 372 -1386 378 -1334
rect 430 -1386 436 -1334
rect 540 -1138 546 -1086
rect 598 -1138 764 -1086
rect 816 -1138 822 -1086
rect 540 -1210 822 -1138
rect 540 -1262 546 -1210
rect 598 -1262 764 -1210
rect 816 -1262 822 -1210
rect 540 -1334 822 -1262
rect 540 -1386 546 -1334
rect 598 -1386 764 -1334
rect 816 -1386 822 -1334
rect 926 -1138 932 -1086
rect 984 -1138 990 -1086
rect 926 -1195 990 -1138
rect 1320 -1166 1340 -1114
rect 1392 -1166 1412 -1114
rect 1706 -1166 1726 -1114
rect 1778 -1166 1798 -1114
rect 926 -1210 1314 -1195
rect 926 -1262 932 -1210
rect 984 -1243 1314 -1210
rect 984 -1262 1256 -1243
rect 926 -1295 1256 -1262
rect 1308 -1295 1314 -1243
rect 1418 -1243 1700 -1195
rect 1418 -1295 1424 -1243
rect 1476 -1295 1642 -1243
rect 1694 -1295 1700 -1243
rect 1804 -1243 1868 -1195
rect 1804 -1295 1810 -1243
rect 1862 -1295 1868 -1243
rect 926 -1334 990 -1295
rect 926 -1386 932 -1334
rect 984 -1386 990 -1334
rect 1320 -1376 1340 -1324
rect 1392 -1376 1412 -1324
rect 1706 -1376 1726 -1324
rect 1778 -1376 1798 -1324
rect 442 -1476 462 -1424
rect 514 -1476 534 -1424
rect 828 -1476 848 -1424
rect 900 -1476 920 -1424
rect 1321 -1484 1340 -1432
rect 1392 -1484 1413 -1432
rect 1706 -1484 1726 -1432
rect 1778 -1484 1798 -1432
rect 442 -1584 462 -1532
rect 514 -1584 534 -1532
rect 828 -1584 848 -1532
rect 900 -1584 920 -1532
rect 1250 -1561 1314 -1513
rect 1250 -1613 1256 -1561
rect 1308 -1613 1314 -1561
rect 1418 -1561 1700 -1513
rect 1418 -1613 1424 -1561
rect 1476 -1613 1642 -1561
rect 1694 -1613 1700 -1561
rect 1804 -1561 1868 -1513
rect 1804 -1613 1810 -1561
rect 1862 -1613 1868 -1561
rect 372 -1674 378 -1622
rect 430 -1674 436 -1622
rect 372 -1746 436 -1674
rect 372 -1798 378 -1746
rect 430 -1798 436 -1746
rect 372 -1870 436 -1798
rect 372 -1922 378 -1870
rect 430 -1922 436 -1870
rect 540 -1674 546 -1622
rect 598 -1674 764 -1622
rect 816 -1674 822 -1622
rect 540 -1746 822 -1674
rect 540 -1798 546 -1746
rect 598 -1798 764 -1746
rect 816 -1798 822 -1746
rect 540 -1870 822 -1798
rect 540 -1922 546 -1870
rect 598 -1922 764 -1870
rect 816 -1922 822 -1870
rect 926 -1674 932 -1622
rect 984 -1674 990 -1622
rect 926 -1746 990 -1674
rect 1320 -1694 1340 -1642
rect 1392 -1694 1412 -1642
rect 1706 -1694 1726 -1642
rect 1778 -1694 1798 -1642
rect 926 -1798 932 -1746
rect 984 -1798 990 -1746
rect 926 -1831 990 -1798
rect 1320 -1802 1340 -1750
rect 1392 -1802 1412 -1750
rect 1705 -1802 1726 -1750
rect 1778 -1802 1797 -1750
rect 926 -1870 1314 -1831
rect 926 -1922 932 -1870
rect 984 -1879 1314 -1870
rect 984 -1922 1256 -1879
rect 926 -1931 1256 -1922
rect 1308 -1931 1314 -1879
rect 1418 -1879 1700 -1831
rect 1418 -1931 1424 -1879
rect 1476 -1931 1642 -1879
rect 1694 -1931 1700 -1879
rect 1804 -1879 1868 -1831
rect 1804 -1931 1810 -1879
rect 1862 -1931 1868 -1879
rect 442 -2012 462 -1960
rect 514 -2012 534 -1960
rect 828 -2012 848 -1960
rect 900 -2012 920 -1960
rect 1320 -2012 1340 -1960
rect 1392 -2012 1412 -1960
rect 1706 -2012 1726 -1960
rect 1778 -2012 1798 -1960
rect 456 -2092 462 -2040
rect 514 -2092 1726 -2040
rect 1778 -2092 1784 -2040
rect 242 -2147 378 -2141
rect 242 -2231 278 -2147
rect 312 -2231 378 -2147
rect 430 -2147 1998 -2141
rect 430 -2231 664 -2147
rect 698 -2231 1050 -2147
rect 1084 -2231 1998 -2147
rect 242 -2237 1998 -2231
rect 242 -2271 1810 -2265
rect 242 -2355 1156 -2271
rect 1190 -2355 1542 -2271
rect 1576 -2355 1810 -2271
rect 1862 -2271 1998 -2265
rect 1862 -2355 1928 -2271
rect 1962 -2355 1998 -2271
rect 242 -2361 1998 -2355
<< via1 >>
rect 462 2168 514 2220
rect 848 2168 900 2220
rect 378 2078 430 2130
rect 378 1954 430 2006
rect 378 1830 430 1882
rect 546 2078 598 2130
rect 764 2078 816 2130
rect 546 1954 598 2006
rect 764 1954 816 2006
rect 546 1830 598 1882
rect 764 1830 816 1882
rect 932 2078 984 2130
rect 932 1954 984 2006
rect 932 1830 984 1882
rect 462 1740 514 1792
rect 848 1740 900 1792
rect 462 1632 514 1684
rect 848 1632 900 1684
rect 378 1542 430 1594
rect 378 1418 430 1470
rect 378 1294 430 1346
rect 546 1542 598 1594
rect 764 1542 816 1594
rect 546 1418 598 1470
rect 764 1418 816 1470
rect 546 1294 598 1346
rect 764 1294 816 1346
rect 932 1542 984 1594
rect 932 1418 984 1470
rect 932 1294 984 1346
rect 462 1204 514 1256
rect 848 1204 900 1256
rect 462 1096 514 1148
rect 848 1096 900 1148
rect 378 1006 430 1058
rect 378 882 430 934
rect 378 758 430 810
rect 546 1006 598 1058
rect 764 1006 816 1058
rect 546 882 598 934
rect 764 882 816 934
rect 546 758 598 810
rect 764 758 816 810
rect 932 1006 984 1058
rect 932 882 984 934
rect 932 758 984 810
rect 462 668 514 720
rect 848 668 900 720
rect 462 560 514 612
rect 848 560 900 612
rect 378 470 430 522
rect 378 346 430 398
rect 378 222 430 274
rect 546 470 598 522
rect 764 470 816 522
rect 546 346 598 398
rect 764 346 816 398
rect 546 222 598 274
rect 764 222 816 274
rect 932 470 984 522
rect 1340 424 1392 476
rect 1726 424 1778 476
rect 932 346 984 398
rect 1256 295 1308 347
rect 1424 295 1476 347
rect 1642 295 1694 347
rect 1810 295 1862 347
rect 932 222 984 274
rect 1340 214 1392 266
rect 1726 214 1778 266
rect 462 132 514 184
rect 848 132 900 184
rect 1340 106 1392 158
rect 1726 106 1778 158
rect 462 24 514 76
rect 848 24 900 76
rect 378 -66 430 -14
rect 378 -190 430 -138
rect 378 -314 430 -262
rect 546 -66 598 -14
rect 764 -66 816 -14
rect 546 -190 598 -138
rect 764 -190 816 -138
rect 546 -314 598 -262
rect 764 -314 816 -262
rect 932 -66 984 -14
rect 1256 -23 1308 29
rect 1424 -23 1476 29
rect 1642 -23 1694 29
rect 1810 -23 1862 29
rect 1340 -104 1392 -52
rect 1726 -104 1778 -52
rect 932 -190 984 -138
rect 1340 -212 1392 -160
rect 1726 -212 1778 -160
rect 932 -314 984 -262
rect 1256 -341 1308 -289
rect 1424 -341 1476 -289
rect 1642 -341 1694 -289
rect 1810 -341 1862 -289
rect 462 -404 514 -352
rect 848 -404 900 -352
rect 1340 -422 1392 -370
rect 1726 -422 1778 -370
rect 462 -512 514 -460
rect 848 -512 900 -460
rect 1340 -530 1392 -478
rect 1726 -530 1778 -478
rect 378 -602 430 -550
rect 378 -726 430 -674
rect 378 -850 430 -798
rect 546 -602 598 -550
rect 764 -602 816 -550
rect 546 -726 598 -674
rect 764 -726 816 -674
rect 546 -850 598 -798
rect 764 -850 816 -798
rect 932 -602 984 -550
rect 1256 -659 1308 -607
rect 1424 -659 1476 -607
rect 1642 -659 1694 -607
rect 1810 -659 1862 -607
rect 932 -726 984 -674
rect 1340 -740 1392 -688
rect 1726 -740 1778 -688
rect 932 -850 984 -798
rect 1340 -848 1392 -796
rect 1726 -848 1778 -796
rect 462 -940 514 -888
rect 848 -940 900 -888
rect 1256 -977 1308 -925
rect 1424 -977 1476 -925
rect 1642 -977 1694 -925
rect 1810 -977 1862 -925
rect 462 -1048 514 -996
rect 848 -1048 900 -996
rect 1340 -1058 1392 -1006
rect 1726 -1058 1778 -1006
rect 378 -1138 430 -1086
rect 378 -1262 430 -1210
rect 378 -1386 430 -1334
rect 546 -1138 598 -1086
rect 764 -1138 816 -1086
rect 546 -1262 598 -1210
rect 764 -1262 816 -1210
rect 546 -1386 598 -1334
rect 764 -1386 816 -1334
rect 932 -1138 984 -1086
rect 1340 -1166 1392 -1114
rect 1726 -1166 1778 -1114
rect 932 -1262 984 -1210
rect 1256 -1295 1308 -1243
rect 1424 -1295 1476 -1243
rect 1642 -1295 1694 -1243
rect 1810 -1295 1862 -1243
rect 932 -1386 984 -1334
rect 1340 -1376 1392 -1324
rect 1726 -1376 1778 -1324
rect 462 -1476 514 -1424
rect 848 -1476 900 -1424
rect 1340 -1484 1392 -1432
rect 1726 -1484 1778 -1432
rect 462 -1584 514 -1532
rect 848 -1584 900 -1532
rect 1256 -1613 1308 -1561
rect 1424 -1613 1476 -1561
rect 1642 -1613 1694 -1561
rect 1810 -1613 1862 -1561
rect 378 -1674 430 -1622
rect 378 -1798 430 -1746
rect 378 -1922 430 -1870
rect 546 -1674 598 -1622
rect 764 -1674 816 -1622
rect 546 -1798 598 -1746
rect 764 -1798 816 -1746
rect 546 -1922 598 -1870
rect 764 -1922 816 -1870
rect 932 -1674 984 -1622
rect 1340 -1694 1392 -1642
rect 1726 -1694 1778 -1642
rect 932 -1798 984 -1746
rect 1340 -1802 1392 -1750
rect 1726 -1802 1778 -1750
rect 932 -1922 984 -1870
rect 1256 -1931 1308 -1879
rect 1424 -1931 1476 -1879
rect 1642 -1931 1694 -1879
rect 1810 -1931 1862 -1879
rect 462 -2012 514 -1960
rect 848 -2012 900 -1960
rect 1340 -2012 1392 -1960
rect 1726 -2012 1778 -1960
rect 462 -2092 514 -2040
rect 1726 -2092 1778 -2040
rect 378 -2231 430 -2141
rect 1810 -2355 1862 -2265
<< metal2 >>
rect 460 2220 516 2226
rect 460 2168 462 2220
rect 514 2168 516 2220
rect 376 2130 432 2136
rect 376 2078 378 2130
rect 430 2078 432 2130
rect 376 2006 432 2078
rect 376 1954 378 2006
rect 430 1954 432 2006
rect 376 1882 432 1954
rect 376 1830 378 1882
rect 430 1830 432 1882
rect 376 1594 432 1830
rect 376 1542 378 1594
rect 430 1542 432 1594
rect 376 1470 432 1542
rect 376 1418 378 1470
rect 430 1418 432 1470
rect 376 1346 432 1418
rect 376 1294 378 1346
rect 430 1294 432 1346
rect 376 1058 432 1294
rect 376 1006 378 1058
rect 430 1006 432 1058
rect 376 934 432 1006
rect 376 882 378 934
rect 430 882 432 934
rect 376 810 432 882
rect 376 758 378 810
rect 430 758 432 810
rect 376 522 432 758
rect 376 470 378 522
rect 430 470 432 522
rect 376 398 432 470
rect 376 346 378 398
rect 430 346 432 398
rect 376 274 432 346
rect 376 222 378 274
rect 430 222 432 274
rect 376 -14 432 222
rect 376 -66 378 -14
rect 430 -66 432 -14
rect 376 -138 432 -66
rect 376 -190 378 -138
rect 430 -190 432 -138
rect 376 -262 432 -190
rect 376 -314 378 -262
rect 430 -314 432 -262
rect 376 -550 432 -314
rect 376 -602 378 -550
rect 430 -602 432 -550
rect 376 -674 432 -602
rect 376 -726 378 -674
rect 430 -726 432 -674
rect 376 -798 432 -726
rect 376 -850 378 -798
rect 430 -850 432 -798
rect 376 -1086 432 -850
rect 376 -1138 378 -1086
rect 430 -1138 432 -1086
rect 376 -1210 432 -1138
rect 376 -1262 378 -1210
rect 430 -1262 432 -1210
rect 376 -1334 432 -1262
rect 376 -1386 378 -1334
rect 430 -1386 432 -1334
rect 376 -1622 432 -1386
rect 376 -1674 378 -1622
rect 430 -1674 432 -1622
rect 376 -1746 432 -1674
rect 376 -1798 378 -1746
rect 430 -1798 432 -1746
rect 376 -1870 432 -1798
rect 376 -1922 378 -1870
rect 430 -1922 432 -1870
rect 376 -2141 432 -1922
rect 460 1792 516 2168
rect 846 2220 902 2226
rect 846 2168 848 2220
rect 900 2168 902 2220
rect 460 1740 462 1792
rect 514 1740 516 1792
rect 460 1684 516 1740
rect 460 1632 462 1684
rect 514 1632 516 1684
rect 460 1256 516 1632
rect 460 1204 462 1256
rect 514 1204 516 1256
rect 460 1148 516 1204
rect 460 1096 462 1148
rect 514 1096 516 1148
rect 460 720 516 1096
rect 460 668 462 720
rect 514 668 516 720
rect 460 612 516 668
rect 460 560 462 612
rect 514 560 516 612
rect 460 184 516 560
rect 460 132 462 184
rect 514 132 516 184
rect 460 76 516 132
rect 460 24 462 76
rect 514 24 516 76
rect 460 -352 516 24
rect 460 -404 462 -352
rect 514 -404 516 -352
rect 460 -460 516 -404
rect 460 -512 462 -460
rect 514 -512 516 -460
rect 460 -888 516 -512
rect 460 -940 462 -888
rect 514 -940 516 -888
rect 460 -996 516 -940
rect 460 -1048 462 -996
rect 514 -1048 516 -996
rect 460 -1424 516 -1048
rect 460 -1476 462 -1424
rect 514 -1476 516 -1424
rect 460 -1532 516 -1476
rect 460 -1584 462 -1532
rect 514 -1584 516 -1532
rect 460 -1960 516 -1584
rect 544 2130 600 2136
rect 544 2078 546 2130
rect 598 2078 600 2130
rect 544 2006 600 2078
rect 544 1954 546 2006
rect 598 1954 600 2006
rect 544 1882 600 1954
rect 544 1830 546 1882
rect 598 1830 600 1882
rect 544 1594 600 1830
rect 544 1542 546 1594
rect 598 1542 600 1594
rect 544 1470 600 1542
rect 544 1418 546 1470
rect 598 1418 600 1470
rect 544 1346 600 1418
rect 544 1294 546 1346
rect 598 1294 600 1346
rect 544 1058 600 1294
rect 544 1006 546 1058
rect 598 1006 600 1058
rect 544 934 600 1006
rect 544 882 546 934
rect 598 882 600 934
rect 544 810 600 882
rect 544 758 546 810
rect 598 758 600 810
rect 544 522 600 758
rect 544 470 546 522
rect 598 470 600 522
rect 544 398 600 470
rect 544 346 546 398
rect 598 346 600 398
rect 544 274 600 346
rect 544 222 546 274
rect 598 222 600 274
rect 544 -14 600 222
rect 544 -66 546 -14
rect 598 -66 600 -14
rect 544 -138 600 -66
rect 544 -190 546 -138
rect 598 -190 600 -138
rect 544 -262 600 -190
rect 544 -314 546 -262
rect 598 -314 600 -262
rect 544 -550 600 -314
rect 544 -602 546 -550
rect 598 -602 600 -550
rect 544 -674 600 -602
rect 544 -726 546 -674
rect 598 -726 600 -674
rect 544 -798 600 -726
rect 544 -850 546 -798
rect 598 -850 600 -798
rect 544 -1086 600 -850
rect 544 -1138 546 -1086
rect 598 -1138 600 -1086
rect 544 -1210 600 -1138
rect 544 -1262 546 -1210
rect 598 -1262 600 -1210
rect 544 -1334 600 -1262
rect 544 -1386 546 -1334
rect 598 -1386 600 -1334
rect 544 -1622 600 -1386
rect 544 -1674 546 -1622
rect 598 -1674 600 -1622
rect 544 -1746 600 -1674
rect 544 -1798 546 -1746
rect 598 -1798 600 -1746
rect 544 -1870 600 -1798
rect 544 -1922 546 -1870
rect 598 -1922 600 -1870
rect 544 -1928 600 -1922
rect 762 2130 818 2136
rect 762 2078 764 2130
rect 816 2078 818 2130
rect 762 2006 818 2078
rect 762 1954 764 2006
rect 816 1954 818 2006
rect 762 1882 818 1954
rect 762 1830 764 1882
rect 816 1830 818 1882
rect 762 1594 818 1830
rect 762 1542 764 1594
rect 816 1542 818 1594
rect 762 1470 818 1542
rect 762 1418 764 1470
rect 816 1418 818 1470
rect 762 1346 818 1418
rect 762 1294 764 1346
rect 816 1294 818 1346
rect 762 1058 818 1294
rect 762 1006 764 1058
rect 816 1006 818 1058
rect 762 934 818 1006
rect 762 882 764 934
rect 816 882 818 934
rect 762 810 818 882
rect 762 758 764 810
rect 816 758 818 810
rect 762 522 818 758
rect 762 470 764 522
rect 816 470 818 522
rect 762 398 818 470
rect 762 346 764 398
rect 816 346 818 398
rect 762 274 818 346
rect 762 222 764 274
rect 816 222 818 274
rect 762 -14 818 222
rect 762 -66 764 -14
rect 816 -66 818 -14
rect 762 -138 818 -66
rect 762 -190 764 -138
rect 816 -190 818 -138
rect 762 -262 818 -190
rect 762 -314 764 -262
rect 816 -314 818 -262
rect 762 -550 818 -314
rect 762 -602 764 -550
rect 816 -602 818 -550
rect 762 -674 818 -602
rect 762 -726 764 -674
rect 816 -726 818 -674
rect 762 -798 818 -726
rect 762 -850 764 -798
rect 816 -850 818 -798
rect 762 -1086 818 -850
rect 762 -1138 764 -1086
rect 816 -1138 818 -1086
rect 762 -1210 818 -1138
rect 762 -1262 764 -1210
rect 816 -1262 818 -1210
rect 762 -1334 818 -1262
rect 762 -1386 764 -1334
rect 816 -1386 818 -1334
rect 762 -1622 818 -1386
rect 762 -1674 764 -1622
rect 816 -1674 818 -1622
rect 762 -1746 818 -1674
rect 762 -1798 764 -1746
rect 816 -1798 818 -1746
rect 762 -1870 818 -1798
rect 762 -1922 764 -1870
rect 816 -1922 818 -1870
rect 762 -1928 818 -1922
rect 846 1792 902 2168
rect 846 1740 848 1792
rect 900 1740 902 1792
rect 846 1684 902 1740
rect 846 1632 848 1684
rect 900 1632 902 1684
rect 846 1256 902 1632
rect 846 1204 848 1256
rect 900 1204 902 1256
rect 846 1148 902 1204
rect 846 1096 848 1148
rect 900 1096 902 1148
rect 846 720 902 1096
rect 846 668 848 720
rect 900 668 902 720
rect 846 612 902 668
rect 846 560 848 612
rect 900 560 902 612
rect 846 184 902 560
rect 846 132 848 184
rect 900 132 902 184
rect 846 76 902 132
rect 846 24 848 76
rect 900 24 902 76
rect 846 -352 902 24
rect 846 -404 848 -352
rect 900 -404 902 -352
rect 846 -460 902 -404
rect 846 -512 848 -460
rect 900 -512 902 -460
rect 846 -888 902 -512
rect 846 -940 848 -888
rect 900 -940 902 -888
rect 846 -996 902 -940
rect 846 -1048 848 -996
rect 900 -1048 902 -996
rect 846 -1424 902 -1048
rect 846 -1476 848 -1424
rect 900 -1476 902 -1424
rect 846 -1532 902 -1476
rect 846 -1584 848 -1532
rect 900 -1584 902 -1532
rect 460 -2012 462 -1960
rect 514 -2012 516 -1960
rect 460 -2040 516 -2012
rect 846 -1960 902 -1584
rect 930 2130 986 2136
rect 930 2078 932 2130
rect 984 2078 986 2130
rect 930 2006 986 2078
rect 930 1954 932 2006
rect 984 1954 986 2006
rect 930 1882 986 1954
rect 930 1830 932 1882
rect 984 1830 986 1882
rect 930 1594 986 1830
rect 930 1542 932 1594
rect 984 1542 986 1594
rect 930 1470 986 1542
rect 930 1418 932 1470
rect 984 1418 986 1470
rect 930 1346 986 1418
rect 930 1294 932 1346
rect 984 1294 986 1346
rect 930 1058 986 1294
rect 930 1006 932 1058
rect 984 1006 986 1058
rect 930 934 986 1006
rect 930 882 932 934
rect 984 882 986 934
rect 930 810 986 882
rect 930 758 932 810
rect 984 758 986 810
rect 930 522 986 758
rect 930 470 932 522
rect 984 470 986 522
rect 930 398 986 470
rect 1338 476 1394 482
rect 1338 424 1340 476
rect 1392 424 1394 476
rect 930 346 932 398
rect 984 346 986 398
rect 930 274 986 346
rect 930 222 932 274
rect 984 222 986 274
rect 930 -14 986 222
rect 930 -66 932 -14
rect 984 -66 986 -14
rect 930 -138 986 -66
rect 930 -190 932 -138
rect 984 -190 986 -138
rect 930 -262 986 -190
rect 930 -314 932 -262
rect 984 -314 986 -262
rect 930 -550 986 -314
rect 930 -602 932 -550
rect 984 -602 986 -550
rect 930 -674 986 -602
rect 930 -726 932 -674
rect 984 -726 986 -674
rect 930 -798 986 -726
rect 930 -850 932 -798
rect 984 -850 986 -798
rect 930 -1086 986 -850
rect 930 -1138 932 -1086
rect 984 -1138 986 -1086
rect 930 -1210 986 -1138
rect 930 -1262 932 -1210
rect 984 -1262 986 -1210
rect 930 -1334 986 -1262
rect 930 -1386 932 -1334
rect 984 -1386 986 -1334
rect 930 -1622 986 -1386
rect 930 -1674 932 -1622
rect 984 -1674 986 -1622
rect 930 -1746 986 -1674
rect 930 -1798 932 -1746
rect 984 -1798 986 -1746
rect 930 -1870 986 -1798
rect 930 -1922 932 -1870
rect 984 -1922 986 -1870
rect 930 -1928 986 -1922
rect 1254 347 1310 401
rect 1254 295 1256 347
rect 1308 295 1310 347
rect 1254 29 1310 295
rect 1254 -23 1256 29
rect 1308 -23 1310 29
rect 1254 -289 1310 -23
rect 1254 -341 1256 -289
rect 1308 -341 1310 -289
rect 1254 -607 1310 -341
rect 1254 -659 1256 -607
rect 1308 -659 1310 -607
rect 1254 -925 1310 -659
rect 1254 -977 1256 -925
rect 1308 -977 1310 -925
rect 1254 -1243 1310 -977
rect 1254 -1295 1256 -1243
rect 1308 -1295 1310 -1243
rect 1254 -1561 1310 -1295
rect 1254 -1613 1256 -1561
rect 1308 -1613 1310 -1561
rect 1254 -1879 1310 -1613
rect 1254 -1931 1256 -1879
rect 1308 -1931 1310 -1879
rect 1254 -1937 1310 -1931
rect 1338 266 1394 424
rect 1724 476 1780 482
rect 1724 424 1726 476
rect 1778 424 1780 476
rect 1338 214 1340 266
rect 1392 214 1394 266
rect 1338 158 1394 214
rect 1338 106 1340 158
rect 1392 106 1394 158
rect 1338 -52 1394 106
rect 1338 -104 1340 -52
rect 1392 -104 1394 -52
rect 1338 -160 1394 -104
rect 1338 -212 1340 -160
rect 1392 -212 1394 -160
rect 1338 -370 1394 -212
rect 1338 -422 1340 -370
rect 1392 -422 1394 -370
rect 1338 -478 1394 -422
rect 1338 -530 1340 -478
rect 1392 -530 1394 -478
rect 1338 -688 1394 -530
rect 1338 -740 1340 -688
rect 1392 -740 1394 -688
rect 1338 -796 1394 -740
rect 1338 -848 1340 -796
rect 1392 -848 1394 -796
rect 1338 -1006 1394 -848
rect 1338 -1058 1340 -1006
rect 1392 -1058 1394 -1006
rect 1338 -1114 1394 -1058
rect 1338 -1166 1340 -1114
rect 1392 -1166 1394 -1114
rect 1338 -1324 1394 -1166
rect 1338 -1376 1340 -1324
rect 1392 -1376 1394 -1324
rect 1338 -1432 1394 -1376
rect 1338 -1484 1340 -1432
rect 1392 -1484 1394 -1432
rect 1338 -1642 1394 -1484
rect 1338 -1694 1340 -1642
rect 1392 -1694 1394 -1642
rect 1338 -1750 1394 -1694
rect 1338 -1802 1340 -1750
rect 1392 -1802 1394 -1750
rect 846 -2012 848 -1960
rect 900 -2012 902 -1960
rect 846 -2018 902 -2012
rect 1338 -1960 1394 -1802
rect 1422 347 1478 401
rect 1422 295 1424 347
rect 1476 295 1478 347
rect 1422 29 1478 295
rect 1422 -23 1424 29
rect 1476 -23 1478 29
rect 1422 -289 1478 -23
rect 1422 -341 1424 -289
rect 1476 -341 1478 -289
rect 1422 -607 1478 -341
rect 1422 -659 1424 -607
rect 1476 -659 1478 -607
rect 1422 -925 1478 -659
rect 1422 -977 1424 -925
rect 1476 -977 1478 -925
rect 1422 -1243 1478 -977
rect 1422 -1295 1424 -1243
rect 1476 -1295 1478 -1243
rect 1422 -1561 1478 -1295
rect 1422 -1613 1424 -1561
rect 1476 -1613 1478 -1561
rect 1422 -1879 1478 -1613
rect 1422 -1931 1424 -1879
rect 1476 -1931 1478 -1879
rect 1422 -1937 1478 -1931
rect 1640 347 1696 401
rect 1640 295 1642 347
rect 1694 295 1696 347
rect 1640 29 1696 295
rect 1640 -23 1642 29
rect 1694 -23 1696 29
rect 1640 -289 1696 -23
rect 1640 -341 1642 -289
rect 1694 -341 1696 -289
rect 1640 -607 1696 -341
rect 1640 -659 1642 -607
rect 1694 -659 1696 -607
rect 1640 -925 1696 -659
rect 1640 -977 1642 -925
rect 1694 -977 1696 -925
rect 1640 -1243 1696 -977
rect 1640 -1295 1642 -1243
rect 1694 -1295 1696 -1243
rect 1640 -1561 1696 -1295
rect 1640 -1613 1642 -1561
rect 1694 -1613 1696 -1561
rect 1640 -1879 1696 -1613
rect 1640 -1931 1642 -1879
rect 1694 -1931 1696 -1879
rect 1640 -1937 1696 -1931
rect 1724 266 1780 424
rect 1724 214 1726 266
rect 1778 214 1780 266
rect 1724 158 1780 214
rect 1724 106 1726 158
rect 1778 106 1780 158
rect 1724 -52 1780 106
rect 1724 -104 1726 -52
rect 1778 -104 1780 -52
rect 1724 -160 1780 -104
rect 1724 -212 1726 -160
rect 1778 -212 1780 -160
rect 1724 -370 1780 -212
rect 1724 -422 1726 -370
rect 1778 -422 1780 -370
rect 1724 -478 1780 -422
rect 1724 -530 1726 -478
rect 1778 -530 1780 -478
rect 1724 -688 1780 -530
rect 1724 -740 1726 -688
rect 1778 -740 1780 -688
rect 1724 -796 1780 -740
rect 1724 -848 1726 -796
rect 1778 -848 1780 -796
rect 1724 -1006 1780 -848
rect 1724 -1058 1726 -1006
rect 1778 -1058 1780 -1006
rect 1724 -1114 1780 -1058
rect 1724 -1166 1726 -1114
rect 1778 -1166 1780 -1114
rect 1724 -1324 1780 -1166
rect 1724 -1376 1726 -1324
rect 1778 -1376 1780 -1324
rect 1724 -1432 1780 -1376
rect 1724 -1484 1726 -1432
rect 1778 -1484 1780 -1432
rect 1724 -1642 1780 -1484
rect 1724 -1694 1726 -1642
rect 1778 -1694 1780 -1642
rect 1724 -1750 1780 -1694
rect 1724 -1802 1726 -1750
rect 1778 -1802 1780 -1750
rect 1338 -2012 1340 -1960
rect 1392 -2012 1394 -1960
rect 1338 -2018 1394 -2012
rect 1724 -1960 1780 -1802
rect 1724 -2012 1726 -1960
rect 1778 -2012 1780 -1960
rect 460 -2092 462 -2040
rect 514 -2092 516 -2040
rect 460 -2098 516 -2092
rect 1724 -2040 1780 -2012
rect 1724 -2092 1726 -2040
rect 1778 -2092 1780 -2040
rect 1724 -2098 1780 -2092
rect 1808 347 1864 401
rect 1808 295 1810 347
rect 1862 295 1864 347
rect 1808 29 1864 295
rect 1808 -23 1810 29
rect 1862 -23 1864 29
rect 1808 -289 1864 -23
rect 1808 -341 1810 -289
rect 1862 -341 1864 -289
rect 1808 -607 1864 -341
rect 1808 -659 1810 -607
rect 1862 -659 1864 -607
rect 1808 -925 1864 -659
rect 1808 -977 1810 -925
rect 1862 -977 1864 -925
rect 1808 -1243 1864 -977
rect 1808 -1295 1810 -1243
rect 1862 -1295 1864 -1243
rect 1808 -1561 1864 -1295
rect 1808 -1613 1810 -1561
rect 1862 -1613 1864 -1561
rect 1808 -1879 1864 -1613
rect 1808 -1931 1810 -1879
rect 1862 -1931 1864 -1879
rect 376 -2231 378 -2141
rect 430 -2231 432 -2141
rect 376 -2237 432 -2231
rect 1808 -2265 1864 -1931
rect 1808 -2355 1810 -2265
rect 1862 -2355 1864 -2265
rect 1808 -2361 1864 -2355
use sky130_fd_pr__pfet_01v8_TMYUV5  XM1
timestamp 1730624594
transform 1 0 488 0 1 104
box -246 -2245 246 2245
use sky130_fd_pr__pfet_01v8_TMYUV5  XM2
timestamp 1730624594
transform 1 0 874 0 1 104
box -246 -2245 246 2245
use sky130_fd_pr__nfet_01v8_KDBLWN  XM3
timestamp 1730624594
transform 1 0 1366 0 1 -768
box -246 -1373 246 1373
use sky130_fd_pr__nfet_01v8_KDBLWN  XM4
timestamp 1730624594
transform 1 0 1752 0 1 -768
box -246 -1373 246 1373
<< labels >>
flabel metal1 242 -2237 338 -2141 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel metal1 242 -2361 338 -2265 0 FreeSans 320 0 0 0 vssa
port 5 nsew
flabel via1 848 -2012 900 -1960 0 FreeSans 320 0 0 0 ckb
port 4 nsew
flabel via1 1340 -2012 1392 -1960 0 FreeSans 320 0 0 0 ck
port 3 nsew
flabel via1 932 2078 984 2130 0 FreeSans 320 0 0 0 out
port 6 nsew
flabel via1 1726 424 1778 476 0 FreeSans 320 0 0 0 in
port 2 nsew
<< end >>
