magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect 105 -1958 139 -1882
rect 105 -2048 139 -2042
rect 491 -1958 525 -1882
rect 491 -2048 525 -2042
rect 597 -2082 631 -1882
rect 597 -2172 631 -2166
rect 983 -2082 1017 -1882
rect 983 -2172 1017 -2166
<< viali >>
rect 105 -2042 139 -1958
rect 491 -2042 525 -1958
rect 597 -2166 631 -2082
rect 983 -2166 1017 -2082
<< metal1 >>
rect 269 2357 289 2409
rect 341 2357 361 2409
rect 199 2267 205 2319
rect 257 2267 263 2319
rect 199 2195 263 2267
rect 199 2143 205 2195
rect 257 2143 263 2195
rect 199 2071 263 2143
rect 199 2019 205 2071
rect 257 2019 263 2071
rect 367 2267 373 2319
rect 425 2267 431 2319
rect 367 2195 431 2267
rect 367 2143 373 2195
rect 425 2143 431 2195
rect 367 2071 431 2143
rect 367 2019 373 2071
rect 425 2019 431 2071
rect 269 1929 289 1981
rect 341 1929 361 1981
rect 269 1821 289 1873
rect 341 1821 361 1873
rect 199 1731 205 1783
rect 257 1731 263 1783
rect 199 1659 263 1731
rect 199 1607 205 1659
rect 257 1607 263 1659
rect 199 1535 263 1607
rect 199 1483 205 1535
rect 257 1483 263 1535
rect 367 1731 373 1783
rect 425 1731 431 1783
rect 367 1659 431 1731
rect 367 1607 373 1659
rect 425 1607 431 1659
rect 367 1535 431 1607
rect 367 1483 373 1535
rect 425 1483 431 1535
rect 269 1393 289 1445
rect 341 1393 361 1445
rect 269 1285 289 1337
rect 341 1285 361 1337
rect 199 1195 205 1247
rect 257 1195 263 1247
rect 199 1123 263 1195
rect 199 1071 205 1123
rect 257 1071 263 1123
rect 199 999 263 1071
rect 199 947 205 999
rect 257 947 263 999
rect 367 1195 373 1247
rect 425 1195 431 1247
rect 367 1123 431 1195
rect 367 1071 373 1123
rect 425 1071 431 1123
rect 367 999 431 1071
rect 367 947 373 999
rect 425 947 431 999
rect 269 857 289 909
rect 341 857 361 909
rect 269 749 289 801
rect 341 749 361 801
rect 199 659 205 711
rect 257 659 263 711
rect 199 587 263 659
rect 199 535 205 587
rect 257 535 263 587
rect 199 463 263 535
rect 199 411 205 463
rect 257 411 263 463
rect 367 659 373 711
rect 425 659 431 711
rect 367 587 431 659
rect 761 613 781 665
rect 833 613 853 665
rect 367 535 373 587
rect 425 535 431 587
rect 367 463 431 535
rect 691 536 755 584
rect 691 484 697 536
rect 749 484 755 536
rect 859 536 923 584
rect 859 484 865 536
rect 917 484 923 536
rect 367 411 373 463
rect 425 411 431 463
rect 367 402 431 411
rect 761 403 781 455
rect 833 403 853 455
rect 269 321 289 373
rect 341 321 361 373
rect 761 295 781 347
rect 833 295 853 347
rect 269 213 289 265
rect 341 213 361 265
rect 691 218 755 266
rect 199 123 205 175
rect 257 123 263 175
rect 199 51 263 123
rect 199 -1 205 51
rect 257 -1 263 51
rect 199 -73 263 -1
rect 199 -125 205 -73
rect 257 -125 263 -73
rect 367 123 373 175
rect 425 123 431 175
rect 691 166 697 218
rect 749 166 755 218
rect 859 218 923 266
rect 859 166 865 218
rect 917 166 923 218
rect 367 51 431 123
rect 761 85 781 137
rect 833 85 853 137
rect 367 -1 373 51
rect 425 -1 431 51
rect 367 -73 431 -1
rect 761 -23 781 29
rect 833 -23 853 29
rect 367 -125 373 -73
rect 425 -125 431 -73
rect 691 -100 755 -52
rect 691 -152 697 -100
rect 749 -152 755 -100
rect 859 -100 923 -52
rect 859 -152 865 -100
rect 917 -152 923 -100
rect 269 -215 289 -163
rect 341 -215 361 -163
rect 761 -233 781 -181
rect 833 -233 853 -181
rect 269 -323 289 -271
rect 341 -323 361 -271
rect 761 -341 781 -289
rect 833 -341 853 -289
rect 199 -413 205 -361
rect 257 -413 263 -361
rect 199 -485 263 -413
rect 199 -537 205 -485
rect 257 -537 263 -485
rect 199 -609 263 -537
rect 199 -661 205 -609
rect 257 -661 263 -609
rect 367 -413 373 -361
rect 425 -413 431 -361
rect 367 -485 431 -413
rect 691 -418 755 -370
rect 691 -470 697 -418
rect 749 -470 755 -418
rect 859 -418 923 -370
rect 859 -470 865 -418
rect 917 -470 923 -418
rect 367 -537 373 -485
rect 425 -537 431 -485
rect 367 -609 431 -537
rect 761 -551 781 -499
rect 833 -551 853 -499
rect 367 -661 373 -609
rect 425 -661 431 -609
rect 761 -659 781 -607
rect 833 -659 853 -607
rect 269 -751 289 -699
rect 341 -751 361 -699
rect 691 -736 755 -688
rect 691 -788 697 -736
rect 749 -788 755 -736
rect 859 -736 923 -688
rect 859 -788 865 -736
rect 917 -788 923 -736
rect 269 -859 289 -807
rect 341 -859 361 -807
rect 761 -869 781 -817
rect 833 -869 853 -817
rect 199 -949 205 -897
rect 257 -949 263 -897
rect 199 -1021 263 -949
rect 199 -1073 205 -1021
rect 257 -1073 263 -1021
rect 199 -1145 263 -1073
rect 199 -1197 205 -1145
rect 257 -1197 263 -1145
rect 367 -949 373 -897
rect 425 -949 431 -897
rect 367 -1006 431 -949
rect 761 -977 781 -925
rect 833 -977 853 -925
rect 367 -1021 755 -1006
rect 367 -1073 373 -1021
rect 425 -1054 755 -1021
rect 425 -1073 697 -1054
rect 367 -1106 697 -1073
rect 749 -1106 755 -1054
rect 859 -1054 923 -1006
rect 859 -1106 865 -1054
rect 917 -1106 923 -1054
rect 367 -1145 431 -1106
rect 367 -1197 373 -1145
rect 425 -1197 431 -1145
rect 761 -1187 781 -1135
rect 833 -1187 853 -1135
rect 269 -1287 289 -1235
rect 341 -1287 361 -1235
rect 761 -1295 781 -1243
rect 833 -1295 853 -1243
rect 269 -1395 289 -1343
rect 341 -1395 361 -1343
rect 691 -1372 755 -1324
rect 691 -1424 697 -1372
rect 749 -1424 755 -1372
rect 859 -1372 923 -1324
rect 859 -1424 865 -1372
rect 917 -1424 923 -1372
rect 199 -1485 205 -1433
rect 257 -1485 263 -1433
rect 199 -1557 263 -1485
rect 199 -1609 205 -1557
rect 257 -1609 263 -1557
rect 199 -1681 263 -1609
rect 199 -1733 205 -1681
rect 257 -1733 263 -1681
rect 367 -1485 373 -1433
rect 425 -1485 431 -1433
rect 367 -1557 431 -1485
rect 761 -1505 781 -1453
rect 833 -1505 853 -1453
rect 367 -1609 373 -1557
rect 425 -1609 431 -1557
rect 367 -1642 431 -1609
rect 761 -1613 781 -1561
rect 833 -1613 853 -1561
rect 367 -1681 755 -1642
rect 367 -1733 373 -1681
rect 425 -1690 755 -1681
rect 425 -1733 697 -1690
rect 367 -1742 697 -1733
rect 749 -1742 755 -1690
rect 859 -1690 923 -1642
rect 859 -1742 865 -1690
rect 917 -1742 923 -1690
rect 269 -1823 289 -1771
rect 341 -1823 361 -1771
rect 761 -1823 781 -1771
rect 833 -1823 853 -1771
rect 199 -1909 205 -1857
rect 257 -1909 865 -1857
rect 917 -1909 923 -1857
rect 69 -1958 1053 -1952
rect 69 -2042 105 -1958
rect 139 -2042 491 -1958
rect 525 -2042 1053 -1958
rect 69 -2048 1053 -2042
rect 69 -2082 1053 -2076
rect 69 -2166 597 -2082
rect 631 -2166 983 -2082
rect 1017 -2166 1053 -2082
rect 69 -2172 1053 -2166
rect 69 -2252 205 -2200
rect 257 -2252 1053 -2200
rect 69 -2258 1053 -2252
<< via1 >>
rect 289 2357 341 2409
rect 205 2267 257 2319
rect 205 2143 257 2195
rect 205 2019 257 2071
rect 373 2267 425 2319
rect 373 2143 425 2195
rect 373 2019 425 2071
rect 289 1929 341 1981
rect 289 1821 341 1873
rect 205 1731 257 1783
rect 205 1607 257 1659
rect 205 1483 257 1535
rect 373 1731 425 1783
rect 373 1607 425 1659
rect 373 1483 425 1535
rect 289 1393 341 1445
rect 289 1285 341 1337
rect 205 1195 257 1247
rect 205 1071 257 1123
rect 205 947 257 999
rect 373 1195 425 1247
rect 373 1071 425 1123
rect 373 947 425 999
rect 289 857 341 909
rect 289 749 341 801
rect 205 659 257 711
rect 205 535 257 587
rect 205 411 257 463
rect 373 659 425 711
rect 781 613 833 665
rect 373 535 425 587
rect 697 484 749 536
rect 865 484 917 536
rect 373 411 425 463
rect 781 403 833 455
rect 289 321 341 373
rect 781 295 833 347
rect 289 213 341 265
rect 205 123 257 175
rect 205 -1 257 51
rect 205 -125 257 -73
rect 373 123 425 175
rect 697 166 749 218
rect 865 166 917 218
rect 781 85 833 137
rect 373 -1 425 51
rect 781 -23 833 29
rect 373 -125 425 -73
rect 697 -152 749 -100
rect 865 -152 917 -100
rect 289 -215 341 -163
rect 781 -233 833 -181
rect 289 -323 341 -271
rect 781 -341 833 -289
rect 205 -413 257 -361
rect 205 -537 257 -485
rect 205 -661 257 -609
rect 373 -413 425 -361
rect 697 -470 749 -418
rect 865 -470 917 -418
rect 373 -537 425 -485
rect 781 -551 833 -499
rect 373 -661 425 -609
rect 781 -659 833 -607
rect 289 -751 341 -699
rect 697 -788 749 -736
rect 865 -788 917 -736
rect 289 -859 341 -807
rect 781 -869 833 -817
rect 205 -949 257 -897
rect 205 -1073 257 -1021
rect 205 -1197 257 -1145
rect 373 -949 425 -897
rect 781 -977 833 -925
rect 373 -1073 425 -1021
rect 697 -1106 749 -1054
rect 865 -1106 917 -1054
rect 373 -1197 425 -1145
rect 781 -1187 833 -1135
rect 289 -1287 341 -1235
rect 781 -1295 833 -1243
rect 289 -1395 341 -1343
rect 697 -1424 749 -1372
rect 865 -1424 917 -1372
rect 205 -1485 257 -1433
rect 205 -1609 257 -1557
rect 205 -1733 257 -1681
rect 373 -1485 425 -1433
rect 781 -1505 833 -1453
rect 373 -1609 425 -1557
rect 781 -1613 833 -1561
rect 373 -1733 425 -1681
rect 697 -1742 749 -1690
rect 865 -1742 917 -1690
rect 289 -1823 341 -1771
rect 781 -1823 833 -1771
rect 205 -1909 257 -1857
rect 865 -1909 917 -1857
rect 205 -2252 257 -2200
<< metal2 >>
rect 287 2409 343 2415
rect 287 2357 289 2409
rect 341 2357 343 2409
rect 203 2319 259 2325
rect 203 2267 205 2319
rect 257 2267 259 2319
rect 203 2195 259 2267
rect 203 2143 205 2195
rect 257 2143 259 2195
rect 203 2071 259 2143
rect 203 2019 205 2071
rect 257 2019 259 2071
rect 203 1783 259 2019
rect 203 1731 205 1783
rect 257 1731 259 1783
rect 203 1659 259 1731
rect 203 1607 205 1659
rect 257 1607 259 1659
rect 203 1535 259 1607
rect 203 1483 205 1535
rect 257 1483 259 1535
rect 203 1247 259 1483
rect 203 1195 205 1247
rect 257 1195 259 1247
rect 203 1123 259 1195
rect 203 1071 205 1123
rect 257 1071 259 1123
rect 203 999 259 1071
rect 203 947 205 999
rect 257 947 259 999
rect 203 711 259 947
rect 203 659 205 711
rect 257 659 259 711
rect 203 587 259 659
rect 203 535 205 587
rect 257 535 259 587
rect 203 463 259 535
rect 203 411 205 463
rect 257 411 259 463
rect 203 175 259 411
rect 203 123 205 175
rect 257 123 259 175
rect 203 51 259 123
rect 203 -1 205 51
rect 257 -1 259 51
rect 203 -73 259 -1
rect 203 -125 205 -73
rect 257 -125 259 -73
rect 203 -361 259 -125
rect 203 -413 205 -361
rect 257 -413 259 -361
rect 203 -485 259 -413
rect 203 -537 205 -485
rect 257 -537 259 -485
rect 203 -609 259 -537
rect 203 -661 205 -609
rect 257 -661 259 -609
rect 203 -897 259 -661
rect 203 -949 205 -897
rect 257 -949 259 -897
rect 203 -1021 259 -949
rect 203 -1073 205 -1021
rect 257 -1073 259 -1021
rect 203 -1145 259 -1073
rect 203 -1197 205 -1145
rect 257 -1197 259 -1145
rect 203 -1433 259 -1197
rect 203 -1485 205 -1433
rect 257 -1485 259 -1433
rect 203 -1557 259 -1485
rect 203 -1609 205 -1557
rect 257 -1609 259 -1557
rect 203 -1681 259 -1609
rect 203 -1733 205 -1681
rect 257 -1733 259 -1681
rect 203 -1857 259 -1733
rect 287 1981 343 2357
rect 287 1929 289 1981
rect 341 1929 343 1981
rect 287 1873 343 1929
rect 287 1821 289 1873
rect 341 1821 343 1873
rect 287 1445 343 1821
rect 287 1393 289 1445
rect 341 1393 343 1445
rect 287 1337 343 1393
rect 287 1285 289 1337
rect 341 1285 343 1337
rect 287 909 343 1285
rect 287 857 289 909
rect 341 857 343 909
rect 287 801 343 857
rect 287 749 289 801
rect 341 749 343 801
rect 287 373 343 749
rect 287 321 289 373
rect 341 321 343 373
rect 287 265 343 321
rect 287 213 289 265
rect 341 213 343 265
rect 287 -163 343 213
rect 287 -215 289 -163
rect 341 -215 343 -163
rect 287 -271 343 -215
rect 287 -323 289 -271
rect 341 -323 343 -271
rect 287 -699 343 -323
rect 287 -751 289 -699
rect 341 -751 343 -699
rect 287 -807 343 -751
rect 287 -859 289 -807
rect 341 -859 343 -807
rect 287 -1235 343 -859
rect 287 -1287 289 -1235
rect 341 -1287 343 -1235
rect 287 -1343 343 -1287
rect 287 -1395 289 -1343
rect 341 -1395 343 -1343
rect 287 -1771 343 -1395
rect 371 2319 427 2325
rect 371 2267 373 2319
rect 425 2267 427 2319
rect 371 2195 427 2267
rect 371 2143 373 2195
rect 425 2143 427 2195
rect 371 2071 427 2143
rect 371 2019 373 2071
rect 425 2019 427 2071
rect 371 1783 427 2019
rect 371 1731 373 1783
rect 425 1731 427 1783
rect 371 1659 427 1731
rect 371 1607 373 1659
rect 425 1607 427 1659
rect 371 1535 427 1607
rect 371 1483 373 1535
rect 425 1483 427 1535
rect 371 1247 427 1483
rect 371 1195 373 1247
rect 425 1195 427 1247
rect 371 1123 427 1195
rect 371 1071 373 1123
rect 425 1071 427 1123
rect 371 999 427 1071
rect 371 947 373 999
rect 425 947 427 999
rect 371 711 427 947
rect 371 659 373 711
rect 425 659 427 711
rect 371 587 427 659
rect 779 665 835 671
rect 779 613 781 665
rect 833 613 835 665
rect 371 535 373 587
rect 425 535 427 587
rect 371 463 427 535
rect 371 411 373 463
rect 425 411 427 463
rect 371 175 427 411
rect 371 123 373 175
rect 425 123 427 175
rect 371 51 427 123
rect 371 -1 373 51
rect 425 -1 427 51
rect 371 -73 427 -1
rect 371 -125 373 -73
rect 425 -125 427 -73
rect 371 -361 427 -125
rect 371 -413 373 -361
rect 425 -413 427 -361
rect 371 -485 427 -413
rect 371 -537 373 -485
rect 425 -537 427 -485
rect 371 -609 427 -537
rect 371 -661 373 -609
rect 425 -661 427 -609
rect 371 -897 427 -661
rect 371 -949 373 -897
rect 425 -949 427 -897
rect 371 -1021 427 -949
rect 371 -1073 373 -1021
rect 425 -1073 427 -1021
rect 371 -1145 427 -1073
rect 371 -1197 373 -1145
rect 425 -1197 427 -1145
rect 371 -1433 427 -1197
rect 371 -1485 373 -1433
rect 425 -1485 427 -1433
rect 371 -1557 427 -1485
rect 371 -1609 373 -1557
rect 425 -1609 427 -1557
rect 371 -1681 427 -1609
rect 371 -1733 373 -1681
rect 425 -1733 427 -1681
rect 371 -1739 427 -1733
rect 695 536 751 590
rect 695 484 697 536
rect 749 484 751 536
rect 695 218 751 484
rect 695 166 697 218
rect 749 166 751 218
rect 695 -100 751 166
rect 695 -152 697 -100
rect 749 -152 751 -100
rect 695 -418 751 -152
rect 695 -470 697 -418
rect 749 -470 751 -418
rect 695 -736 751 -470
rect 695 -788 697 -736
rect 749 -788 751 -736
rect 695 -1054 751 -788
rect 695 -1106 697 -1054
rect 749 -1106 751 -1054
rect 695 -1372 751 -1106
rect 695 -1424 697 -1372
rect 749 -1424 751 -1372
rect 695 -1690 751 -1424
rect 695 -1742 697 -1690
rect 749 -1742 751 -1690
rect 695 -1748 751 -1742
rect 779 455 835 613
rect 779 403 781 455
rect 833 403 835 455
rect 779 347 835 403
rect 779 295 781 347
rect 833 295 835 347
rect 779 137 835 295
rect 779 85 781 137
rect 833 85 835 137
rect 779 29 835 85
rect 779 -23 781 29
rect 833 -23 835 29
rect 779 -181 835 -23
rect 779 -233 781 -181
rect 833 -233 835 -181
rect 779 -289 835 -233
rect 779 -341 781 -289
rect 833 -341 835 -289
rect 779 -499 835 -341
rect 779 -551 781 -499
rect 833 -551 835 -499
rect 779 -607 835 -551
rect 779 -659 781 -607
rect 833 -659 835 -607
rect 779 -817 835 -659
rect 779 -869 781 -817
rect 833 -869 835 -817
rect 779 -925 835 -869
rect 779 -977 781 -925
rect 833 -977 835 -925
rect 779 -1135 835 -977
rect 779 -1187 781 -1135
rect 833 -1187 835 -1135
rect 779 -1243 835 -1187
rect 779 -1295 781 -1243
rect 833 -1295 835 -1243
rect 779 -1453 835 -1295
rect 779 -1505 781 -1453
rect 833 -1505 835 -1453
rect 779 -1561 835 -1505
rect 779 -1613 781 -1561
rect 833 -1613 835 -1561
rect 287 -1823 289 -1771
rect 341 -1823 343 -1771
rect 287 -1829 343 -1823
rect 779 -1771 835 -1613
rect 779 -1823 781 -1771
rect 833 -1823 835 -1771
rect 779 -1829 835 -1823
rect 863 536 919 590
rect 863 484 865 536
rect 917 484 919 536
rect 863 218 919 484
rect 863 166 865 218
rect 917 166 919 218
rect 863 -100 919 166
rect 863 -152 865 -100
rect 917 -152 919 -100
rect 863 -418 919 -152
rect 863 -470 865 -418
rect 917 -470 919 -418
rect 863 -736 919 -470
rect 863 -788 865 -736
rect 917 -788 919 -736
rect 863 -1054 919 -788
rect 863 -1106 865 -1054
rect 917 -1106 919 -1054
rect 863 -1372 919 -1106
rect 863 -1424 865 -1372
rect 917 -1424 919 -1372
rect 863 -1690 919 -1424
rect 863 -1742 865 -1690
rect 917 -1742 919 -1690
rect 203 -1909 205 -1857
rect 257 -1909 259 -1857
rect 203 -2200 259 -1909
rect 863 -1857 919 -1742
rect 863 -1909 865 -1857
rect 917 -1909 919 -1857
rect 863 -1915 919 -1909
rect 203 -2252 205 -2200
rect 257 -2252 259 -2200
rect 203 -2258 259 -2252
use sky130_fd_pr__pfet_01v8_TMYUV5  XM1
timestamp 1730624594
transform 1 0 315 0 1 293
box -246 -2245 246 2245
use sky130_fd_pr__nfet_01v8_KDBLWN  XM2
timestamp 1730624594
transform 1 0 807 0 1 -579
box -246 -1373 246 1373
<< labels >>
flabel metal1 69 -2048 165 -1952 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel metal1 69 -2172 165 -2076 0 FreeSans 320 0 0 0 vssa
port 4 nsew
flabel metal1 69 -2258 127 -2200 0 FreeSans 320 0 0 0 in
port 5 nsew
flabel via1 781 -1823 833 -1771 0 FreeSans 320 0 0 0 swn
port 3 nsew
flabel via1 289 -1823 341 -1771 0 FreeSans 320 0 0 0 swp
port 2 nsew
flabel via1 373 2267 425 2319 0 FreeSans 320 0 0 0 out
port 6 nsew
<< end >>
