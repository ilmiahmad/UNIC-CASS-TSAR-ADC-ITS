magic
tech sky130A
magscale 1 2
timestamp 1730903028
<< viali >>
rect 3893 12189 3927 12223
rect 4169 12121 4203 12155
rect 5641 12053 5675 12087
rect 4169 11849 4203 11883
rect 5917 11781 5951 11815
rect 2421 11713 2455 11747
rect 2697 11645 2731 11679
rect 6193 11645 6227 11679
rect 6469 11645 6503 11679
rect 6745 11645 6779 11679
rect 4445 11509 4479 11543
rect 8217 11509 8251 11543
rect 3525 11305 3559 11339
rect 5254 11305 5288 11339
rect 6745 11305 6779 11339
rect 10701 11305 10735 11339
rect 1777 11169 1811 11203
rect 4997 11169 5031 11203
rect 6929 11169 6963 11203
rect 8953 11169 8987 11203
rect 9229 11169 9263 11203
rect 2053 11033 2087 11067
rect 7205 11033 7239 11067
rect 8677 10965 8711 10999
rect 6791 10761 6825 10795
rect 9781 10761 9815 10795
rect 2421 10693 2455 10727
rect 8309 10693 8343 10727
rect 5917 10625 5951 10659
rect 6883 10625 6917 10659
rect 8033 10625 8067 10659
rect 2145 10557 2179 10591
rect 3893 10557 3927 10591
rect 5641 10557 5675 10591
rect 4169 10421 4203 10455
rect 1869 10217 1903 10251
rect 6469 10217 6503 10251
rect 11161 10217 11195 10251
rect 3341 10081 3375 10115
rect 3617 10081 3651 10115
rect 4721 10013 4755 10047
rect 4997 10013 5031 10047
rect 5089 10013 5123 10047
rect 9413 10013 9447 10047
rect 7757 9945 7791 9979
rect 9689 9945 9723 9979
rect 4721 9877 4755 9911
rect 4721 9537 4755 9571
rect 8217 9537 8251 9571
rect 7849 9469 7883 9503
rect 9413 9469 9447 9503
rect 9689 9469 9723 9503
rect 11161 9469 11195 9503
rect 4813 9333 4847 9367
rect 1501 9129 1535 9163
rect 3893 9129 3927 9163
rect 6837 9129 6871 9163
rect 10701 9129 10735 9163
rect 8309 8993 8343 9027
rect 8953 8993 8987 9027
rect 3249 8925 3283 8959
rect 5641 8925 5675 8959
rect 8585 8925 8619 8959
rect 10920 8925 10954 8959
rect 2973 8857 3007 8891
rect 5365 8857 5399 8891
rect 9229 8857 9263 8891
rect 11023 8789 11057 8823
rect 3801 8585 3835 8619
rect 8125 8585 8159 8619
rect 5273 8517 5307 8551
rect 6653 8517 6687 8551
rect 9321 8449 9355 8483
rect 1501 8381 1535 8415
rect 2973 8381 3007 8415
rect 3249 8381 3283 8415
rect 5549 8381 5583 8415
rect 6377 8381 6411 8415
rect 8493 8381 8527 8415
rect 1869 8041 1903 8075
rect 4077 8041 4111 8075
rect 7665 8041 7699 8075
rect 10701 8041 10735 8075
rect 3617 7905 3651 7939
rect 6193 7905 6227 7939
rect 9229 7905 9263 7939
rect 5825 7837 5859 7871
rect 5917 7837 5951 7871
rect 8953 7837 8987 7871
rect 3341 7769 3375 7803
rect 5549 7769 5583 7803
rect 8769 7769 8803 7803
rect 7205 7497 7239 7531
rect 8493 7429 8527 7463
rect 6193 7361 6227 7395
rect 8769 7361 8803 7395
rect 5825 7293 5859 7327
rect 8585 7293 8619 7327
rect 9045 7293 9079 7327
rect 9321 7293 9355 7327
rect 10793 7293 10827 7327
rect 8953 7157 8987 7191
rect 7769 6953 7803 6987
rect 8677 6953 8711 6987
rect 9952 6953 9986 6987
rect 3893 6817 3927 6851
rect 6285 6817 6319 6851
rect 8309 6817 8343 6851
rect 5641 6749 5675 6783
rect 8033 6749 8067 6783
rect 8493 6749 8527 6783
rect 9689 6749 9723 6783
rect 5365 6681 5399 6715
rect 11437 6613 11471 6647
rect 2053 6409 2087 6443
rect 4445 6409 4479 6443
rect 3525 6341 3559 6375
rect 7297 6341 7331 6375
rect 7021 6273 7055 6307
rect 3801 6205 3835 6239
rect 5917 6205 5951 6239
rect 6193 6205 6227 6239
rect 9505 6205 9539 6239
rect 9781 6205 9815 6239
rect 8769 6069 8803 6103
rect 11253 6069 11287 6103
rect 1869 5865 1903 5899
rect 3341 5729 3375 5763
rect 6561 5729 6595 5763
rect 9873 5729 9907 5763
rect 3617 5661 3651 5695
rect 6929 5661 6963 5695
rect 9597 5661 9631 5695
rect 6285 5593 6319 5627
rect 7205 5593 7239 5627
rect 4813 5525 4847 5559
rect 8677 5525 8711 5559
rect 11345 5525 11379 5559
rect 3617 5321 3651 5355
rect 5089 5253 5123 5287
rect 7573 5253 7607 5287
rect 3433 5185 3467 5219
rect 5365 5185 5399 5219
rect 3157 5117 3191 5151
rect 9413 5117 9447 5151
rect 9689 5117 9723 5151
rect 1685 4981 1719 5015
rect 9045 4981 9079 5015
rect 11161 4981 11195 5015
rect 3893 4777 3927 4811
rect 5383 4777 5417 4811
rect 7008 4777 7042 4811
rect 3341 4641 3375 4675
rect 3617 4641 3651 4675
rect 5641 4641 5675 4675
rect 6745 4641 6779 4675
rect 1869 4437 1903 4471
rect 8493 4437 8527 4471
rect 4537 4165 4571 4199
rect 7481 4165 7515 4199
rect 4261 4029 4295 4063
rect 6009 4029 6043 4063
rect 7205 4029 7239 4063
rect 9505 4029 9539 4063
rect 9781 4029 9815 4063
rect 8953 3893 8987 3927
rect 11253 3893 11287 3927
rect 6561 3553 6595 3587
rect 6837 3553 6871 3587
rect 6929 3553 6963 3587
rect 9597 3553 9631 3587
rect 9873 3553 9907 3587
rect 7192 3417 7226 3451
rect 5089 3349 5123 3383
rect 8677 3349 8711 3383
rect 11345 3349 11379 3383
rect 4445 3145 4479 3179
rect 6837 3145 6871 3179
rect 11253 3145 11287 3179
rect 8309 3077 8343 3111
rect 6193 3009 6227 3043
rect 8585 3009 8619 3043
rect 9505 3009 9539 3043
rect 5917 2941 5951 2975
rect 9781 2941 9815 2975
<< metal1 >>
rect 1104 12538 11868 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 6214 12538
rect 6266 12486 6278 12538
rect 6330 12486 6342 12538
rect 6394 12486 6406 12538
rect 6458 12486 6470 12538
rect 6522 12486 8214 12538
rect 8266 12486 8278 12538
rect 8330 12486 8342 12538
rect 8394 12486 8406 12538
rect 8458 12486 8470 12538
rect 8522 12486 10214 12538
rect 10266 12486 10278 12538
rect 10330 12486 10342 12538
rect 10394 12486 10406 12538
rect 10458 12486 10470 12538
rect 10522 12486 11868 12538
rect 1104 12464 11868 12486
rect 3602 12180 3608 12232
rect 3660 12220 3666 12232
rect 3881 12223 3939 12229
rect 3881 12220 3893 12223
rect 3660 12192 3893 12220
rect 3660 12180 3666 12192
rect 3881 12189 3893 12192
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 4154 12112 4160 12164
rect 4212 12112 4218 12164
rect 4540 12124 4646 12152
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 4062 12084 4068 12096
rect 2832 12056 4068 12084
rect 2832 12044 2838 12056
rect 4062 12044 4068 12056
rect 4120 12084 4126 12096
rect 4540 12084 4568 12124
rect 4120 12056 4568 12084
rect 5629 12087 5687 12093
rect 4120 12044 4126 12056
rect 5629 12053 5641 12087
rect 5675 12084 5687 12087
rect 5902 12084 5908 12096
rect 5675 12056 5908 12084
rect 5675 12053 5687 12056
rect 5629 12047 5687 12053
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 1104 11994 11868 12016
rect 1104 11942 4894 11994
rect 4946 11942 4958 11994
rect 5010 11942 5022 11994
rect 5074 11942 5086 11994
rect 5138 11942 5150 11994
rect 5202 11942 6894 11994
rect 6946 11942 6958 11994
rect 7010 11942 7022 11994
rect 7074 11942 7086 11994
rect 7138 11942 7150 11994
rect 7202 11942 8894 11994
rect 8946 11942 8958 11994
rect 9010 11942 9022 11994
rect 9074 11942 9086 11994
rect 9138 11942 9150 11994
rect 9202 11942 10894 11994
rect 10946 11942 10958 11994
rect 11010 11942 11022 11994
rect 11074 11942 11086 11994
rect 11138 11942 11150 11994
rect 11202 11942 11868 11994
rect 1104 11920 11868 11942
rect 3602 11880 3608 11892
rect 2424 11852 3608 11880
rect 2424 11753 2452 11852
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4154 11840 4160 11892
rect 4212 11840 4218 11892
rect 7650 11880 7656 11892
rect 4632 11852 7656 11880
rect 2774 11772 2780 11824
rect 2832 11812 2838 11824
rect 2832 11784 3174 11812
rect 2832 11772 2838 11784
rect 4062 11772 4068 11824
rect 4120 11812 4126 11824
rect 4632 11812 4660 11852
rect 4120 11784 4738 11812
rect 4120 11772 4126 11784
rect 5902 11772 5908 11824
rect 5960 11772 5966 11824
rect 6932 11812 6960 11852
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 6932 11784 7222 11812
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11713 2467 11747
rect 2409 11707 2467 11713
rect 2682 11636 2688 11688
rect 2740 11636 2746 11688
rect 6181 11679 6239 11685
rect 6181 11645 6193 11679
rect 6227 11676 6239 11679
rect 6454 11676 6460 11688
rect 6227 11648 6460 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 6730 11636 6736 11688
rect 6788 11636 6794 11688
rect 4433 11543 4491 11549
rect 4433 11509 4445 11543
rect 4479 11540 4491 11543
rect 4890 11540 4896 11552
rect 4479 11512 4896 11540
rect 4479 11509 4491 11512
rect 4433 11503 4491 11509
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7248 11512 8217 11540
rect 7248 11500 7254 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 1104 11450 11868 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 6214 11450
rect 6266 11398 6278 11450
rect 6330 11398 6342 11450
rect 6394 11398 6406 11450
rect 6458 11398 6470 11450
rect 6522 11398 8214 11450
rect 8266 11398 8278 11450
rect 8330 11398 8342 11450
rect 8394 11398 8406 11450
rect 8458 11398 8470 11450
rect 8522 11398 10214 11450
rect 10266 11398 10278 11450
rect 10330 11398 10342 11450
rect 10394 11398 10406 11450
rect 10458 11398 10470 11450
rect 10522 11398 11868 11450
rect 1104 11376 11868 11398
rect 2682 11296 2688 11348
rect 2740 11336 2746 11348
rect 3513 11339 3571 11345
rect 3513 11336 3525 11339
rect 2740 11308 3525 11336
rect 2740 11296 2746 11308
rect 3513 11305 3525 11308
rect 3559 11305 3571 11339
rect 3513 11299 3571 11305
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 5242 11339 5300 11345
rect 5242 11336 5254 11339
rect 4948 11308 5254 11336
rect 4948 11296 4954 11308
rect 5242 11305 5254 11308
rect 5288 11305 5300 11339
rect 5242 11299 5300 11305
rect 6730 11296 6736 11348
rect 6788 11296 6794 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 10689 11339 10747 11345
rect 10689 11336 10701 11339
rect 7340 11308 10701 11336
rect 7340 11296 7346 11308
rect 10689 11305 10701 11308
rect 10735 11305 10747 11339
rect 10689 11299 10747 11305
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11200 1823 11203
rect 3602 11200 3608 11212
rect 1811 11172 3608 11200
rect 1811 11169 1823 11172
rect 1765 11163 1823 11169
rect 3602 11160 3608 11172
rect 3660 11200 3666 11212
rect 4985 11203 5043 11209
rect 4985 11200 4997 11203
rect 3660 11172 4997 11200
rect 3660 11160 3666 11172
rect 4985 11169 4997 11172
rect 5031 11200 5043 11203
rect 6546 11200 6552 11212
rect 5031 11172 6552 11200
rect 5031 11169 5043 11172
rect 4985 11163 5043 11169
rect 6546 11160 6552 11172
rect 6604 11200 6610 11212
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6604 11172 6929 11200
rect 6604 11160 6610 11172
rect 6917 11169 6929 11172
rect 6963 11200 6975 11203
rect 8202 11200 8208 11212
rect 6963 11172 8208 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 8202 11160 8208 11172
rect 8260 11200 8266 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8260 11172 8953 11200
rect 8260 11160 8266 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11200 9275 11203
rect 9766 11200 9772 11212
rect 9263 11172 9772 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 2038 11024 2044 11076
rect 2096 11024 2102 11076
rect 2774 11024 2780 11076
rect 2832 11024 2838 11076
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4120 11036 5750 11064
rect 4120 11024 4126 11036
rect 7190 11024 7196 11076
rect 7248 11024 7254 11076
rect 7650 11024 7656 11076
rect 7708 11024 7714 11076
rect 9674 11024 9680 11076
rect 9732 11024 9738 11076
rect 8570 10956 8576 11008
rect 8628 10996 8634 11008
rect 8665 10999 8723 11005
rect 8665 10996 8677 10999
rect 8628 10968 8677 10996
rect 8628 10956 8634 10968
rect 8665 10965 8677 10968
rect 8711 10965 8723 10999
rect 8665 10959 8723 10965
rect 1104 10906 11868 10928
rect 1104 10854 4894 10906
rect 4946 10854 4958 10906
rect 5010 10854 5022 10906
rect 5074 10854 5086 10906
rect 5138 10854 5150 10906
rect 5202 10854 6894 10906
rect 6946 10854 6958 10906
rect 7010 10854 7022 10906
rect 7074 10854 7086 10906
rect 7138 10854 7150 10906
rect 7202 10854 8894 10906
rect 8946 10854 8958 10906
rect 9010 10854 9022 10906
rect 9074 10854 9086 10906
rect 9138 10854 9150 10906
rect 9202 10854 10894 10906
rect 10946 10854 10958 10906
rect 11010 10854 11022 10906
rect 11074 10854 11086 10906
rect 11138 10854 11150 10906
rect 11202 10854 11868 10906
rect 1104 10832 11868 10854
rect 6779 10795 6837 10801
rect 6779 10792 6791 10795
rect 2424 10764 6791 10792
rect 2424 10733 2452 10764
rect 6779 10761 6791 10764
rect 6825 10761 6837 10795
rect 6779 10755 6837 10761
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 9674 10792 9680 10804
rect 7708 10764 9680 10792
rect 7708 10752 7714 10764
rect 2409 10727 2467 10733
rect 2409 10693 2421 10727
rect 2455 10693 2467 10727
rect 2409 10687 2467 10693
rect 2682 10684 2688 10736
rect 2740 10724 2746 10736
rect 8202 10724 8208 10736
rect 2740 10696 2898 10724
rect 8036 10696 8208 10724
rect 2740 10684 2746 10696
rect 5905 10659 5963 10665
rect 3804 10628 4554 10656
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 2179 10560 2268 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2240 10452 2268 10560
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 3142 10588 3148 10600
rect 2832 10560 3148 10588
rect 2832 10548 2838 10560
rect 3142 10548 3148 10560
rect 3200 10588 3206 10600
rect 3804 10588 3832 10628
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 6546 10656 6552 10668
rect 5951 10628 6552 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 6871 10659 6929 10665
rect 6871 10625 6883 10659
rect 6917 10656 6929 10659
rect 7282 10656 7288 10668
rect 6917 10628 7288 10656
rect 6917 10625 6929 10628
rect 6871 10619 6929 10625
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 8036 10665 8064 10696
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 8297 10727 8355 10733
rect 8297 10693 8309 10727
rect 8343 10724 8355 10727
rect 8570 10724 8576 10736
rect 8343 10696 8576 10724
rect 8343 10693 8355 10696
rect 8297 10687 8355 10693
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 8680 10724 8708 10764
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 9766 10752 9772 10804
rect 9824 10752 9830 10804
rect 9692 10724 9720 10752
rect 10134 10724 10140 10736
rect 8680 10696 8786 10724
rect 9692 10696 10140 10724
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 3200 10560 3832 10588
rect 3881 10591 3939 10597
rect 3200 10548 3206 10560
rect 3881 10557 3893 10591
rect 3927 10588 3939 10591
rect 5074 10588 5080 10600
rect 3927 10560 5080 10588
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 5074 10548 5080 10560
rect 5132 10588 5138 10600
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5132 10560 5641 10588
rect 5132 10548 5138 10560
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 3602 10452 3608 10464
rect 2240 10424 3608 10452
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4157 10455 4215 10461
rect 4157 10452 4169 10455
rect 4028 10424 4169 10452
rect 4028 10412 4034 10424
rect 4157 10421 4169 10424
rect 4203 10421 4215 10455
rect 4157 10415 4215 10421
rect 1104 10362 11868 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 6214 10362
rect 6266 10310 6278 10362
rect 6330 10310 6342 10362
rect 6394 10310 6406 10362
rect 6458 10310 6470 10362
rect 6522 10310 8214 10362
rect 8266 10310 8278 10362
rect 8330 10310 8342 10362
rect 8394 10310 8406 10362
rect 8458 10310 8470 10362
rect 8522 10310 10214 10362
rect 10266 10310 10278 10362
rect 10330 10310 10342 10362
rect 10394 10310 10406 10362
rect 10458 10310 10470 10362
rect 10522 10310 11868 10362
rect 1104 10288 11868 10310
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 2038 10248 2044 10260
rect 1903 10220 2044 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 6546 10248 6552 10260
rect 6503 10220 6552 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 11149 10251 11207 10257
rect 11149 10217 11161 10251
rect 11195 10248 11207 10251
rect 11238 10248 11244 10260
rect 11195 10220 11244 10248
rect 11195 10217 11207 10220
rect 11149 10211 11207 10217
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 3970 10180 3976 10192
rect 3528 10152 3976 10180
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 3528 10112 3556 10152
rect 3970 10140 3976 10152
rect 4028 10140 4034 10192
rect 3375 10084 3556 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 3602 10072 3608 10124
rect 3660 10072 3666 10124
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10044 4767 10047
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 4755 10016 4997 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5074 10004 5080 10056
rect 5132 10004 5138 10056
rect 9398 10004 9404 10056
rect 9456 10004 9462 10056
rect 2682 9936 2688 9988
rect 2740 9936 2746 9988
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 7745 9979 7803 9985
rect 7745 9976 7757 9979
rect 7340 9948 7757 9976
rect 7340 9936 7346 9948
rect 7745 9945 7757 9948
rect 7791 9945 7803 9979
rect 7745 9939 7803 9945
rect 9677 9979 9735 9985
rect 9677 9945 9689 9979
rect 9723 9976 9735 9979
rect 9723 9948 9904 9976
rect 9723 9945 9735 9948
rect 9677 9939 9735 9945
rect 9876 9920 9904 9948
rect 10134 9936 10140 9988
rect 10192 9936 10198 9988
rect 4706 9868 4712 9920
rect 4764 9868 4770 9920
rect 9858 9868 9864 9920
rect 9916 9868 9922 9920
rect 1104 9818 11868 9840
rect 1104 9766 4894 9818
rect 4946 9766 4958 9818
rect 5010 9766 5022 9818
rect 5074 9766 5086 9818
rect 5138 9766 5150 9818
rect 5202 9766 6894 9818
rect 6946 9766 6958 9818
rect 7010 9766 7022 9818
rect 7074 9766 7086 9818
rect 7138 9766 7150 9818
rect 7202 9766 8894 9818
rect 8946 9766 8958 9818
rect 9010 9766 9022 9818
rect 9074 9766 9086 9818
rect 9138 9766 9150 9818
rect 9202 9766 10894 9818
rect 10946 9766 10958 9818
rect 11010 9766 11022 9818
rect 11074 9766 11086 9818
rect 11138 9766 11150 9818
rect 11202 9766 11868 9818
rect 1104 9744 11868 9766
rect 10134 9596 10140 9648
rect 10192 9596 10198 9648
rect 4706 9528 4712 9580
rect 4764 9528 4770 9580
rect 8202 9528 8208 9580
rect 8260 9528 8266 9580
rect 7834 9460 7840 9512
rect 7892 9460 7898 9512
rect 8662 9460 8668 9512
rect 8720 9500 8726 9512
rect 9398 9500 9404 9512
rect 8720 9472 9404 9500
rect 8720 9460 8726 9472
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 9766 9500 9772 9512
rect 9723 9472 9772 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 11330 9500 11336 9512
rect 11195 9472 11336 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 4798 9324 4804 9376
rect 4856 9324 4862 9376
rect 1104 9274 11868 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 6214 9274
rect 6266 9222 6278 9274
rect 6330 9222 6342 9274
rect 6394 9222 6406 9274
rect 6458 9222 6470 9274
rect 6522 9222 8214 9274
rect 8266 9222 8278 9274
rect 8330 9222 8342 9274
rect 8394 9222 8406 9274
rect 8458 9222 8470 9274
rect 8522 9222 10214 9274
rect 10266 9222 10278 9274
rect 10330 9222 10342 9274
rect 10394 9222 10406 9274
rect 10458 9222 10470 9274
rect 10522 9222 11868 9274
rect 1104 9200 11868 9222
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 2866 9160 2872 9172
rect 1535 9132 2872 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 3878 9120 3884 9172
rect 3936 9120 3942 9172
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 6825 9163 6883 9169
rect 6825 9160 6837 9163
rect 6788 9132 6837 9160
rect 6788 9120 6794 9132
rect 6825 9129 6837 9132
rect 6871 9129 6883 9163
rect 6825 9123 6883 9129
rect 10689 9163 10747 9169
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 10778 9160 10784 9172
rect 10735 9132 10784 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 8297 9027 8355 9033
rect 8297 9024 8309 9027
rect 7892 8996 8309 9024
rect 7892 8984 7898 8996
rect 8297 8993 8309 8996
rect 8343 8993 8355 9027
rect 8297 8987 8355 8993
rect 8662 8984 8668 9036
rect 8720 9024 8726 9036
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 8720 8996 8953 9024
rect 8720 8984 8726 8996
rect 8941 8993 8953 8996
rect 8987 8993 8999 9027
rect 8941 8987 8999 8993
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 3326 8956 3332 8968
rect 3283 8928 3332 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8956 5687 8959
rect 6546 8956 6552 8968
rect 5675 8928 6552 8956
rect 5675 8925 5687 8928
rect 5629 8919 5687 8925
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 8754 8956 8760 8968
rect 8619 8928 8760 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 10778 8916 10784 8968
rect 10836 8956 10842 8968
rect 10908 8959 10966 8965
rect 10908 8956 10920 8959
rect 10836 8928 10920 8956
rect 10836 8916 10842 8928
rect 10908 8925 10920 8928
rect 10954 8925 10966 8959
rect 10908 8919 10966 8925
rect 2498 8848 2504 8900
rect 2556 8848 2562 8900
rect 2961 8891 3019 8897
rect 2961 8857 2973 8891
rect 3007 8888 3019 8891
rect 3050 8888 3056 8900
rect 3007 8860 3056 8888
rect 3007 8857 3019 8860
rect 2961 8851 3019 8857
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 4798 8848 4804 8900
rect 4856 8848 4862 8900
rect 5353 8891 5411 8897
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 5442 8888 5448 8900
rect 5399 8860 5448 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 8018 8888 8024 8900
rect 7866 8860 8024 8888
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 9217 8891 9275 8897
rect 9217 8857 9229 8891
rect 9263 8857 9275 8891
rect 9217 8851 9275 8857
rect 9232 8820 9260 8851
rect 10226 8848 10232 8900
rect 10284 8848 10290 8900
rect 9398 8820 9404 8832
rect 9232 8792 9404 8820
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 10962 8780 10968 8832
rect 11020 8829 11026 8832
rect 11020 8823 11069 8829
rect 11020 8789 11023 8823
rect 11057 8789 11069 8823
rect 11020 8783 11069 8789
rect 11020 8780 11026 8783
rect 1104 8730 11868 8752
rect 1104 8678 4894 8730
rect 4946 8678 4958 8730
rect 5010 8678 5022 8730
rect 5074 8678 5086 8730
rect 5138 8678 5150 8730
rect 5202 8678 6894 8730
rect 6946 8678 6958 8730
rect 7010 8678 7022 8730
rect 7074 8678 7086 8730
rect 7138 8678 7150 8730
rect 7202 8678 8894 8730
rect 8946 8678 8958 8730
rect 9010 8678 9022 8730
rect 9074 8678 9086 8730
rect 9138 8678 9150 8730
rect 9202 8678 10894 8730
rect 10946 8678 10958 8730
rect 11010 8678 11022 8730
rect 11074 8678 11086 8730
rect 11138 8678 11150 8730
rect 11202 8678 11868 8730
rect 1104 8656 11868 8678
rect 1302 8576 1308 8628
rect 1360 8616 1366 8628
rect 3789 8619 3847 8625
rect 3789 8616 3801 8619
rect 1360 8588 3801 8616
rect 1360 8576 1366 8588
rect 3789 8585 3801 8588
rect 3835 8585 3847 8619
rect 3789 8579 3847 8585
rect 8110 8576 8116 8628
rect 8168 8576 8174 8628
rect 2498 8508 2504 8560
rect 2556 8508 2562 8560
rect 4798 8508 4804 8560
rect 4856 8508 4862 8560
rect 5261 8551 5319 8557
rect 5261 8517 5273 8551
rect 5307 8548 5319 8551
rect 5350 8548 5356 8560
rect 5307 8520 5356 8548
rect 5307 8517 5319 8520
rect 5261 8511 5319 8517
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 6641 8551 6699 8557
rect 6641 8548 6653 8551
rect 6052 8520 6653 8548
rect 6052 8508 6058 8520
rect 6641 8517 6653 8520
rect 6687 8517 6699 8551
rect 6641 8511 6699 8517
rect 7650 8508 7656 8560
rect 7708 8508 7714 8560
rect 9306 8440 9312 8492
rect 9364 8440 9370 8492
rect 1489 8415 1547 8421
rect 1489 8381 1501 8415
rect 1535 8412 1547 8415
rect 2590 8412 2596 8424
rect 1535 8384 2596 8412
rect 1535 8381 1547 8384
rect 1489 8375 1547 8381
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 2866 8372 2872 8424
rect 2924 8412 2930 8424
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2924 8384 2973 8412
rect 2924 8372 2930 8384
rect 2961 8381 2973 8384
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 3326 8412 3332 8424
rect 3283 8384 3332 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 3252 8276 3280 8375
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 5534 8372 5540 8424
rect 5592 8372 5598 8424
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8412 6423 8415
rect 6411 8384 6500 8412
rect 6411 8381 6423 8384
rect 6365 8375 6423 8381
rect 3602 8276 3608 8288
rect 3252 8248 3608 8276
rect 3602 8236 3608 8248
rect 3660 8276 3666 8288
rect 5902 8276 5908 8288
rect 3660 8248 5908 8276
rect 3660 8236 3666 8248
rect 5902 8236 5908 8248
rect 5960 8276 5966 8288
rect 6472 8276 6500 8384
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 8481 8415 8539 8421
rect 8481 8412 8493 8415
rect 7432 8384 8493 8412
rect 7432 8372 7438 8384
rect 8481 8381 8493 8384
rect 8527 8381 8539 8415
rect 8481 8375 8539 8381
rect 8662 8276 8668 8288
rect 5960 8248 8668 8276
rect 5960 8236 5966 8248
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 1104 8186 11868 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 6214 8186
rect 6266 8134 6278 8186
rect 6330 8134 6342 8186
rect 6394 8134 6406 8186
rect 6458 8134 6470 8186
rect 6522 8134 8214 8186
rect 8266 8134 8278 8186
rect 8330 8134 8342 8186
rect 8394 8134 8406 8186
rect 8458 8134 8470 8186
rect 8522 8134 10214 8186
rect 10266 8134 10278 8186
rect 10330 8134 10342 8186
rect 10394 8134 10406 8186
rect 10458 8134 10470 8186
rect 10522 8134 11868 8186
rect 1104 8112 11868 8134
rect 1857 8075 1915 8081
rect 1857 8041 1869 8075
rect 1903 8072 1915 8075
rect 3234 8072 3240 8084
rect 1903 8044 3240 8072
rect 1903 8041 1915 8044
rect 1857 8035 1915 8041
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 4062 8032 4068 8084
rect 4120 8032 4126 8084
rect 7653 8075 7711 8081
rect 7653 8041 7665 8075
rect 7699 8072 7711 8075
rect 9214 8072 9220 8084
rect 7699 8044 9220 8072
rect 7699 8041 7711 8044
rect 7653 8035 7711 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 3602 7896 3608 7948
rect 3660 7896 3666 7948
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 4120 7908 6193 7936
rect 4120 7896 4126 7908
rect 6181 7905 6193 7908
rect 6227 7905 6239 7939
rect 6181 7899 6239 7905
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 6328 7908 9229 7936
rect 6328 7896 6334 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 5902 7828 5908 7880
rect 5960 7828 5966 7880
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8720 7840 8953 7868
rect 8720 7828 8726 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 2682 7760 2688 7812
rect 2740 7760 2746 7812
rect 3329 7803 3387 7809
rect 3329 7769 3341 7803
rect 3375 7769 3387 7803
rect 3329 7763 3387 7769
rect 3344 7732 3372 7763
rect 4798 7760 4804 7812
rect 4856 7760 4862 7812
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 5537 7803 5595 7809
rect 5537 7800 5549 7803
rect 5500 7772 5549 7800
rect 5500 7760 5506 7772
rect 5537 7769 5549 7772
rect 5583 7800 5595 7803
rect 7650 7800 7656 7812
rect 5583 7772 5764 7800
rect 7406 7772 7656 7800
rect 5583 7769 5595 7772
rect 5537 7763 5595 7769
rect 5626 7732 5632 7744
rect 3344 7704 5632 7732
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 5736 7732 5764 7772
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 8757 7803 8815 7809
rect 8757 7769 8769 7803
rect 8803 7800 8815 7803
rect 9490 7800 9496 7812
rect 8803 7772 9496 7800
rect 8803 7769 8815 7772
rect 8757 7763 8815 7769
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 10226 7760 10232 7812
rect 10284 7760 10290 7812
rect 7834 7732 7840 7744
rect 5736 7704 7840 7732
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 1104 7642 11868 7664
rect 1104 7590 4894 7642
rect 4946 7590 4958 7642
rect 5010 7590 5022 7642
rect 5074 7590 5086 7642
rect 5138 7590 5150 7642
rect 5202 7590 6894 7642
rect 6946 7590 6958 7642
rect 7010 7590 7022 7642
rect 7074 7590 7086 7642
rect 7138 7590 7150 7642
rect 7202 7590 8894 7642
rect 8946 7590 8958 7642
rect 9010 7590 9022 7642
rect 9074 7590 9086 7642
rect 9138 7590 9150 7642
rect 9202 7590 10894 7642
rect 10946 7590 10958 7642
rect 11010 7590 11022 7642
rect 11074 7590 11086 7642
rect 11138 7590 11150 7642
rect 11202 7590 11868 7642
rect 1104 7568 11868 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3142 7528 3148 7540
rect 2740 7500 3148 7528
rect 2740 7488 2746 7500
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 6270 7528 6276 7540
rect 5316 7500 6276 7528
rect 5316 7488 5322 7500
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 7193 7531 7251 7537
rect 7193 7497 7205 7531
rect 7239 7528 7251 7531
rect 7282 7528 7288 7540
rect 7239 7500 7288 7528
rect 7239 7497 7251 7500
rect 7193 7491 7251 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 11330 7528 11336 7540
rect 8496 7500 11336 7528
rect 8496 7469 8524 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 8481 7463 8539 7469
rect 8481 7429 8493 7463
rect 8527 7429 8539 7463
rect 8481 7423 8539 7429
rect 10042 7420 10048 7472
rect 10100 7420 10106 7472
rect 6181 7395 6239 7401
rect 6181 7361 6193 7395
rect 6227 7392 6239 7395
rect 6546 7392 6552 7404
rect 6227 7364 6552 7392
rect 6227 7361 6239 7364
rect 6181 7355 6239 7361
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8076 7364 8769 7392
rect 8076 7352 8082 7364
rect 8757 7361 8769 7364
rect 8803 7392 8815 7395
rect 8846 7392 8852 7404
rect 8803 7364 8852 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7324 5871 7327
rect 8570 7324 8576 7336
rect 5859 7296 8576 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8720 7296 9045 7324
rect 8720 7284 8726 7296
rect 8956 7200 8984 7296
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 9306 7284 9312 7336
rect 9364 7284 9370 7336
rect 10594 7284 10600 7336
rect 10652 7324 10658 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 10652 7296 10793 7324
rect 10652 7284 10658 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 8938 7148 8944 7200
rect 8996 7148 9002 7200
rect 1104 7098 11868 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 6214 7098
rect 6266 7046 6278 7098
rect 6330 7046 6342 7098
rect 6394 7046 6406 7098
rect 6458 7046 6470 7098
rect 6522 7046 8214 7098
rect 8266 7046 8278 7098
rect 8330 7046 8342 7098
rect 8394 7046 8406 7098
rect 8458 7046 8470 7098
rect 8522 7046 10214 7098
rect 10266 7046 10278 7098
rect 10330 7046 10342 7098
rect 10394 7046 10406 7098
rect 10458 7046 10470 7098
rect 10522 7046 11868 7098
rect 1104 7024 11868 7046
rect 7742 6944 7748 6996
rect 7800 6993 7806 6996
rect 7800 6987 7815 6993
rect 7803 6953 7815 6987
rect 7800 6947 7815 6953
rect 8665 6987 8723 6993
rect 8665 6953 8677 6987
rect 8711 6984 8723 6987
rect 8938 6984 8944 6996
rect 8711 6956 8944 6984
rect 8711 6953 8723 6956
rect 8665 6947 8723 6953
rect 7800 6944 7806 6947
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 9940 6987 9998 6993
rect 9940 6953 9952 6987
rect 9986 6984 9998 6987
rect 10042 6984 10048 6996
rect 9986 6956 10048 6984
rect 9986 6953 9998 6956
rect 9940 6947 9998 6953
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 3878 6808 3884 6860
rect 3936 6808 3942 6860
rect 4798 6848 4804 6860
rect 4264 6820 4804 6848
rect 4264 6766 4292 6820
rect 4798 6808 4804 6820
rect 4856 6848 4862 6860
rect 5350 6848 5356 6860
rect 4856 6820 5356 6848
rect 4856 6808 4862 6820
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6273 6851 6331 6857
rect 6273 6848 6285 6851
rect 6144 6820 6285 6848
rect 6144 6808 6150 6820
rect 6273 6817 6285 6820
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 8297 6851 8355 6857
rect 8297 6817 8309 6851
rect 8343 6848 8355 6851
rect 8570 6848 8576 6860
rect 8343 6820 8576 6848
rect 8343 6817 8355 6820
rect 8297 6811 8355 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 8846 6848 8852 6860
rect 8680 6820 8852 6848
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6780 5687 6783
rect 5810 6780 5816 6792
rect 5675 6752 5816 6780
rect 5675 6749 5687 6752
rect 5629 6743 5687 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 8018 6740 8024 6792
rect 8076 6740 8082 6792
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6780 8539 6783
rect 8680 6780 8708 6820
rect 8846 6808 8852 6820
rect 8904 6848 8910 6860
rect 10686 6848 10692 6860
rect 8904 6820 10692 6848
rect 8904 6808 8910 6820
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 8527 6752 8708 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 8588 6724 8616 6752
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9548 6752 9689 6780
rect 9548 6740 9554 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 5353 6715 5411 6721
rect 5353 6681 5365 6715
rect 5399 6712 5411 6715
rect 5442 6712 5448 6724
rect 5399 6684 5448 6712
rect 5399 6681 5411 6684
rect 5353 6675 5411 6681
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 8570 6712 8576 6724
rect 7314 6684 8576 6712
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 10686 6672 10692 6724
rect 10744 6672 10750 6724
rect 11422 6604 11428 6656
rect 11480 6604 11486 6656
rect 1104 6554 11868 6576
rect 1104 6502 4894 6554
rect 4946 6502 4958 6554
rect 5010 6502 5022 6554
rect 5074 6502 5086 6554
rect 5138 6502 5150 6554
rect 5202 6502 6894 6554
rect 6946 6502 6958 6554
rect 7010 6502 7022 6554
rect 7074 6502 7086 6554
rect 7138 6502 7150 6554
rect 7202 6502 8894 6554
rect 8946 6502 8958 6554
rect 9010 6502 9022 6554
rect 9074 6502 9086 6554
rect 9138 6502 9150 6554
rect 9202 6502 10894 6554
rect 10946 6502 10958 6554
rect 11010 6502 11022 6554
rect 11074 6502 11086 6554
rect 11138 6502 11150 6554
rect 11202 6502 11868 6554
rect 1104 6480 11868 6502
rect 1210 6400 1216 6452
rect 1268 6440 1274 6452
rect 2041 6443 2099 6449
rect 2041 6440 2053 6443
rect 1268 6412 2053 6440
rect 1268 6400 1274 6412
rect 2041 6409 2053 6412
rect 2087 6409 2099 6443
rect 2041 6403 2099 6409
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 4614 6440 4620 6452
rect 4479 6412 4620 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 6546 6400 6552 6452
rect 6604 6440 6610 6452
rect 8662 6440 8668 6452
rect 6604 6412 8668 6440
rect 6604 6400 6610 6412
rect 2498 6332 2504 6384
rect 2556 6332 2562 6384
rect 3513 6375 3571 6381
rect 3513 6341 3525 6375
rect 3559 6372 3571 6375
rect 3559 6344 4660 6372
rect 3559 6341 3571 6344
rect 3513 6335 3571 6341
rect 4632 6316 4660 6344
rect 5350 6332 5356 6384
rect 5408 6332 5414 6384
rect 4614 6264 4620 6316
rect 4672 6304 4678 6316
rect 7024 6313 7052 6412
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 7190 6332 7196 6384
rect 7248 6372 7254 6384
rect 7285 6375 7343 6381
rect 7285 6372 7297 6375
rect 7248 6344 7297 6372
rect 7248 6332 7254 6344
rect 7285 6341 7297 6344
rect 7331 6372 7343 6375
rect 7374 6372 7380 6384
rect 7331 6344 7380 6372
rect 7331 6341 7343 6344
rect 7285 6335 7343 6341
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 8570 6372 8576 6384
rect 8510 6344 8576 6372
rect 8570 6332 8576 6344
rect 8628 6332 8634 6384
rect 10778 6332 10784 6384
rect 10836 6332 10842 6384
rect 7009 6307 7067 6313
rect 4672 6276 4752 6304
rect 4672 6264 4678 6276
rect 3786 6196 3792 6248
rect 3844 6196 3850 6248
rect 4724 6236 4752 6276
rect 7009 6273 7021 6307
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 5442 6236 5448 6248
rect 4724 6208 5448 6236
rect 5442 6196 5448 6208
rect 5500 6236 5506 6248
rect 5905 6239 5963 6245
rect 5905 6236 5917 6239
rect 5500 6208 5917 6236
rect 5500 6196 5506 6208
rect 5905 6205 5917 6208
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6236 6239 6239
rect 6730 6236 6736 6248
rect 6227 6208 6736 6236
rect 6227 6205 6239 6208
rect 6181 6199 6239 6205
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7374 6236 7380 6248
rect 6972 6208 7380 6236
rect 6972 6196 6978 6208
rect 7374 6196 7380 6208
rect 7432 6236 7438 6248
rect 8018 6236 8024 6248
rect 7432 6208 8024 6236
rect 7432 6196 7438 6208
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 9490 6196 9496 6248
rect 9548 6196 9554 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9600 6208 9781 6236
rect 9600 6168 9628 6208
rect 9769 6205 9781 6208
rect 9815 6236 9827 6239
rect 11422 6236 11428 6248
rect 9815 6208 11428 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 11422 6196 11428 6208
rect 11480 6196 11486 6248
rect 8312 6140 9628 6168
rect 6546 6060 6552 6112
rect 6604 6100 6610 6112
rect 8312 6100 8340 6140
rect 6604 6072 8340 6100
rect 6604 6060 6610 6072
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8628 6072 8769 6100
rect 8628 6060 8634 6072
rect 8757 6069 8769 6072
rect 8803 6100 8815 6103
rect 9766 6100 9772 6112
rect 8803 6072 9772 6100
rect 8803 6069 8815 6072
rect 8757 6063 8815 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 11241 6103 11299 6109
rect 11241 6069 11253 6103
rect 11287 6100 11299 6103
rect 11422 6100 11428 6112
rect 11287 6072 11428 6100
rect 11287 6069 11299 6072
rect 11241 6063 11299 6069
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 1104 6010 11868 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 6214 6010
rect 6266 5958 6278 6010
rect 6330 5958 6342 6010
rect 6394 5958 6406 6010
rect 6458 5958 6470 6010
rect 6522 5958 8214 6010
rect 8266 5958 8278 6010
rect 8330 5958 8342 6010
rect 8394 5958 8406 6010
rect 8458 5958 8470 6010
rect 8522 5958 10214 6010
rect 10266 5958 10278 6010
rect 10330 5958 10342 6010
rect 10394 5958 10406 6010
rect 10458 5958 10470 6010
rect 10522 5958 11868 6010
rect 1104 5936 11868 5958
rect 1857 5899 1915 5905
rect 1857 5865 1869 5899
rect 1903 5896 1915 5899
rect 2774 5896 2780 5908
rect 1903 5868 2780 5896
rect 1903 5865 1915 5868
rect 1857 5859 1915 5865
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 3786 5896 3792 5908
rect 3568 5868 3792 5896
rect 3568 5856 3574 5868
rect 3786 5856 3792 5868
rect 3844 5896 3850 5908
rect 3844 5868 7052 5896
rect 3844 5856 3850 5868
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5760 3387 5763
rect 4614 5760 4620 5772
rect 3375 5732 4620 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 6546 5720 6552 5772
rect 6604 5720 6610 5772
rect 7024 5760 7052 5868
rect 9861 5763 9919 5769
rect 9861 5760 9873 5763
rect 7024 5732 9873 5760
rect 9861 5729 9873 5732
rect 9907 5760 9919 5763
rect 11422 5760 11428 5772
rect 9907 5732 11428 5760
rect 9907 5729 9919 5732
rect 9861 5723 9919 5729
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 3694 5692 3700 5704
rect 3651 5664 3700 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 4798 5652 4804 5704
rect 4856 5692 4862 5704
rect 4856 5664 5198 5692
rect 4856 5652 4862 5664
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 9585 5695 9643 5701
rect 9585 5692 9597 5695
rect 9548 5664 9597 5692
rect 9548 5652 9554 5664
rect 9585 5661 9597 5664
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 10928 5664 10994 5692
rect 10928 5652 10934 5664
rect 2682 5584 2688 5636
rect 2740 5584 2746 5636
rect 6273 5627 6331 5633
rect 6273 5593 6285 5627
rect 6319 5624 6331 5627
rect 7190 5624 7196 5636
rect 6319 5596 7196 5624
rect 6319 5593 6331 5596
rect 6273 5587 6331 5593
rect 7190 5584 7196 5596
rect 7248 5624 7254 5636
rect 7466 5624 7472 5636
rect 7248 5596 7472 5624
rect 7248 5584 7254 5596
rect 7466 5584 7472 5596
rect 7524 5584 7530 5636
rect 8418 5596 9996 5624
rect 4801 5559 4859 5565
rect 4801 5525 4813 5559
rect 4847 5556 4859 5559
rect 5626 5556 5632 5568
rect 4847 5528 5632 5556
rect 4847 5525 4859 5528
rect 4801 5519 4859 5525
rect 5626 5516 5632 5528
rect 5684 5556 5690 5568
rect 6086 5556 6092 5568
rect 5684 5528 6092 5556
rect 5684 5516 5690 5528
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 8665 5559 8723 5565
rect 8665 5556 8677 5559
rect 8536 5528 8677 5556
rect 8536 5516 8542 5528
rect 8665 5525 8677 5528
rect 8711 5556 8723 5559
rect 9858 5556 9864 5568
rect 8711 5528 9864 5556
rect 8711 5525 8723 5528
rect 8665 5519 8723 5525
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 9968 5556 9996 5596
rect 10686 5556 10692 5568
rect 9968 5528 10692 5556
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 11330 5516 11336 5568
rect 11388 5516 11394 5568
rect 1104 5466 11868 5488
rect 1104 5414 4894 5466
rect 4946 5414 4958 5466
rect 5010 5414 5022 5466
rect 5074 5414 5086 5466
rect 5138 5414 5150 5466
rect 5202 5414 6894 5466
rect 6946 5414 6958 5466
rect 7010 5414 7022 5466
rect 7074 5414 7086 5466
rect 7138 5414 7150 5466
rect 7202 5414 8894 5466
rect 8946 5414 8958 5466
rect 9010 5414 9022 5466
rect 9074 5414 9086 5466
rect 9138 5414 9150 5466
rect 9202 5414 10894 5466
rect 10946 5414 10958 5466
rect 11010 5414 11022 5466
rect 11074 5414 11086 5466
rect 11138 5414 11150 5466
rect 11202 5414 11868 5466
rect 1104 5392 11868 5414
rect 3602 5312 3608 5364
rect 3660 5312 3666 5364
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 9674 5352 9680 5364
rect 3752 5324 9680 5352
rect 3752 5312 3758 5324
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 2682 5244 2688 5296
rect 2740 5284 2746 5296
rect 4798 5284 4804 5296
rect 2740 5256 3832 5284
rect 4646 5256 4804 5284
rect 2740 5244 2746 5256
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5216 3479 5219
rect 3510 5216 3516 5228
rect 3467 5188 3516 5216
rect 3467 5185 3479 5188
rect 3421 5179 3479 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 3142 5108 3148 5160
rect 3200 5108 3206 5160
rect 1673 5015 1731 5021
rect 1673 4981 1685 5015
rect 1719 5012 1731 5015
rect 3050 5012 3056 5024
rect 1719 4984 3056 5012
rect 1719 4981 1731 4984
rect 1673 4975 1731 4981
rect 3050 4972 3056 4984
rect 3108 4972 3114 5024
rect 3804 5012 3832 5256
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 5077 5287 5135 5293
rect 5077 5253 5089 5287
rect 5123 5284 5135 5287
rect 5442 5284 5448 5296
rect 5123 5256 5448 5284
rect 5123 5253 5135 5256
rect 5077 5247 5135 5253
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 7282 5244 7288 5296
rect 7340 5284 7346 5296
rect 7561 5287 7619 5293
rect 7561 5284 7573 5287
rect 7340 5256 7573 5284
rect 7340 5244 7346 5256
rect 7561 5253 7573 5256
rect 7607 5253 7619 5287
rect 7561 5247 7619 5253
rect 10686 5244 10692 5296
rect 10744 5244 10750 5296
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5216 5411 5219
rect 6546 5216 6552 5228
rect 5399 5188 6552 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5117 9459 5151
rect 9401 5111 9459 5117
rect 4890 5012 4896 5024
rect 3804 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 9033 5015 9091 5021
rect 9033 4981 9045 5015
rect 9079 5012 9091 5015
rect 9416 5012 9444 5111
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 11330 5148 11336 5160
rect 9732 5120 11336 5148
rect 9732 5108 9738 5120
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 9490 5012 9496 5024
rect 9079 4984 9496 5012
rect 9079 4981 9091 4984
rect 9033 4975 9091 4981
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 11149 5015 11207 5021
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11238 5012 11244 5024
rect 11195 4984 11244 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 1104 4922 11868 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 6214 4922
rect 6266 4870 6278 4922
rect 6330 4870 6342 4922
rect 6394 4870 6406 4922
rect 6458 4870 6470 4922
rect 6522 4870 8214 4922
rect 8266 4870 8278 4922
rect 8330 4870 8342 4922
rect 8394 4870 8406 4922
rect 8458 4870 8470 4922
rect 8522 4870 10214 4922
rect 10266 4870 10278 4922
rect 10330 4870 10342 4922
rect 10394 4870 10406 4922
rect 10458 4870 10470 4922
rect 10522 4870 11868 4922
rect 1104 4848 11868 4870
rect 3142 4768 3148 4820
rect 3200 4808 3206 4820
rect 3200 4780 3556 4808
rect 3200 4768 3206 4780
rect 3528 4740 3556 4780
rect 3878 4768 3884 4820
rect 3936 4808 3942 4820
rect 4062 4808 4068 4820
rect 3936 4780 4068 4808
rect 3936 4768 3942 4780
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 4614 4808 4620 4820
rect 4356 4780 4620 4808
rect 4356 4740 4384 4780
rect 4614 4768 4620 4780
rect 4672 4808 4678 4820
rect 5371 4811 5429 4817
rect 5371 4808 5383 4811
rect 4672 4780 5383 4808
rect 4672 4768 4678 4780
rect 5371 4777 5383 4780
rect 5417 4808 5429 4811
rect 6996 4811 7054 4817
rect 6996 4808 7008 4811
rect 5417 4780 7008 4808
rect 5417 4777 5429 4780
rect 5371 4771 5429 4777
rect 6996 4777 7008 4780
rect 7042 4808 7054 4811
rect 7466 4808 7472 4820
rect 7042 4780 7472 4808
rect 7042 4777 7054 4780
rect 6996 4771 7054 4777
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 5810 4740 5816 4752
rect 3528 4712 4384 4740
rect 5644 4712 5816 4740
rect 3329 4675 3387 4681
rect 3329 4641 3341 4675
rect 3375 4672 3387 4675
rect 3528 4672 3556 4712
rect 3375 4644 3556 4672
rect 3605 4675 3663 4681
rect 3375 4641 3387 4644
rect 3329 4635 3387 4641
rect 3605 4641 3617 4675
rect 3651 4672 3663 4675
rect 3694 4672 3700 4684
rect 3651 4644 3700 4672
rect 3651 4641 3663 4644
rect 3605 4635 3663 4641
rect 3694 4632 3700 4644
rect 3752 4632 3758 4684
rect 5644 4681 5672 4712
rect 5810 4700 5816 4712
rect 5868 4740 5874 4752
rect 5868 4712 6868 4740
rect 5868 4700 5874 4712
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4641 5687 4675
rect 5629 4635 5687 4641
rect 6730 4632 6736 4684
rect 6788 4632 6794 4684
rect 6840 4672 6868 4712
rect 9766 4672 9772 4684
rect 6840 4644 9772 4672
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 2590 4496 2596 4548
rect 2648 4496 2654 4548
rect 4890 4496 4896 4548
rect 4948 4536 4954 4548
rect 5442 4536 5448 4548
rect 4948 4508 5448 4536
rect 4948 4496 4954 4508
rect 5442 4496 5448 4508
rect 5500 4496 5506 4548
rect 8294 4536 8300 4548
rect 8234 4508 8300 4536
rect 8294 4496 8300 4508
rect 8352 4496 8358 4548
rect 1857 4471 1915 4477
rect 1857 4437 1869 4471
rect 1903 4468 1915 4471
rect 2682 4468 2688 4480
rect 1903 4440 2688 4468
rect 1903 4437 1915 4440
rect 1857 4431 1915 4437
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 8478 4428 8484 4480
rect 8536 4468 8542 4480
rect 9398 4468 9404 4480
rect 8536 4440 9404 4468
rect 8536 4428 8542 4440
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 1104 4378 11868 4400
rect 1104 4326 4894 4378
rect 4946 4326 4958 4378
rect 5010 4326 5022 4378
rect 5074 4326 5086 4378
rect 5138 4326 5150 4378
rect 5202 4326 6894 4378
rect 6946 4326 6958 4378
rect 7010 4326 7022 4378
rect 7074 4326 7086 4378
rect 7138 4326 7150 4378
rect 7202 4326 8894 4378
rect 8946 4326 8958 4378
rect 9010 4326 9022 4378
rect 9074 4326 9086 4378
rect 9138 4326 9150 4378
rect 9202 4326 10894 4378
rect 10946 4326 10958 4378
rect 11010 4326 11022 4378
rect 11074 4326 11086 4378
rect 11138 4326 11150 4378
rect 11202 4326 11868 4378
rect 1104 4304 11868 4326
rect 5442 4224 5448 4276
rect 5500 4264 5506 4276
rect 8294 4264 8300 4276
rect 5500 4236 5672 4264
rect 5500 4224 5506 4236
rect 4525 4199 4583 4205
rect 4525 4165 4537 4199
rect 4571 4196 4583 4199
rect 4614 4196 4620 4208
rect 4571 4168 4620 4196
rect 4571 4165 4583 4168
rect 4525 4159 4583 4165
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 5644 4128 5672 4236
rect 6932 4236 8300 4264
rect 6932 4128 6960 4236
rect 8294 4224 8300 4236
rect 8352 4264 8358 4276
rect 10686 4264 10692 4276
rect 8352 4236 10692 4264
rect 8352 4224 8358 4236
rect 7466 4156 7472 4208
rect 7524 4156 7530 4208
rect 8772 4196 8800 4236
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 11238 4196 11244 4208
rect 8694 4168 8800 4196
rect 11072 4168 11244 4196
rect 5644 4114 6960 4128
rect 5658 4100 6960 4114
rect 10778 4088 10784 4140
rect 10836 4128 10842 4140
rect 11072 4128 11100 4168
rect 11238 4156 11244 4168
rect 11296 4156 11302 4208
rect 10836 4100 10902 4128
rect 10980 4100 11100 4128
rect 10836 4088 10842 4100
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4060 4307 4063
rect 5534 4060 5540 4072
rect 4295 4032 5540 4060
rect 4295 4029 4307 4032
rect 4249 4023 4307 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 5994 4060 6000 4072
rect 5868 4032 6000 4060
rect 5868 4020 5874 4032
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 5552 3992 5580 4020
rect 6822 3992 6828 4004
rect 5552 3964 6828 3992
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 7208 3924 7236 4023
rect 9490 4020 9496 4072
rect 9548 4020 9554 4072
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 10980 4060 11008 4100
rect 9824 4032 11008 4060
rect 9824 4020 9830 4032
rect 8754 3924 8760 3936
rect 7208 3896 8760 3924
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9306 3924 9312 3936
rect 8996 3896 9312 3924
rect 8996 3884 9002 3896
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 11238 3884 11244 3936
rect 11296 3884 11302 3936
rect 1104 3834 11868 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 6214 3834
rect 6266 3782 6278 3834
rect 6330 3782 6342 3834
rect 6394 3782 6406 3834
rect 6458 3782 6470 3834
rect 6522 3782 8214 3834
rect 8266 3782 8278 3834
rect 8330 3782 8342 3834
rect 8394 3782 8406 3834
rect 8458 3782 8470 3834
rect 8522 3782 10214 3834
rect 10266 3782 10278 3834
rect 10330 3782 10342 3834
rect 10394 3782 10406 3834
rect 10458 3782 10470 3834
rect 10522 3782 11868 3834
rect 1104 3760 11868 3782
rect 6730 3680 6736 3732
rect 6788 3680 6794 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 6880 3692 8800 3720
rect 6880 3680 6886 3692
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6748 3584 6776 3680
rect 8772 3652 8800 3692
rect 8772 3624 9720 3652
rect 6595 3556 6776 3584
rect 6825 3587 6883 3593
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 6871 3556 6929 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 6917 3553 6929 3556
rect 6963 3584 6975 3587
rect 8570 3584 8576 3596
rect 6963 3556 8576 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 8570 3544 8576 3556
rect 8628 3584 8634 3596
rect 9490 3584 9496 3596
rect 8628 3556 9496 3584
rect 8628 3544 8634 3556
rect 9490 3544 9496 3556
rect 9548 3584 9554 3596
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 9548 3556 9597 3584
rect 9548 3544 9554 3556
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9692 3584 9720 3624
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9692 3556 9873 3584
rect 9585 3547 9643 3553
rect 9861 3553 9873 3556
rect 9907 3584 9919 3587
rect 11238 3584 11244 3596
rect 9907 3556 11244 3584
rect 9907 3553 9919 3556
rect 9861 3547 9919 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 5442 3476 5448 3528
rect 5500 3476 5506 3528
rect 7180 3451 7238 3457
rect 7180 3448 7192 3451
rect 7116 3420 7192 3448
rect 5077 3383 5135 3389
rect 5077 3349 5089 3383
rect 5123 3380 5135 3383
rect 7116 3380 7144 3420
rect 7180 3417 7192 3420
rect 7226 3448 7238 3451
rect 7282 3448 7288 3460
rect 7226 3420 7288 3448
rect 7226 3417 7238 3420
rect 7180 3411 7238 3417
rect 7282 3408 7288 3420
rect 7340 3408 7346 3460
rect 8418 3420 9352 3448
rect 5123 3352 7144 3380
rect 5123 3349 5135 3352
rect 5077 3343 5135 3349
rect 7834 3340 7840 3392
rect 7892 3380 7898 3392
rect 8496 3380 8524 3420
rect 7892 3352 8524 3380
rect 7892 3340 7898 3352
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 9214 3380 9220 3392
rect 8720 3352 9220 3380
rect 8720 3340 8726 3352
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 9324 3380 9352 3420
rect 10870 3408 10876 3460
rect 10928 3408 10934 3460
rect 10778 3380 10784 3392
rect 9324 3352 10784 3380
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 11330 3340 11336 3392
rect 11388 3340 11394 3392
rect 1104 3290 11868 3312
rect 1104 3238 4894 3290
rect 4946 3238 4958 3290
rect 5010 3238 5022 3290
rect 5074 3238 5086 3290
rect 5138 3238 5150 3290
rect 5202 3238 6894 3290
rect 6946 3238 6958 3290
rect 7010 3238 7022 3290
rect 7074 3238 7086 3290
rect 7138 3238 7150 3290
rect 7202 3238 8894 3290
rect 8946 3238 8958 3290
rect 9010 3238 9022 3290
rect 9074 3238 9086 3290
rect 9138 3238 9150 3290
rect 9202 3238 10894 3290
rect 10946 3238 10958 3290
rect 11010 3238 11022 3290
rect 11074 3238 11086 3290
rect 11138 3238 11150 3290
rect 11202 3238 11868 3290
rect 1104 3216 11868 3238
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 5258 3176 5264 3188
rect 4488 3148 5264 3176
rect 4488 3136 4494 3148
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 6788 3148 6837 3176
rect 6788 3136 6794 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 11241 3179 11299 3185
rect 11241 3176 11253 3179
rect 6825 3139 6883 3145
rect 8772 3148 11253 3176
rect 8772 3120 8800 3148
rect 11241 3145 11253 3148
rect 11287 3176 11299 3179
rect 11422 3176 11428 3188
rect 11287 3148 11428 3176
rect 11287 3145 11299 3148
rect 11241 3139 11299 3145
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 5442 3068 5448 3120
rect 5500 3068 5506 3120
rect 5902 3068 5908 3120
rect 5960 3108 5966 3120
rect 5960 3080 6224 3108
rect 5960 3068 5966 3080
rect 6196 3049 6224 3080
rect 7834 3068 7840 3120
rect 7892 3068 7898 3120
rect 8297 3111 8355 3117
rect 8297 3077 8309 3111
rect 8343 3108 8355 3111
rect 8754 3108 8760 3120
rect 8343 3080 8760 3108
rect 8343 3077 8355 3080
rect 8297 3071 8355 3077
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 10778 3068 10784 3120
rect 10836 3068 10842 3120
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 5905 2975 5963 2981
rect 5905 2972 5917 2975
rect 4672 2944 5917 2972
rect 4672 2932 4678 2944
rect 5905 2941 5917 2944
rect 5951 2941 5963 2975
rect 6196 2972 6224 3003
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 8628 3012 9505 3040
rect 8628 3000 8634 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 6196 2944 9781 2972
rect 5905 2935 5963 2941
rect 9769 2941 9781 2944
rect 9815 2972 9827 2975
rect 11330 2972 11336 2984
rect 9815 2944 11336 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 1104 2746 11868 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 6214 2746
rect 6266 2694 6278 2746
rect 6330 2694 6342 2746
rect 6394 2694 6406 2746
rect 6458 2694 6470 2746
rect 6522 2694 8214 2746
rect 8266 2694 8278 2746
rect 8330 2694 8342 2746
rect 8394 2694 8406 2746
rect 8458 2694 8470 2746
rect 8522 2694 10214 2746
rect 10266 2694 10278 2746
rect 10330 2694 10342 2746
rect 10394 2694 10406 2746
rect 10458 2694 10470 2746
rect 10522 2694 11868 2746
rect 1104 2672 11868 2694
rect 1104 2202 11868 2224
rect 1104 2150 4894 2202
rect 4946 2150 4958 2202
rect 5010 2150 5022 2202
rect 5074 2150 5086 2202
rect 5138 2150 5150 2202
rect 5202 2150 6894 2202
rect 6946 2150 6958 2202
rect 7010 2150 7022 2202
rect 7074 2150 7086 2202
rect 7138 2150 7150 2202
rect 7202 2150 8894 2202
rect 8946 2150 8958 2202
rect 9010 2150 9022 2202
rect 9074 2150 9086 2202
rect 9138 2150 9150 2202
rect 9202 2150 10894 2202
rect 10946 2150 10958 2202
rect 11010 2150 11022 2202
rect 11074 2150 11086 2202
rect 11138 2150 11150 2202
rect 11202 2150 11868 2202
rect 1104 2128 11868 2150
<< via1 >>
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 6214 12486 6266 12538
rect 6278 12486 6330 12538
rect 6342 12486 6394 12538
rect 6406 12486 6458 12538
rect 6470 12486 6522 12538
rect 8214 12486 8266 12538
rect 8278 12486 8330 12538
rect 8342 12486 8394 12538
rect 8406 12486 8458 12538
rect 8470 12486 8522 12538
rect 10214 12486 10266 12538
rect 10278 12486 10330 12538
rect 10342 12486 10394 12538
rect 10406 12486 10458 12538
rect 10470 12486 10522 12538
rect 3608 12180 3660 12232
rect 4160 12155 4212 12164
rect 4160 12121 4169 12155
rect 4169 12121 4203 12155
rect 4203 12121 4212 12155
rect 4160 12112 4212 12121
rect 2780 12044 2832 12096
rect 4068 12044 4120 12096
rect 5908 12044 5960 12096
rect 4894 11942 4946 11994
rect 4958 11942 5010 11994
rect 5022 11942 5074 11994
rect 5086 11942 5138 11994
rect 5150 11942 5202 11994
rect 6894 11942 6946 11994
rect 6958 11942 7010 11994
rect 7022 11942 7074 11994
rect 7086 11942 7138 11994
rect 7150 11942 7202 11994
rect 8894 11942 8946 11994
rect 8958 11942 9010 11994
rect 9022 11942 9074 11994
rect 9086 11942 9138 11994
rect 9150 11942 9202 11994
rect 10894 11942 10946 11994
rect 10958 11942 11010 11994
rect 11022 11942 11074 11994
rect 11086 11942 11138 11994
rect 11150 11942 11202 11994
rect 3608 11840 3660 11892
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 4160 11840 4212 11849
rect 2780 11772 2832 11824
rect 4068 11772 4120 11824
rect 5908 11815 5960 11824
rect 5908 11781 5917 11815
rect 5917 11781 5951 11815
rect 5951 11781 5960 11815
rect 5908 11772 5960 11781
rect 7656 11840 7708 11892
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 6460 11679 6512 11688
rect 6460 11645 6469 11679
rect 6469 11645 6503 11679
rect 6503 11645 6512 11679
rect 6460 11636 6512 11645
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 4896 11500 4948 11552
rect 7196 11500 7248 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 6214 11398 6266 11450
rect 6278 11398 6330 11450
rect 6342 11398 6394 11450
rect 6406 11398 6458 11450
rect 6470 11398 6522 11450
rect 8214 11398 8266 11450
rect 8278 11398 8330 11450
rect 8342 11398 8394 11450
rect 8406 11398 8458 11450
rect 8470 11398 8522 11450
rect 10214 11398 10266 11450
rect 10278 11398 10330 11450
rect 10342 11398 10394 11450
rect 10406 11398 10458 11450
rect 10470 11398 10522 11450
rect 2688 11296 2740 11348
rect 4896 11296 4948 11348
rect 6736 11339 6788 11348
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 7288 11296 7340 11348
rect 3608 11160 3660 11212
rect 6552 11160 6604 11212
rect 8208 11160 8260 11212
rect 9772 11160 9824 11212
rect 2044 11067 2096 11076
rect 2044 11033 2053 11067
rect 2053 11033 2087 11067
rect 2087 11033 2096 11067
rect 2044 11024 2096 11033
rect 2780 11024 2832 11076
rect 4068 11024 4120 11076
rect 7196 11067 7248 11076
rect 7196 11033 7205 11067
rect 7205 11033 7239 11067
rect 7239 11033 7248 11067
rect 7196 11024 7248 11033
rect 7656 11024 7708 11076
rect 9680 11024 9732 11076
rect 8576 10956 8628 11008
rect 4894 10854 4946 10906
rect 4958 10854 5010 10906
rect 5022 10854 5074 10906
rect 5086 10854 5138 10906
rect 5150 10854 5202 10906
rect 6894 10854 6946 10906
rect 6958 10854 7010 10906
rect 7022 10854 7074 10906
rect 7086 10854 7138 10906
rect 7150 10854 7202 10906
rect 8894 10854 8946 10906
rect 8958 10854 9010 10906
rect 9022 10854 9074 10906
rect 9086 10854 9138 10906
rect 9150 10854 9202 10906
rect 10894 10854 10946 10906
rect 10958 10854 11010 10906
rect 11022 10854 11074 10906
rect 11086 10854 11138 10906
rect 11150 10854 11202 10906
rect 7656 10752 7708 10804
rect 2688 10684 2740 10736
rect 2780 10548 2832 10600
rect 3148 10548 3200 10600
rect 6552 10616 6604 10668
rect 7288 10616 7340 10668
rect 8208 10684 8260 10736
rect 8576 10684 8628 10736
rect 9680 10752 9732 10804
rect 9772 10795 9824 10804
rect 9772 10761 9781 10795
rect 9781 10761 9815 10795
rect 9815 10761 9824 10795
rect 9772 10752 9824 10761
rect 10140 10684 10192 10736
rect 5080 10548 5132 10600
rect 3608 10412 3660 10464
rect 3976 10412 4028 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 6214 10310 6266 10362
rect 6278 10310 6330 10362
rect 6342 10310 6394 10362
rect 6406 10310 6458 10362
rect 6470 10310 6522 10362
rect 8214 10310 8266 10362
rect 8278 10310 8330 10362
rect 8342 10310 8394 10362
rect 8406 10310 8458 10362
rect 8470 10310 8522 10362
rect 10214 10310 10266 10362
rect 10278 10310 10330 10362
rect 10342 10310 10394 10362
rect 10406 10310 10458 10362
rect 10470 10310 10522 10362
rect 2044 10208 2096 10260
rect 6552 10208 6604 10260
rect 11244 10208 11296 10260
rect 3976 10140 4028 10192
rect 3608 10115 3660 10124
rect 3608 10081 3617 10115
rect 3617 10081 3651 10115
rect 3651 10081 3660 10115
rect 3608 10072 3660 10081
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 2688 9936 2740 9988
rect 7288 9936 7340 9988
rect 10140 9936 10192 9988
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 9864 9868 9916 9920
rect 4894 9766 4946 9818
rect 4958 9766 5010 9818
rect 5022 9766 5074 9818
rect 5086 9766 5138 9818
rect 5150 9766 5202 9818
rect 6894 9766 6946 9818
rect 6958 9766 7010 9818
rect 7022 9766 7074 9818
rect 7086 9766 7138 9818
rect 7150 9766 7202 9818
rect 8894 9766 8946 9818
rect 8958 9766 9010 9818
rect 9022 9766 9074 9818
rect 9086 9766 9138 9818
rect 9150 9766 9202 9818
rect 10894 9766 10946 9818
rect 10958 9766 11010 9818
rect 11022 9766 11074 9818
rect 11086 9766 11138 9818
rect 11150 9766 11202 9818
rect 10140 9596 10192 9648
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 7840 9503 7892 9512
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 8668 9460 8720 9512
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 9772 9460 9824 9512
rect 11336 9460 11388 9512
rect 4804 9367 4856 9376
rect 4804 9333 4813 9367
rect 4813 9333 4847 9367
rect 4847 9333 4856 9367
rect 4804 9324 4856 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 6214 9222 6266 9274
rect 6278 9222 6330 9274
rect 6342 9222 6394 9274
rect 6406 9222 6458 9274
rect 6470 9222 6522 9274
rect 8214 9222 8266 9274
rect 8278 9222 8330 9274
rect 8342 9222 8394 9274
rect 8406 9222 8458 9274
rect 8470 9222 8522 9274
rect 10214 9222 10266 9274
rect 10278 9222 10330 9274
rect 10342 9222 10394 9274
rect 10406 9222 10458 9274
rect 10470 9222 10522 9274
rect 2872 9120 2924 9172
rect 3884 9163 3936 9172
rect 3884 9129 3893 9163
rect 3893 9129 3927 9163
rect 3927 9129 3936 9163
rect 3884 9120 3936 9129
rect 6736 9120 6788 9172
rect 10784 9120 10836 9172
rect 7840 8984 7892 9036
rect 8668 8984 8720 9036
rect 3332 8916 3384 8968
rect 6552 8916 6604 8968
rect 8760 8916 8812 8968
rect 10784 8916 10836 8968
rect 2504 8848 2556 8900
rect 3056 8848 3108 8900
rect 4804 8848 4856 8900
rect 5448 8848 5500 8900
rect 8024 8848 8076 8900
rect 10232 8848 10284 8900
rect 9404 8780 9456 8832
rect 10968 8780 11020 8832
rect 4894 8678 4946 8730
rect 4958 8678 5010 8730
rect 5022 8678 5074 8730
rect 5086 8678 5138 8730
rect 5150 8678 5202 8730
rect 6894 8678 6946 8730
rect 6958 8678 7010 8730
rect 7022 8678 7074 8730
rect 7086 8678 7138 8730
rect 7150 8678 7202 8730
rect 8894 8678 8946 8730
rect 8958 8678 9010 8730
rect 9022 8678 9074 8730
rect 9086 8678 9138 8730
rect 9150 8678 9202 8730
rect 10894 8678 10946 8730
rect 10958 8678 11010 8730
rect 11022 8678 11074 8730
rect 11086 8678 11138 8730
rect 11150 8678 11202 8730
rect 1308 8576 1360 8628
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 2504 8508 2556 8560
rect 4804 8508 4856 8560
rect 5356 8508 5408 8560
rect 6000 8508 6052 8560
rect 7656 8508 7708 8560
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 2596 8372 2648 8424
rect 2872 8372 2924 8424
rect 3332 8372 3384 8424
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 3608 8236 3660 8288
rect 5908 8236 5960 8288
rect 7380 8372 7432 8424
rect 8668 8236 8720 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 6214 8134 6266 8186
rect 6278 8134 6330 8186
rect 6342 8134 6394 8186
rect 6406 8134 6458 8186
rect 6470 8134 6522 8186
rect 8214 8134 8266 8186
rect 8278 8134 8330 8186
rect 8342 8134 8394 8186
rect 8406 8134 8458 8186
rect 8470 8134 8522 8186
rect 10214 8134 10266 8186
rect 10278 8134 10330 8186
rect 10342 8134 10394 8186
rect 10406 8134 10458 8186
rect 10470 8134 10522 8186
rect 3240 8032 3292 8084
rect 4068 8075 4120 8084
rect 4068 8041 4077 8075
rect 4077 8041 4111 8075
rect 4111 8041 4120 8075
rect 4068 8032 4120 8041
rect 9220 8032 9272 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 3608 7939 3660 7948
rect 3608 7905 3617 7939
rect 3617 7905 3651 7939
rect 3651 7905 3660 7939
rect 3608 7896 3660 7905
rect 4068 7896 4120 7948
rect 6276 7896 6328 7948
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 8668 7828 8720 7880
rect 2688 7760 2740 7812
rect 4804 7760 4856 7812
rect 5448 7760 5500 7812
rect 5632 7692 5684 7744
rect 7656 7760 7708 7812
rect 9496 7760 9548 7812
rect 10232 7760 10284 7812
rect 7840 7692 7892 7744
rect 4894 7590 4946 7642
rect 4958 7590 5010 7642
rect 5022 7590 5074 7642
rect 5086 7590 5138 7642
rect 5150 7590 5202 7642
rect 6894 7590 6946 7642
rect 6958 7590 7010 7642
rect 7022 7590 7074 7642
rect 7086 7590 7138 7642
rect 7150 7590 7202 7642
rect 8894 7590 8946 7642
rect 8958 7590 9010 7642
rect 9022 7590 9074 7642
rect 9086 7590 9138 7642
rect 9150 7590 9202 7642
rect 10894 7590 10946 7642
rect 10958 7590 11010 7642
rect 11022 7590 11074 7642
rect 11086 7590 11138 7642
rect 11150 7590 11202 7642
rect 2688 7488 2740 7540
rect 3148 7488 3200 7540
rect 5264 7488 5316 7540
rect 6276 7488 6328 7540
rect 7288 7488 7340 7540
rect 11336 7488 11388 7540
rect 10048 7420 10100 7472
rect 6552 7352 6604 7404
rect 8024 7352 8076 7404
rect 8852 7352 8904 7404
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 8668 7284 8720 7336
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 10600 7284 10652 7336
rect 8944 7191 8996 7200
rect 8944 7157 8953 7191
rect 8953 7157 8987 7191
rect 8987 7157 8996 7191
rect 8944 7148 8996 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 6214 7046 6266 7098
rect 6278 7046 6330 7098
rect 6342 7046 6394 7098
rect 6406 7046 6458 7098
rect 6470 7046 6522 7098
rect 8214 7046 8266 7098
rect 8278 7046 8330 7098
rect 8342 7046 8394 7098
rect 8406 7046 8458 7098
rect 8470 7046 8522 7098
rect 10214 7046 10266 7098
rect 10278 7046 10330 7098
rect 10342 7046 10394 7098
rect 10406 7046 10458 7098
rect 10470 7046 10522 7098
rect 7748 6987 7800 6996
rect 7748 6953 7769 6987
rect 7769 6953 7800 6987
rect 7748 6944 7800 6953
rect 8944 6944 8996 6996
rect 10048 6944 10100 6996
rect 3884 6851 3936 6860
rect 3884 6817 3893 6851
rect 3893 6817 3927 6851
rect 3927 6817 3936 6851
rect 3884 6808 3936 6817
rect 4804 6808 4856 6860
rect 5356 6808 5408 6860
rect 6092 6808 6144 6860
rect 8576 6808 8628 6860
rect 5816 6740 5868 6792
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8852 6808 8904 6860
rect 10692 6808 10744 6860
rect 9496 6740 9548 6792
rect 5448 6672 5500 6724
rect 8576 6672 8628 6724
rect 10692 6672 10744 6724
rect 11428 6647 11480 6656
rect 11428 6613 11437 6647
rect 11437 6613 11471 6647
rect 11471 6613 11480 6647
rect 11428 6604 11480 6613
rect 4894 6502 4946 6554
rect 4958 6502 5010 6554
rect 5022 6502 5074 6554
rect 5086 6502 5138 6554
rect 5150 6502 5202 6554
rect 6894 6502 6946 6554
rect 6958 6502 7010 6554
rect 7022 6502 7074 6554
rect 7086 6502 7138 6554
rect 7150 6502 7202 6554
rect 8894 6502 8946 6554
rect 8958 6502 9010 6554
rect 9022 6502 9074 6554
rect 9086 6502 9138 6554
rect 9150 6502 9202 6554
rect 10894 6502 10946 6554
rect 10958 6502 11010 6554
rect 11022 6502 11074 6554
rect 11086 6502 11138 6554
rect 11150 6502 11202 6554
rect 1216 6400 1268 6452
rect 4620 6400 4672 6452
rect 6552 6400 6604 6452
rect 2504 6332 2556 6384
rect 5356 6332 5408 6384
rect 4620 6264 4672 6316
rect 8668 6400 8720 6452
rect 7196 6332 7248 6384
rect 7380 6332 7432 6384
rect 8576 6332 8628 6384
rect 10784 6332 10836 6384
rect 3792 6239 3844 6248
rect 3792 6205 3801 6239
rect 3801 6205 3835 6239
rect 3835 6205 3844 6239
rect 3792 6196 3844 6205
rect 5448 6196 5500 6248
rect 6736 6196 6788 6248
rect 6920 6196 6972 6248
rect 7380 6196 7432 6248
rect 8024 6196 8076 6248
rect 9496 6239 9548 6248
rect 9496 6205 9505 6239
rect 9505 6205 9539 6239
rect 9539 6205 9548 6239
rect 9496 6196 9548 6205
rect 11428 6196 11480 6248
rect 6552 6060 6604 6112
rect 8576 6060 8628 6112
rect 9772 6060 9824 6112
rect 11428 6060 11480 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 6214 5958 6266 6010
rect 6278 5958 6330 6010
rect 6342 5958 6394 6010
rect 6406 5958 6458 6010
rect 6470 5958 6522 6010
rect 8214 5958 8266 6010
rect 8278 5958 8330 6010
rect 8342 5958 8394 6010
rect 8406 5958 8458 6010
rect 8470 5958 8522 6010
rect 10214 5958 10266 6010
rect 10278 5958 10330 6010
rect 10342 5958 10394 6010
rect 10406 5958 10458 6010
rect 10470 5958 10522 6010
rect 2780 5856 2832 5908
rect 3516 5856 3568 5908
rect 3792 5856 3844 5908
rect 4620 5720 4672 5772
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 11428 5720 11480 5772
rect 3700 5652 3752 5704
rect 4804 5652 4856 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 9496 5652 9548 5704
rect 10876 5652 10928 5704
rect 2688 5584 2740 5636
rect 7196 5627 7248 5636
rect 7196 5593 7205 5627
rect 7205 5593 7239 5627
rect 7239 5593 7248 5627
rect 7196 5584 7248 5593
rect 7472 5584 7524 5636
rect 5632 5516 5684 5568
rect 6092 5516 6144 5568
rect 8484 5516 8536 5568
rect 9864 5516 9916 5568
rect 10692 5516 10744 5568
rect 11336 5559 11388 5568
rect 11336 5525 11345 5559
rect 11345 5525 11379 5559
rect 11379 5525 11388 5559
rect 11336 5516 11388 5525
rect 4894 5414 4946 5466
rect 4958 5414 5010 5466
rect 5022 5414 5074 5466
rect 5086 5414 5138 5466
rect 5150 5414 5202 5466
rect 6894 5414 6946 5466
rect 6958 5414 7010 5466
rect 7022 5414 7074 5466
rect 7086 5414 7138 5466
rect 7150 5414 7202 5466
rect 8894 5414 8946 5466
rect 8958 5414 9010 5466
rect 9022 5414 9074 5466
rect 9086 5414 9138 5466
rect 9150 5414 9202 5466
rect 10894 5414 10946 5466
rect 10958 5414 11010 5466
rect 11022 5414 11074 5466
rect 11086 5414 11138 5466
rect 11150 5414 11202 5466
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 3700 5312 3752 5364
rect 9680 5312 9732 5364
rect 2688 5244 2740 5296
rect 3516 5176 3568 5228
rect 3148 5151 3200 5160
rect 3148 5117 3157 5151
rect 3157 5117 3191 5151
rect 3191 5117 3200 5151
rect 3148 5108 3200 5117
rect 3056 4972 3108 5024
rect 4804 5244 4856 5296
rect 5448 5244 5500 5296
rect 7288 5244 7340 5296
rect 10692 5244 10744 5296
rect 6552 5176 6604 5228
rect 4896 4972 4948 5024
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 11336 5108 11388 5160
rect 9496 4972 9548 5024
rect 11244 4972 11296 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 6214 4870 6266 4922
rect 6278 4870 6330 4922
rect 6342 4870 6394 4922
rect 6406 4870 6458 4922
rect 6470 4870 6522 4922
rect 8214 4870 8266 4922
rect 8278 4870 8330 4922
rect 8342 4870 8394 4922
rect 8406 4870 8458 4922
rect 8470 4870 8522 4922
rect 10214 4870 10266 4922
rect 10278 4870 10330 4922
rect 10342 4870 10394 4922
rect 10406 4870 10458 4922
rect 10470 4870 10522 4922
rect 3148 4768 3200 4820
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 4068 4768 4120 4820
rect 4620 4768 4672 4820
rect 7472 4768 7524 4820
rect 3700 4632 3752 4684
rect 5816 4700 5868 4752
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 9772 4632 9824 4684
rect 2596 4496 2648 4548
rect 4896 4496 4948 4548
rect 5448 4496 5500 4548
rect 8300 4496 8352 4548
rect 2688 4428 2740 4480
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 8484 4428 8536 4437
rect 9404 4428 9456 4480
rect 4894 4326 4946 4378
rect 4958 4326 5010 4378
rect 5022 4326 5074 4378
rect 5086 4326 5138 4378
rect 5150 4326 5202 4378
rect 6894 4326 6946 4378
rect 6958 4326 7010 4378
rect 7022 4326 7074 4378
rect 7086 4326 7138 4378
rect 7150 4326 7202 4378
rect 8894 4326 8946 4378
rect 8958 4326 9010 4378
rect 9022 4326 9074 4378
rect 9086 4326 9138 4378
rect 9150 4326 9202 4378
rect 10894 4326 10946 4378
rect 10958 4326 11010 4378
rect 11022 4326 11074 4378
rect 11086 4326 11138 4378
rect 11150 4326 11202 4378
rect 5448 4224 5500 4276
rect 4620 4156 4672 4208
rect 8300 4224 8352 4276
rect 7472 4199 7524 4208
rect 7472 4165 7481 4199
rect 7481 4165 7515 4199
rect 7515 4165 7524 4199
rect 7472 4156 7524 4165
rect 10692 4224 10744 4276
rect 10784 4088 10836 4140
rect 11244 4156 11296 4208
rect 5540 4020 5592 4072
rect 5816 4020 5868 4072
rect 6000 4063 6052 4072
rect 6000 4029 6009 4063
rect 6009 4029 6043 4063
rect 6043 4029 6052 4063
rect 6000 4020 6052 4029
rect 6828 3952 6880 4004
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 8760 3884 8812 3936
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 8944 3884 8996 3893
rect 9312 3884 9364 3936
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 6214 3782 6266 3834
rect 6278 3782 6330 3834
rect 6342 3782 6394 3834
rect 6406 3782 6458 3834
rect 6470 3782 6522 3834
rect 8214 3782 8266 3834
rect 8278 3782 8330 3834
rect 8342 3782 8394 3834
rect 8406 3782 8458 3834
rect 8470 3782 8522 3834
rect 10214 3782 10266 3834
rect 10278 3782 10330 3834
rect 10342 3782 10394 3834
rect 10406 3782 10458 3834
rect 10470 3782 10522 3834
rect 6736 3680 6788 3732
rect 6828 3680 6880 3732
rect 8576 3544 8628 3596
rect 9496 3544 9548 3596
rect 11244 3544 11296 3596
rect 5448 3476 5500 3528
rect 7288 3408 7340 3460
rect 7840 3340 7892 3392
rect 8668 3383 8720 3392
rect 8668 3349 8677 3383
rect 8677 3349 8711 3383
rect 8711 3349 8720 3383
rect 8668 3340 8720 3349
rect 9220 3340 9272 3392
rect 10876 3408 10928 3460
rect 10784 3340 10836 3392
rect 11336 3383 11388 3392
rect 11336 3349 11345 3383
rect 11345 3349 11379 3383
rect 11379 3349 11388 3383
rect 11336 3340 11388 3349
rect 4894 3238 4946 3290
rect 4958 3238 5010 3290
rect 5022 3238 5074 3290
rect 5086 3238 5138 3290
rect 5150 3238 5202 3290
rect 6894 3238 6946 3290
rect 6958 3238 7010 3290
rect 7022 3238 7074 3290
rect 7086 3238 7138 3290
rect 7150 3238 7202 3290
rect 8894 3238 8946 3290
rect 8958 3238 9010 3290
rect 9022 3238 9074 3290
rect 9086 3238 9138 3290
rect 9150 3238 9202 3290
rect 10894 3238 10946 3290
rect 10958 3238 11010 3290
rect 11022 3238 11074 3290
rect 11086 3238 11138 3290
rect 11150 3238 11202 3290
rect 4436 3179 4488 3188
rect 4436 3145 4445 3179
rect 4445 3145 4479 3179
rect 4479 3145 4488 3179
rect 4436 3136 4488 3145
rect 5264 3136 5316 3188
rect 6736 3136 6788 3188
rect 11428 3136 11480 3188
rect 5448 3068 5500 3120
rect 5908 3068 5960 3120
rect 7840 3068 7892 3120
rect 8760 3068 8812 3120
rect 10784 3068 10836 3120
rect 4620 2932 4672 2984
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 11336 2932 11388 2984
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 6214 2694 6266 2746
rect 6278 2694 6330 2746
rect 6342 2694 6394 2746
rect 6406 2694 6458 2746
rect 6470 2694 6522 2746
rect 8214 2694 8266 2746
rect 8278 2694 8330 2746
rect 8342 2694 8394 2746
rect 8406 2694 8458 2746
rect 8470 2694 8522 2746
rect 10214 2694 10266 2746
rect 10278 2694 10330 2746
rect 10342 2694 10394 2746
rect 10406 2694 10458 2746
rect 10470 2694 10522 2746
rect 4894 2150 4946 2202
rect 4958 2150 5010 2202
rect 5022 2150 5074 2202
rect 5086 2150 5138 2202
rect 5150 2150 5202 2202
rect 6894 2150 6946 2202
rect 6958 2150 7010 2202
rect 7022 2150 7074 2202
rect 7086 2150 7138 2202
rect 7150 2150 7202 2202
rect 8894 2150 8946 2202
rect 8958 2150 9010 2202
rect 9022 2150 9074 2202
rect 9086 2150 9138 2202
rect 9150 2150 9202 2202
rect 10894 2150 10946 2202
rect 10958 2150 11010 2202
rect 11022 2150 11074 2202
rect 11086 2150 11138 2202
rect 11150 2150 11202 2202
<< metal2 >>
rect 2962 15056 3018 15065
rect 2962 14991 3018 15000
rect 9218 15056 9274 15065
rect 9218 14991 9274 15000
rect 2870 14376 2926 14385
rect 2870 14311 2926 14320
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 2792 12102 2820 12951
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2792 11830 2820 12038
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2700 11354 2728 11630
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2792 11082 2820 11766
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2056 10266 2084 11018
rect 2792 10826 2820 11018
rect 2700 10798 2820 10826
rect 2700 10742 2728 10798
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2700 9994 2728 10678
rect 2792 10606 2820 10798
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2884 9178 2912 14311
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 1306 8936 1362 8945
rect 1306 8871 1362 8880
rect 2504 8900 2556 8906
rect 1320 8634 1348 8871
rect 2504 8842 2556 8848
rect 1308 8628 1360 8634
rect 1308 8570 1360 8576
rect 2516 8566 2544 8842
rect 2976 8650 3004 14991
rect 8114 14376 8170 14385
rect 8114 14311 8170 14320
rect 3146 13696 3202 13705
rect 3146 13631 3202 13640
rect 3160 12434 3188 13631
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 6214 12540 6522 12549
rect 6214 12538 6220 12540
rect 6276 12538 6300 12540
rect 6356 12538 6380 12540
rect 6436 12538 6460 12540
rect 6516 12538 6522 12540
rect 6276 12486 6278 12538
rect 6458 12486 6460 12538
rect 6214 12484 6220 12486
rect 6276 12484 6300 12486
rect 6356 12484 6380 12486
rect 6436 12484 6460 12486
rect 6516 12484 6522 12486
rect 6214 12475 6522 12484
rect 3160 12406 3280 12434
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2792 8622 3004 8650
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2516 8242 2544 8502
rect 2596 8424 2648 8430
rect 2792 8378 2820 8622
rect 2648 8372 2820 8378
rect 2596 8366 2820 8372
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2608 8350 2820 8366
rect 2516 8214 2728 8242
rect 2700 7818 2728 8214
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2700 7546 2728 7754
rect 2778 7576 2834 7585
rect 2688 7540 2740 7546
rect 2778 7511 2834 7520
rect 2688 7482 2740 7488
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1228 6458 1256 6831
rect 1216 6452 1268 6458
rect 1216 6394 1268 6400
rect 2504 6384 2556 6390
rect 2504 6326 2556 6332
rect 2516 5624 2544 6326
rect 2792 5914 2820 7511
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2688 5636 2740 5642
rect 2516 5596 2688 5624
rect 2688 5578 2740 5584
rect 2700 5302 2728 5578
rect 2688 5296 2740 5302
rect 2608 5256 2688 5284
rect 2608 4554 2636 5256
rect 2688 5238 2740 5244
rect 2596 4548 2648 4554
rect 2596 4490 2648 4496
rect 2688 4480 2740 4486
rect 2884 4434 2912 8366
rect 3068 5030 3096 8842
rect 3160 7546 3188 10542
rect 3252 8090 3280 12406
rect 3882 12336 3938 12345
rect 3882 12271 3938 12280
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3620 11898 3648 12174
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3620 11218 3648 11834
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3620 10470 3648 11154
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3620 10130 3648 10406
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3896 9178 3924 12271
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11830 4108 12038
rect 4172 11898 4200 12106
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 4894 11996 5202 12005
rect 4894 11994 4900 11996
rect 4956 11994 4980 11996
rect 5036 11994 5060 11996
rect 5116 11994 5140 11996
rect 5196 11994 5202 11996
rect 4956 11942 4958 11994
rect 5138 11942 5140 11994
rect 4894 11940 4900 11942
rect 4956 11940 4980 11942
rect 5036 11940 5060 11942
rect 5116 11940 5140 11942
rect 5196 11940 5202 11942
rect 4894 11931 5202 11940
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 5920 11830 5948 12038
rect 6894 11996 7202 12005
rect 6894 11994 6900 11996
rect 6956 11994 6980 11996
rect 7036 11994 7060 11996
rect 7116 11994 7140 11996
rect 7196 11994 7202 11996
rect 6956 11942 6958 11994
rect 7138 11942 7140 11994
rect 6894 11940 6900 11942
rect 6956 11940 6980 11942
rect 7036 11940 7060 11942
rect 7116 11940 7140 11942
rect 7196 11940 7202 11942
rect 6894 11931 7202 11940
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 4080 11082 4108 11766
rect 6460 11688 6512 11694
rect 6090 11656 6146 11665
rect 6736 11688 6788 11694
rect 6512 11648 6592 11676
rect 6460 11630 6512 11636
rect 6090 11591 6146 11600
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4908 11354 4936 11494
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4618 10976 4674 10985
rect 4618 10911 4674 10920
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10198 4016 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 4066 9616 4122 9625
rect 4066 9551 4122 9560
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3344 8430 3372 8910
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3882 8256 3938 8265
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3620 7954 3648 8230
rect 3882 8191 3938 8200
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3896 6866 3924 8191
rect 4080 8090 4108 9551
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3792 6248 3844 6254
rect 3606 6216 3662 6225
rect 3792 6190 3844 6196
rect 3606 6151 3662 6160
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3528 5234 3556 5850
rect 3620 5370 3648 6151
rect 3804 5914 3832 6190
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3712 5370 3740 5646
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2740 4428 2912 4434
rect 2688 4422 2912 4428
rect 2700 4406 2912 4422
rect 2792 785 2820 4406
rect 3068 2774 3096 4966
rect 3160 4826 3188 5102
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3712 4690 3740 5306
rect 4080 4826 4108 7890
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6458 4660 10911
rect 4894 10908 5202 10917
rect 4894 10906 4900 10908
rect 4956 10906 4980 10908
rect 5036 10906 5060 10908
rect 5116 10906 5140 10908
rect 5196 10906 5202 10908
rect 4956 10854 4958 10906
rect 5138 10854 5140 10906
rect 4894 10852 4900 10854
rect 4956 10852 4980 10854
rect 5036 10852 5060 10854
rect 5116 10852 5140 10854
rect 5196 10852 5202 10854
rect 4894 10843 5202 10852
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5092 10062 5120 10542
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9586 4752 9862
rect 4894 9820 5202 9829
rect 4894 9818 4900 9820
rect 4956 9818 4980 9820
rect 5036 9818 5060 9820
rect 5116 9818 5140 9820
rect 5196 9818 5202 9820
rect 4956 9766 4958 9818
rect 5138 9766 5140 9818
rect 4894 9764 4900 9766
rect 4956 9764 4980 9766
rect 5036 9764 5060 9766
rect 5116 9764 5140 9766
rect 5196 9764 5202 9766
rect 4894 9755 5202 9764
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4816 8906 4844 9318
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 4816 8566 4844 8842
rect 4894 8732 5202 8741
rect 4894 8730 4900 8732
rect 4956 8730 4980 8732
rect 5036 8730 5060 8732
rect 5116 8730 5140 8732
rect 5196 8730 5202 8732
rect 4956 8678 4958 8730
rect 5138 8678 5140 8730
rect 4894 8676 4900 8678
rect 4956 8676 4980 8678
rect 5036 8676 5060 8678
rect 5116 8676 5140 8678
rect 5196 8676 5202 8678
rect 4894 8667 5202 8676
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 5356 8560 5408 8566
rect 5460 8548 5488 8842
rect 5408 8520 5488 8548
rect 5356 8502 5408 8508
rect 4816 7818 4844 8502
rect 5460 7818 5488 8520
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 4816 6866 4844 7754
rect 4894 7644 5202 7653
rect 4894 7642 4900 7644
rect 4956 7642 4980 7644
rect 5036 7642 5060 7644
rect 5116 7642 5140 7644
rect 5196 7642 5202 7644
rect 4956 7590 4958 7642
rect 5138 7590 5140 7642
rect 4894 7588 4900 7590
rect 4956 7588 4980 7590
rect 5036 7588 5060 7590
rect 5116 7588 5140 7590
rect 5196 7588 5202 7590
rect 4894 7579 5202 7588
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4894 6556 5202 6565
rect 4894 6554 4900 6556
rect 4956 6554 4980 6556
rect 5036 6554 5060 6556
rect 5116 6554 5140 6556
rect 5196 6554 5202 6556
rect 4956 6502 4958 6554
rect 5138 6502 5140 6554
rect 4894 6500 4900 6502
rect 4956 6500 4980 6502
rect 5036 6500 5060 6502
rect 5116 6500 5140 6502
rect 5196 6500 5202 6502
rect 4894 6491 5202 6500
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5778 4660 6258
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 5302 4844 5646
rect 4894 5468 5202 5477
rect 4894 5466 4900 5468
rect 4956 5466 4980 5468
rect 5036 5466 5060 5468
rect 5116 5466 5140 5468
rect 5196 5466 5202 5468
rect 4956 5414 4958 5466
rect 5138 5414 5140 5466
rect 4894 5412 4900 5414
rect 4956 5412 4980 5414
rect 5036 5412 5060 5414
rect 5116 5412 5140 5414
rect 5196 5412 5202 5414
rect 4894 5403 5202 5412
rect 4804 5296 4856 5302
rect 4856 5256 4936 5284
rect 4804 5238 4856 5244
rect 4908 5030 4936 5256
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 2976 2746 3096 2774
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 2976 105 3004 2746
rect 3896 1465 3924 4762
rect 4632 4214 4660 4762
rect 4908 4554 4936 4966
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4894 4380 5202 4389
rect 4894 4378 4900 4380
rect 4956 4378 4980 4380
rect 5036 4378 5060 4380
rect 5116 4378 5140 4380
rect 5196 4378 5202 4380
rect 4956 4326 4958 4378
rect 5138 4326 5140 4378
rect 4894 4324 4900 4326
rect 4956 4324 4980 4326
rect 5036 4324 5060 4326
rect 5116 4324 5140 4326
rect 5196 4324 5202 4326
rect 4894 4315 5202 4324
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4448 2961 4476 3130
rect 4632 2990 4660 4150
rect 4894 3292 5202 3301
rect 4894 3290 4900 3292
rect 4956 3290 4980 3292
rect 5036 3290 5060 3292
rect 5116 3290 5140 3292
rect 5196 3290 5202 3292
rect 4956 3238 4958 3290
rect 5138 3238 5140 3290
rect 4894 3236 4900 3238
rect 4956 3236 4980 3238
rect 5036 3236 5060 3238
rect 5116 3236 5140 3238
rect 5196 3236 5202 3238
rect 4894 3227 5202 3236
rect 5276 3194 5304 7482
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5368 6390 5396 6802
rect 5460 6730 5488 7754
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5368 4536 5396 6326
rect 5460 6254 5488 6666
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5460 5302 5488 6190
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5448 4548 5500 4554
rect 5368 4508 5448 4536
rect 5448 4490 5500 4496
rect 5460 4282 5488 4490
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5460 3534 5488 4218
rect 5552 4078 5580 8366
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 7886 5948 8230
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 5574 5672 7686
rect 5828 6882 5856 7822
rect 5828 6854 5948 6882
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5828 4758 5856 6734
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5460 3126 5488 3470
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 4620 2984 4672 2990
rect 4434 2952 4490 2961
rect 4620 2926 4672 2932
rect 4434 2887 4490 2896
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5828 2417 5856 4014
rect 5920 3126 5948 6854
rect 6012 4078 6040 8502
rect 6104 6866 6132 11591
rect 6214 11452 6522 11461
rect 6214 11450 6220 11452
rect 6276 11450 6300 11452
rect 6356 11450 6380 11452
rect 6436 11450 6460 11452
rect 6516 11450 6522 11452
rect 6276 11398 6278 11450
rect 6458 11398 6460 11450
rect 6214 11396 6220 11398
rect 6276 11396 6300 11398
rect 6356 11396 6380 11398
rect 6436 11396 6460 11398
rect 6516 11396 6522 11398
rect 6214 11387 6522 11396
rect 6564 11218 6592 11648
rect 6736 11630 6788 11636
rect 6748 11354 6776 11630
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 10674 6592 11154
rect 7208 11082 7236 11494
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 6894 10908 7202 10917
rect 6894 10906 6900 10908
rect 6956 10906 6980 10908
rect 7036 10906 7060 10908
rect 7116 10906 7140 10908
rect 7196 10906 7202 10908
rect 6956 10854 6958 10906
rect 7138 10854 7140 10906
rect 6894 10852 6900 10854
rect 6956 10852 6980 10854
rect 7036 10852 7060 10854
rect 7116 10852 7140 10854
rect 7196 10852 7202 10854
rect 6894 10843 7202 10852
rect 7300 10674 7328 11290
rect 7668 11082 7696 11834
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7668 10810 7696 11018
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 6214 10364 6522 10373
rect 6214 10362 6220 10364
rect 6276 10362 6300 10364
rect 6356 10362 6380 10364
rect 6436 10362 6460 10364
rect 6516 10362 6522 10364
rect 6276 10310 6278 10362
rect 6458 10310 6460 10362
rect 6214 10308 6220 10310
rect 6276 10308 6300 10310
rect 6356 10308 6380 10310
rect 6436 10308 6460 10310
rect 6516 10308 6522 10310
rect 6214 10299 6522 10308
rect 6564 10266 6592 10610
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6734 10160 6790 10169
rect 6734 10095 6790 10104
rect 6214 9276 6522 9285
rect 6214 9274 6220 9276
rect 6276 9274 6300 9276
rect 6356 9274 6380 9276
rect 6436 9274 6460 9276
rect 6516 9274 6522 9276
rect 6276 9222 6278 9274
rect 6458 9222 6460 9274
rect 6214 9220 6220 9222
rect 6276 9220 6300 9222
rect 6356 9220 6380 9222
rect 6436 9220 6460 9222
rect 6516 9220 6522 9222
rect 6214 9211 6522 9220
rect 6748 9178 6776 10095
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 6894 9820 7202 9829
rect 6894 9818 6900 9820
rect 6956 9818 6980 9820
rect 7036 9818 7060 9820
rect 7116 9818 7140 9820
rect 7196 9818 7202 9820
rect 6956 9766 6958 9818
rect 7138 9766 7140 9818
rect 6894 9764 6900 9766
rect 6956 9764 6980 9766
rect 7036 9764 7060 9766
rect 7116 9764 7140 9766
rect 7196 9764 7202 9766
rect 6894 9755 7202 9764
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6214 8188 6522 8197
rect 6214 8186 6220 8188
rect 6276 8186 6300 8188
rect 6356 8186 6380 8188
rect 6436 8186 6460 8188
rect 6516 8186 6522 8188
rect 6276 8134 6278 8186
rect 6458 8134 6460 8186
rect 6214 8132 6220 8134
rect 6276 8132 6300 8134
rect 6356 8132 6380 8134
rect 6436 8132 6460 8134
rect 6516 8132 6522 8134
rect 6214 8123 6522 8132
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6288 7546 6316 7890
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6564 7410 6592 8910
rect 6894 8732 7202 8741
rect 6894 8730 6900 8732
rect 6956 8730 6980 8732
rect 7036 8730 7060 8732
rect 7116 8730 7140 8732
rect 7196 8730 7202 8732
rect 6956 8678 6958 8730
rect 7138 8678 7140 8730
rect 6894 8676 6900 8678
rect 6956 8676 6980 8678
rect 7036 8676 7060 8678
rect 7116 8676 7140 8678
rect 7196 8676 7202 8678
rect 6894 8667 7202 8676
rect 6894 7644 7202 7653
rect 6894 7642 6900 7644
rect 6956 7642 6980 7644
rect 7036 7642 7060 7644
rect 7116 7642 7140 7644
rect 7196 7642 7202 7644
rect 6956 7590 6958 7642
rect 7138 7590 7140 7642
rect 6894 7588 6900 7590
rect 6956 7588 6980 7590
rect 7036 7588 7060 7590
rect 7116 7588 7140 7590
rect 7196 7588 7202 7590
rect 6894 7579 7202 7588
rect 7300 7546 7328 9930
rect 7668 8566 7696 10746
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7852 9042 7880 9454
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6214 7100 6522 7109
rect 6214 7098 6220 7100
rect 6276 7098 6300 7100
rect 6356 7098 6380 7100
rect 6436 7098 6460 7100
rect 6516 7098 6522 7100
rect 6276 7046 6278 7098
rect 6458 7046 6460 7098
rect 6214 7044 6220 7046
rect 6276 7044 6300 7046
rect 6356 7044 6380 7046
rect 6436 7044 6460 7046
rect 6516 7044 6522 7046
rect 6214 7035 6522 7044
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6564 6458 6592 7346
rect 6894 6556 7202 6565
rect 6894 6554 6900 6556
rect 6956 6554 6980 6556
rect 7036 6554 7060 6556
rect 7116 6554 7140 6556
rect 7196 6554 7202 6556
rect 6956 6502 6958 6554
rect 7138 6502 7140 6554
rect 6894 6500 6900 6502
rect 6956 6500 6980 6502
rect 7036 6500 7060 6502
rect 7116 6500 7140 6502
rect 7196 6500 7202 6502
rect 6894 6491 7202 6500
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6214 6012 6522 6021
rect 6214 6010 6220 6012
rect 6276 6010 6300 6012
rect 6356 6010 6380 6012
rect 6436 6010 6460 6012
rect 6516 6010 6522 6012
rect 6276 5958 6278 6010
rect 6458 5958 6460 6010
rect 6214 5956 6220 5958
rect 6276 5956 6300 5958
rect 6356 5956 6380 5958
rect 6436 5956 6460 5958
rect 6516 5956 6522 5958
rect 6214 5947 6522 5956
rect 6564 5778 6592 6054
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 5814 2408 5870 2417
rect 5814 2343 5870 2352
rect 4894 2204 5202 2213
rect 4894 2202 4900 2204
rect 4956 2202 4980 2204
rect 5036 2202 5060 2204
rect 5116 2202 5140 2204
rect 5196 2202 5202 2204
rect 4956 2150 4958 2202
rect 5138 2150 5140 2202
rect 4894 2148 4900 2150
rect 4956 2148 4980 2150
rect 5036 2148 5060 2150
rect 5116 2148 5140 2150
rect 5196 2148 5202 2150
rect 4894 2139 5202 2148
rect 3882 1456 3938 1465
rect 3882 1391 3938 1400
rect 6104 762 6132 5510
rect 6564 5234 6592 5714
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6214 4924 6522 4933
rect 6214 4922 6220 4924
rect 6276 4922 6300 4924
rect 6356 4922 6380 4924
rect 6436 4922 6460 4924
rect 6516 4922 6522 4924
rect 6276 4870 6278 4922
rect 6458 4870 6460 4922
rect 6214 4868 6220 4870
rect 6276 4868 6300 4870
rect 6356 4868 6380 4870
rect 6436 4868 6460 4870
rect 6516 4868 6522 4870
rect 6214 4859 6522 4868
rect 6748 4690 6776 6190
rect 6932 5710 6960 6190
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7208 5642 7236 6326
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 6894 5468 7202 5477
rect 6894 5466 6900 5468
rect 6956 5466 6980 5468
rect 7036 5466 7060 5468
rect 7116 5466 7140 5468
rect 7196 5466 7202 5468
rect 6956 5414 6958 5466
rect 7138 5414 7140 5466
rect 6894 5412 6900 5414
rect 6956 5412 6980 5414
rect 7036 5412 7060 5414
rect 7116 5412 7140 5414
rect 7196 5412 7202 5414
rect 6894 5403 7202 5412
rect 7300 5302 7328 7482
rect 7392 6390 7420 8366
rect 7668 7818 7696 8502
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7852 7750 7880 8978
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7018 7880 7686
rect 8036 7410 8064 8842
rect 8128 8634 8156 14311
rect 8214 12540 8522 12549
rect 8214 12538 8220 12540
rect 8276 12538 8300 12540
rect 8356 12538 8380 12540
rect 8436 12538 8460 12540
rect 8516 12538 8522 12540
rect 8276 12486 8278 12538
rect 8458 12486 8460 12538
rect 8214 12484 8220 12486
rect 8276 12484 8300 12486
rect 8356 12484 8380 12486
rect 8436 12484 8460 12486
rect 8516 12484 8522 12486
rect 8214 12475 8522 12484
rect 8894 11996 9202 12005
rect 8894 11994 8900 11996
rect 8956 11994 8980 11996
rect 9036 11994 9060 11996
rect 9116 11994 9140 11996
rect 9196 11994 9202 11996
rect 8956 11942 8958 11994
rect 9138 11942 9140 11994
rect 8894 11940 8900 11942
rect 8956 11940 8980 11942
rect 9036 11940 9060 11942
rect 9116 11940 9140 11942
rect 9196 11940 9202 11942
rect 8894 11931 9202 11940
rect 8214 11452 8522 11461
rect 8214 11450 8220 11452
rect 8276 11450 8300 11452
rect 8356 11450 8380 11452
rect 8436 11450 8460 11452
rect 8516 11450 8522 11452
rect 8276 11398 8278 11450
rect 8458 11398 8460 11450
rect 8214 11396 8220 11398
rect 8276 11396 8300 11398
rect 8356 11396 8380 11398
rect 8436 11396 8460 11398
rect 8516 11396 8522 11398
rect 8214 11387 8522 11396
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 10742 8248 11154
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 10742 8616 10950
rect 8894 10908 9202 10917
rect 8894 10906 8900 10908
rect 8956 10906 8980 10908
rect 9036 10906 9060 10908
rect 9116 10906 9140 10908
rect 9196 10906 9202 10908
rect 8956 10854 8958 10906
rect 9138 10854 9140 10906
rect 8894 10852 8900 10854
rect 8956 10852 8980 10854
rect 9036 10852 9060 10854
rect 9116 10852 9140 10854
rect 9196 10852 9202 10854
rect 8894 10843 9202 10852
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8214 10364 8522 10373
rect 8214 10362 8220 10364
rect 8276 10362 8300 10364
rect 8356 10362 8380 10364
rect 8436 10362 8460 10364
rect 8516 10362 8522 10364
rect 8276 10310 8278 10362
rect 8458 10310 8460 10362
rect 8214 10308 8220 10310
rect 8276 10308 8300 10310
rect 8356 10308 8380 10310
rect 8436 10308 8460 10310
rect 8516 10308 8522 10310
rect 8214 10299 8522 10308
rect 8894 9820 9202 9829
rect 8894 9818 8900 9820
rect 8956 9818 8980 9820
rect 9036 9818 9060 9820
rect 9116 9818 9140 9820
rect 9196 9818 9202 9820
rect 8956 9766 8958 9818
rect 9138 9766 9140 9818
rect 8894 9764 8900 9766
rect 8956 9764 8980 9766
rect 9036 9764 9060 9766
rect 9116 9764 9140 9766
rect 9196 9764 9202 9766
rect 8894 9755 9202 9764
rect 8206 9616 8262 9625
rect 8206 9551 8208 9560
rect 8260 9551 8262 9560
rect 8208 9522 8260 9528
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8214 9276 8522 9285
rect 8214 9274 8220 9276
rect 8276 9274 8300 9276
rect 8356 9274 8380 9276
rect 8436 9274 8460 9276
rect 8516 9274 8522 9276
rect 8276 9222 8278 9274
rect 8458 9222 8460 9274
rect 8214 9220 8220 9222
rect 8276 9220 8300 9222
rect 8356 9220 8380 9222
rect 8436 9220 8460 9222
rect 8516 9220 8522 9222
rect 8214 9211 8522 9220
rect 8680 9042 8708 9454
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8680 8294 8708 8978
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8214 8188 8522 8197
rect 8214 8186 8220 8188
rect 8276 8186 8300 8188
rect 8356 8186 8380 8188
rect 8436 8186 8460 8188
rect 8516 8186 8522 8188
rect 8276 8134 8278 8186
rect 8458 8134 8460 8186
rect 8214 8132 8220 8134
rect 8276 8132 8300 8134
rect 8356 8132 8380 8134
rect 8436 8132 8460 8134
rect 8516 8132 8522 8134
rect 8214 8123 8522 8132
rect 8680 7886 8708 8230
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8680 7342 8708 7822
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8214 7100 8522 7109
rect 8214 7098 8220 7100
rect 8276 7098 8300 7100
rect 8356 7098 8380 7100
rect 8436 7098 8460 7100
rect 8516 7098 8522 7100
rect 8276 7046 8278 7098
rect 8458 7046 8460 7098
rect 8214 7044 8220 7046
rect 8276 7044 8300 7046
rect 8356 7044 8380 7046
rect 8436 7044 8460 7046
rect 8516 7044 8522 7046
rect 8214 7035 8522 7044
rect 7760 7002 7880 7018
rect 7748 6996 7880 7002
rect 7800 6990 7880 6996
rect 7748 6938 7800 6944
rect 8588 6866 8616 7278
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 8036 6254 8064 6734
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8588 6390 8616 6666
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6214 3836 6522 3845
rect 6214 3834 6220 3836
rect 6276 3834 6300 3836
rect 6356 3834 6380 3836
rect 6436 3834 6460 3836
rect 6516 3834 6522 3836
rect 6276 3782 6278 3834
rect 6458 3782 6460 3834
rect 6214 3780 6220 3782
rect 6276 3780 6300 3782
rect 6356 3780 6380 3782
rect 6436 3780 6460 3782
rect 6516 3780 6522 3782
rect 6214 3771 6522 3780
rect 6748 3738 6776 4626
rect 6894 4380 7202 4389
rect 6894 4378 6900 4380
rect 6956 4378 6980 4380
rect 7036 4378 7060 4380
rect 7116 4378 7140 4380
rect 7196 4378 7202 4380
rect 6956 4326 6958 4378
rect 7138 4326 7140 4378
rect 6894 4324 6900 4326
rect 6956 4324 6980 4326
rect 7036 4324 7060 4326
rect 7116 4324 7140 4326
rect 7196 4324 7202 4326
rect 6894 4315 7202 4324
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6840 3738 6868 3946
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6748 3194 6776 3674
rect 7392 3482 7420 6190
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8214 6012 8522 6021
rect 8214 6010 8220 6012
rect 8276 6010 8300 6012
rect 8356 6010 8380 6012
rect 8436 6010 8460 6012
rect 8516 6010 8522 6012
rect 8276 5958 8278 6010
rect 8458 5958 8460 6010
rect 8214 5956 8220 5958
rect 8276 5956 8300 5958
rect 8356 5956 8380 5958
rect 8436 5956 8460 5958
rect 8516 5956 8522 5958
rect 8214 5947 8522 5956
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7484 4826 7512 5578
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5137 8524 5510
rect 8588 5273 8616 6054
rect 8574 5264 8630 5273
rect 8574 5199 8630 5208
rect 8482 5128 8538 5137
rect 8482 5063 8538 5072
rect 8214 4924 8522 4933
rect 8214 4922 8220 4924
rect 8276 4922 8300 4924
rect 8356 4922 8380 4924
rect 8436 4922 8460 4924
rect 8516 4922 8522 4924
rect 8276 4870 8278 4922
rect 8458 4870 8460 4922
rect 8214 4868 8220 4870
rect 8276 4868 8300 4870
rect 8356 4868 8380 4870
rect 8436 4868 8460 4870
rect 8516 4868 8522 4870
rect 8214 4859 8522 4868
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7484 4214 7512 4762
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8312 4282 8340 4490
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 7472 4208 7524 4214
rect 8496 4185 8524 4422
rect 7472 4150 7524 4156
rect 8482 4176 8538 4185
rect 8482 4111 8538 4120
rect 8214 3836 8522 3845
rect 8214 3834 8220 3836
rect 8276 3834 8300 3836
rect 8356 3834 8380 3836
rect 8436 3834 8460 3836
rect 8516 3834 8522 3836
rect 8276 3782 8278 3834
rect 8458 3782 8460 3834
rect 8214 3780 8220 3782
rect 8276 3780 8300 3782
rect 8356 3780 8380 3782
rect 8436 3780 8460 3782
rect 8516 3780 8522 3782
rect 8214 3771 8522 3780
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 7300 3466 7420 3482
rect 7288 3460 7420 3466
rect 7340 3454 7420 3460
rect 7288 3402 7340 3408
rect 6894 3292 7202 3301
rect 6894 3290 6900 3292
rect 6956 3290 6980 3292
rect 7036 3290 7060 3292
rect 7116 3290 7140 3292
rect 7196 3290 7202 3292
rect 6956 3238 6958 3290
rect 7138 3238 7140 3290
rect 6894 3236 6900 3238
rect 6956 3236 6980 3238
rect 7036 3236 7060 3238
rect 7116 3236 7140 3238
rect 7196 3236 7202 3238
rect 6894 3227 7202 3236
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6214 2748 6522 2757
rect 6214 2746 6220 2748
rect 6276 2746 6300 2748
rect 6356 2746 6380 2748
rect 6436 2746 6460 2748
rect 6516 2746 6522 2748
rect 6276 2694 6278 2746
rect 6458 2694 6460 2746
rect 6214 2692 6220 2694
rect 6276 2692 6300 2694
rect 6356 2692 6380 2694
rect 6436 2692 6460 2694
rect 6516 2692 6522 2694
rect 6214 2683 6522 2692
rect 6748 1465 6776 3130
rect 7392 2774 7420 3454
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7852 3126 7880 3334
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 8588 3058 8616 3538
rect 8680 3398 8708 6394
rect 8772 3942 8800 8910
rect 8894 8732 9202 8741
rect 8894 8730 8900 8732
rect 8956 8730 8980 8732
rect 9036 8730 9060 8732
rect 9116 8730 9140 8732
rect 9196 8730 9202 8732
rect 8956 8678 8958 8730
rect 9138 8678 9140 8730
rect 8894 8676 8900 8678
rect 8956 8676 8980 8678
rect 9036 8676 9060 8678
rect 9116 8676 9140 8678
rect 9196 8676 9202 8678
rect 8894 8667 9202 8676
rect 9232 8090 9260 14991
rect 10782 13696 10838 13705
rect 10782 13631 10838 13640
rect 10598 13016 10654 13025
rect 10598 12951 10654 12960
rect 10214 12540 10522 12549
rect 10214 12538 10220 12540
rect 10276 12538 10300 12540
rect 10356 12538 10380 12540
rect 10436 12538 10460 12540
rect 10516 12538 10522 12540
rect 10276 12486 10278 12538
rect 10458 12486 10460 12538
rect 10214 12484 10220 12486
rect 10276 12484 10300 12486
rect 10356 12484 10380 12486
rect 10436 12484 10460 12486
rect 10516 12484 10522 12486
rect 10214 12475 10522 12484
rect 10214 11452 10522 11461
rect 10214 11450 10220 11452
rect 10276 11450 10300 11452
rect 10356 11450 10380 11452
rect 10436 11450 10460 11452
rect 10516 11450 10522 11452
rect 10276 11398 10278 11450
rect 10458 11398 10460 11450
rect 10214 11396 10220 11398
rect 10276 11396 10300 11398
rect 10356 11396 10380 11398
rect 10436 11396 10460 11398
rect 10516 11396 10522 11398
rect 10214 11387 10522 11396
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10810 9720 11018
rect 9784 10810 9812 11154
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9310 10160 9366 10169
rect 9310 10095 9366 10104
rect 9324 8498 9352 10095
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 9518 9444 9998
rect 10152 9994 10180 10678
rect 10214 10364 10522 10373
rect 10214 10362 10220 10364
rect 10276 10362 10300 10364
rect 10356 10362 10380 10364
rect 10436 10362 10460 10364
rect 10516 10362 10522 10364
rect 10276 10310 10278 10362
rect 10458 10310 10460 10362
rect 10214 10308 10220 10310
rect 10276 10308 10300 10310
rect 10356 10308 10380 10310
rect 10436 10308 10460 10310
rect 10516 10308 10522 10310
rect 10214 10299 10522 10308
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 8894 7644 9202 7653
rect 8894 7642 8900 7644
rect 8956 7642 8980 7644
rect 9036 7642 9060 7644
rect 9116 7642 9140 7644
rect 9196 7642 9202 7644
rect 8956 7590 8958 7642
rect 9138 7590 9140 7642
rect 8894 7588 8900 7590
rect 8956 7588 8980 7590
rect 9036 7588 9060 7590
rect 9116 7588 9140 7590
rect 9196 7588 9202 7590
rect 8894 7579 9202 7588
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8864 6866 8892 7346
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8956 7002 8984 7142
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8956 6905 8984 6938
rect 8942 6896 8998 6905
rect 8852 6860 8904 6866
rect 8942 6831 8998 6840
rect 8852 6802 8904 6808
rect 8894 6556 9202 6565
rect 8894 6554 8900 6556
rect 8956 6554 8980 6556
rect 9036 6554 9060 6556
rect 9116 6554 9140 6556
rect 9196 6554 9202 6556
rect 8956 6502 8958 6554
rect 9138 6502 9140 6554
rect 8894 6500 8900 6502
rect 8956 6500 8980 6502
rect 9036 6500 9060 6502
rect 9116 6500 9140 6502
rect 9196 6500 9202 6502
rect 8894 6491 9202 6500
rect 8894 5468 9202 5477
rect 8894 5466 8900 5468
rect 8956 5466 8980 5468
rect 9036 5466 9060 5468
rect 9116 5466 9140 5468
rect 9196 5466 9202 5468
rect 8956 5414 8958 5466
rect 9138 5414 9140 5466
rect 8894 5412 8900 5414
rect 8956 5412 8980 5414
rect 9036 5412 9060 5414
rect 9116 5412 9140 5414
rect 9196 5412 9202 5414
rect 8894 5403 9202 5412
rect 8894 4380 9202 4389
rect 8894 4378 8900 4380
rect 8956 4378 8980 4380
rect 9036 4378 9060 4380
rect 9116 4378 9140 4380
rect 9196 4378 9202 4380
rect 8956 4326 8958 4378
rect 9138 4326 9140 4378
rect 8894 4324 8900 4326
rect 8956 4324 8980 4326
rect 9036 4324 9060 4326
rect 9116 4324 9140 4326
rect 9196 4324 9202 4326
rect 8894 4315 9202 4324
rect 9324 3942 9352 7278
rect 9416 4486 9444 8774
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9508 6798 9536 7754
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9508 6254 9536 6734
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9508 5710 9536 6190
rect 9784 6118 9812 9454
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9508 5030 9536 5646
rect 9876 5574 9904 9862
rect 10152 9654 10180 9930
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10152 8888 10180 9590
rect 10214 9276 10522 9285
rect 10214 9274 10220 9276
rect 10276 9274 10300 9276
rect 10356 9274 10380 9276
rect 10436 9274 10460 9276
rect 10516 9274 10522 9276
rect 10276 9222 10278 9274
rect 10458 9222 10460 9274
rect 10214 9220 10220 9222
rect 10276 9220 10300 9222
rect 10356 9220 10380 9222
rect 10436 9220 10460 9222
rect 10516 9220 10522 9222
rect 10214 9211 10522 9220
rect 10232 8900 10284 8906
rect 10152 8860 10232 8888
rect 10152 7800 10180 8860
rect 10232 8842 10284 8848
rect 10214 8188 10522 8197
rect 10214 8186 10220 8188
rect 10276 8186 10300 8188
rect 10356 8186 10380 8188
rect 10436 8186 10460 8188
rect 10516 8186 10522 8188
rect 10276 8134 10278 8186
rect 10458 8134 10460 8186
rect 10214 8132 10220 8134
rect 10276 8132 10300 8134
rect 10356 8132 10380 8134
rect 10436 8132 10460 8134
rect 10516 8132 10522 8134
rect 10214 8123 10522 8132
rect 10232 7812 10284 7818
rect 10060 7772 10232 7800
rect 10060 7478 10088 7772
rect 10232 7754 10284 7760
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10060 7002 10088 7414
rect 10612 7342 10640 12951
rect 10796 12434 10824 13631
rect 10704 12406 10824 12434
rect 10704 8090 10732 12406
rect 10782 12336 10838 12345
rect 10782 12271 10838 12280
rect 10796 9178 10824 12271
rect 10894 11996 11202 12005
rect 10894 11994 10900 11996
rect 10956 11994 10980 11996
rect 11036 11994 11060 11996
rect 11116 11994 11140 11996
rect 11196 11994 11202 11996
rect 10956 11942 10958 11994
rect 11138 11942 11140 11994
rect 10894 11940 10900 11942
rect 10956 11940 10980 11942
rect 11036 11940 11060 11942
rect 11116 11940 11140 11942
rect 11196 11940 11202 11942
rect 10894 11931 11202 11940
rect 11242 11656 11298 11665
rect 11242 11591 11298 11600
rect 10894 10908 11202 10917
rect 10894 10906 10900 10908
rect 10956 10906 10980 10908
rect 11036 10906 11060 10908
rect 11116 10906 11140 10908
rect 11196 10906 11202 10908
rect 10956 10854 10958 10906
rect 11138 10854 11140 10906
rect 10894 10852 10900 10854
rect 10956 10852 10980 10854
rect 11036 10852 11060 10854
rect 11116 10852 11140 10854
rect 11196 10852 11202 10854
rect 10894 10843 11202 10852
rect 11256 10266 11284 11591
rect 11334 10976 11390 10985
rect 11334 10911 11390 10920
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 10894 9820 11202 9829
rect 10894 9818 10900 9820
rect 10956 9818 10980 9820
rect 11036 9818 11060 9820
rect 11116 9818 11140 9820
rect 11196 9818 11202 9820
rect 10956 9766 10958 9818
rect 11138 9766 11140 9818
rect 10894 9764 10900 9766
rect 10956 9764 10980 9766
rect 11036 9764 11060 9766
rect 11116 9764 11140 9766
rect 11196 9764 11202 9766
rect 10894 9755 11202 9764
rect 11348 9518 11376 10911
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10966 8936 11022 8945
rect 10796 8265 10824 8910
rect 10966 8871 11022 8880
rect 10980 8838 11008 8871
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10894 8732 11202 8741
rect 10894 8730 10900 8732
rect 10956 8730 10980 8732
rect 11036 8730 11060 8732
rect 11116 8730 11140 8732
rect 11196 8730 11202 8732
rect 10956 8678 10958 8730
rect 11138 8678 11140 8730
rect 10894 8676 10900 8678
rect 10956 8676 10980 8678
rect 11036 8676 11060 8678
rect 11116 8676 11140 8678
rect 11196 8676 11202 8678
rect 10894 8667 11202 8676
rect 10782 8256 10838 8265
rect 10782 8191 10838 8200
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10214 7100 10522 7109
rect 10214 7098 10220 7100
rect 10276 7098 10300 7100
rect 10356 7098 10380 7100
rect 10436 7098 10460 7100
rect 10516 7098 10522 7100
rect 10276 7046 10278 7098
rect 10458 7046 10460 7098
rect 10214 7044 10220 7046
rect 10276 7044 10300 7046
rect 10356 7044 10380 7046
rect 10436 7044 10460 7046
rect 10516 7044 10522 7046
rect 10214 7035 10522 7044
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10796 6882 10824 8191
rect 10894 7644 11202 7653
rect 10894 7642 10900 7644
rect 10956 7642 10980 7644
rect 11036 7642 11060 7644
rect 11116 7642 11140 7644
rect 11196 7642 11202 7644
rect 10956 7590 10958 7642
rect 11138 7590 11140 7642
rect 10894 7588 10900 7590
rect 10956 7588 10980 7590
rect 11036 7588 11060 7590
rect 11116 7588 11140 7590
rect 11196 7588 11202 7590
rect 10894 7579 11202 7588
rect 11334 7576 11390 7585
rect 11334 7511 11336 7520
rect 11388 7511 11390 7520
rect 11336 7482 11388 7488
rect 10704 6866 10824 6882
rect 10692 6860 10824 6866
rect 10744 6854 10824 6860
rect 10692 6802 10744 6808
rect 10704 6730 10732 6802
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10796 6390 10824 6854
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 10894 6556 11202 6565
rect 10894 6554 10900 6556
rect 10956 6554 10980 6556
rect 11036 6554 11060 6556
rect 11116 6554 11140 6556
rect 11196 6554 11202 6556
rect 10956 6502 10958 6554
rect 11138 6502 11140 6554
rect 10894 6500 10900 6502
rect 10956 6500 10980 6502
rect 11036 6500 11060 6502
rect 11116 6500 11140 6502
rect 11196 6500 11202 6502
rect 10894 6491 11202 6500
rect 10784 6384 10836 6390
rect 10836 6344 10916 6372
rect 10784 6326 10836 6332
rect 10214 6012 10522 6021
rect 10214 6010 10220 6012
rect 10276 6010 10300 6012
rect 10356 6010 10380 6012
rect 10436 6010 10460 6012
rect 10516 6010 10522 6012
rect 10276 5958 10278 6010
rect 10458 5958 10460 6010
rect 10214 5956 10220 5958
rect 10276 5956 10300 5958
rect 10356 5956 10380 5958
rect 10436 5956 10460 5958
rect 10516 5956 10522 5958
rect 10214 5947 10522 5956
rect 10888 5710 10916 6344
rect 11440 6254 11468 6598
rect 11428 6248 11480 6254
rect 11426 6216 11428 6225
rect 11480 6216 11482 6225
rect 11426 6151 11482 6160
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5778 11468 6054
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 10876 5704 10928 5710
rect 10704 5652 10876 5658
rect 10704 5646 10928 5652
rect 10704 5630 10916 5646
rect 10704 5574 10732 5630
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 11336 5568 11388 5574
rect 11440 5545 11468 5714
rect 11336 5510 11388 5516
rect 11426 5536 11482 5545
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9692 5166 9720 5306
rect 10704 5302 10732 5510
rect 10894 5468 11202 5477
rect 10894 5466 10900 5468
rect 10956 5466 10980 5468
rect 11036 5466 11060 5468
rect 11116 5466 11140 5468
rect 11196 5466 11202 5468
rect 10956 5414 10958 5466
rect 11138 5414 11140 5466
rect 10894 5412 10900 5414
rect 10956 5412 10980 5414
rect 11036 5412 11060 5414
rect 11116 5412 11140 5414
rect 11196 5412 11202 5414
rect 10894 5403 11202 5412
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9508 4078 9536 4966
rect 10214 4924 10522 4933
rect 10214 4922 10220 4924
rect 10276 4922 10300 4924
rect 10356 4922 10380 4924
rect 10436 4922 10460 4924
rect 10516 4922 10522 4924
rect 10276 4870 10278 4922
rect 10458 4870 10460 4922
rect 10214 4868 10220 4870
rect 10276 4868 10300 4870
rect 10356 4868 10380 4870
rect 10436 4868 10460 4870
rect 10516 4868 10522 4870
rect 10214 4859 10522 4868
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9784 4078 9812 4626
rect 10704 4282 10732 5238
rect 11348 5166 11376 5510
rect 11426 5471 11482 5480
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 10894 4380 11202 4389
rect 10894 4378 10900 4380
rect 10956 4378 10980 4380
rect 11036 4378 11060 4380
rect 11116 4378 11140 4380
rect 11196 4378 11202 4380
rect 10956 4326 10958 4378
rect 11138 4326 11140 4378
rect 10894 4324 10900 4326
rect 10956 4324 10980 4326
rect 11036 4324 11060 4326
rect 11116 4324 11140 4326
rect 11196 4324 11202 4326
rect 10894 4315 11202 4324
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10704 4162 10732 4218
rect 11256 4214 11284 4966
rect 11348 4865 11376 5102
rect 11334 4856 11390 4865
rect 11334 4791 11390 4800
rect 11244 4208 11296 4214
rect 11242 4176 11244 4185
rect 11296 4176 11298 4185
rect 10704 4146 10824 4162
rect 10704 4140 10836 4146
rect 10704 4134 10784 4140
rect 11242 4111 11298 4120
rect 10784 4082 10836 4088
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8772 3126 8800 3878
rect 8956 3505 8984 3878
rect 9508 3602 9536 4014
rect 10214 3836 10522 3845
rect 10214 3834 10220 3836
rect 10276 3834 10300 3836
rect 10356 3834 10380 3836
rect 10436 3834 10460 3836
rect 10516 3834 10522 3836
rect 10276 3782 10278 3834
rect 10458 3782 10460 3834
rect 10214 3780 10220 3782
rect 10276 3780 10300 3782
rect 10356 3780 10380 3782
rect 10436 3780 10460 3782
rect 10516 3780 10522 3782
rect 10214 3771 10522 3780
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 8942 3496 8998 3505
rect 8942 3431 8998 3440
rect 10796 3482 10824 4082
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11256 3602 11284 3878
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11256 3505 11284 3538
rect 11242 3496 11298 3505
rect 10796 3466 10916 3482
rect 10796 3460 10928 3466
rect 10796 3454 10876 3460
rect 10796 3398 10824 3454
rect 11242 3431 11298 3440
rect 10876 3402 10928 3408
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 8894 3292 9202 3301
rect 8894 3290 8900 3292
rect 8956 3290 8980 3292
rect 9036 3290 9060 3292
rect 9116 3290 9140 3292
rect 9196 3290 9202 3292
rect 8956 3238 8958 3290
rect 9138 3238 9140 3290
rect 8894 3236 8900 3238
rect 8956 3236 8980 3238
rect 9036 3236 9060 3238
rect 9116 3236 9140 3238
rect 9196 3236 9202 3238
rect 8894 3227 9202 3236
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 7300 2746 7420 2774
rect 8214 2748 8522 2757
rect 8214 2746 8220 2748
rect 8276 2746 8300 2748
rect 8356 2746 8380 2748
rect 8436 2746 8460 2748
rect 8516 2746 8522 2748
rect 6894 2204 7202 2213
rect 6894 2202 6900 2204
rect 6956 2202 6980 2204
rect 7036 2202 7060 2204
rect 7116 2202 7140 2204
rect 7196 2202 7202 2204
rect 6956 2150 6958 2202
rect 7138 2150 7140 2202
rect 6894 2148 6900 2150
rect 6956 2148 6980 2150
rect 7036 2148 7060 2150
rect 7116 2148 7140 2150
rect 7196 2148 7202 2150
rect 6894 2139 7202 2148
rect 6734 1456 6790 1465
rect 6734 1391 6790 1400
rect 6380 870 6500 898
rect 6380 762 6408 870
rect 6472 800 6500 870
rect 6104 734 6408 762
rect 2962 96 3018 105
rect 2962 31 3018 40
rect 6458 0 6514 800
rect 7300 785 7328 2746
rect 8276 2694 8278 2746
rect 8458 2694 8460 2746
rect 8214 2692 8220 2694
rect 8276 2692 8300 2694
rect 8356 2692 8380 2694
rect 8436 2692 8460 2694
rect 8516 2692 8522 2694
rect 8214 2683 8522 2692
rect 8894 2204 9202 2213
rect 8894 2202 8900 2204
rect 8956 2202 8980 2204
rect 9036 2202 9060 2204
rect 9116 2202 9140 2204
rect 9196 2202 9202 2204
rect 8956 2150 8958 2202
rect 9138 2150 9140 2202
rect 8894 2148 8900 2150
rect 8956 2148 8980 2150
rect 9036 2148 9060 2150
rect 9116 2148 9140 2150
rect 9196 2148 9202 2150
rect 8894 2139 9202 2148
rect 7286 776 7342 785
rect 7286 711 7342 720
rect 9232 105 9260 3334
rect 10796 3126 10824 3334
rect 10894 3292 11202 3301
rect 10894 3290 10900 3292
rect 10956 3290 10980 3292
rect 11036 3290 11060 3292
rect 11116 3290 11140 3292
rect 11196 3290 11202 3292
rect 10956 3238 10958 3290
rect 11138 3238 11140 3290
rect 10894 3236 10900 3238
rect 10956 3236 10980 3238
rect 11036 3236 11060 3238
rect 11116 3236 11140 3238
rect 11196 3236 11202 3238
rect 10894 3227 11202 3236
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 11348 2990 11376 3334
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11348 2825 11376 2926
rect 11334 2816 11390 2825
rect 10214 2748 10522 2757
rect 11334 2751 11390 2760
rect 10214 2746 10220 2748
rect 10276 2746 10300 2748
rect 10356 2746 10380 2748
rect 10436 2746 10460 2748
rect 10516 2746 10522 2748
rect 10276 2694 10278 2746
rect 10458 2694 10460 2746
rect 10214 2692 10220 2694
rect 10276 2692 10300 2694
rect 10356 2692 10380 2694
rect 10436 2692 10460 2694
rect 10516 2692 10522 2694
rect 10214 2683 10522 2692
rect 10894 2204 11202 2213
rect 10894 2202 10900 2204
rect 10956 2202 10980 2204
rect 11036 2202 11060 2204
rect 11116 2202 11140 2204
rect 11196 2202 11202 2204
rect 10956 2150 10958 2202
rect 11138 2150 11140 2202
rect 10894 2148 10900 2150
rect 10956 2148 10980 2150
rect 11036 2148 11060 2150
rect 11116 2148 11140 2150
rect 11196 2148 11202 2150
rect 10894 2139 11202 2148
rect 11440 2145 11468 3130
rect 11426 2136 11482 2145
rect 11426 2071 11482 2080
rect 9218 96 9274 105
rect 9218 31 9274 40
<< via2 >>
rect 2962 15000 3018 15056
rect 9218 15000 9274 15056
rect 2870 14320 2926 14376
rect 2778 12960 2834 13016
rect 1306 8880 1362 8936
rect 8114 14320 8170 14376
rect 3146 13640 3202 13696
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 6220 12538 6276 12540
rect 6300 12538 6356 12540
rect 6380 12538 6436 12540
rect 6460 12538 6516 12540
rect 6220 12486 6266 12538
rect 6266 12486 6276 12538
rect 6300 12486 6330 12538
rect 6330 12486 6342 12538
rect 6342 12486 6356 12538
rect 6380 12486 6394 12538
rect 6394 12486 6406 12538
rect 6406 12486 6436 12538
rect 6460 12486 6470 12538
rect 6470 12486 6516 12538
rect 6220 12484 6276 12486
rect 6300 12484 6356 12486
rect 6380 12484 6436 12486
rect 6460 12484 6516 12486
rect 2778 7520 2834 7576
rect 1214 6840 1270 6896
rect 3882 12280 3938 12336
rect 4900 11994 4956 11996
rect 4980 11994 5036 11996
rect 5060 11994 5116 11996
rect 5140 11994 5196 11996
rect 4900 11942 4946 11994
rect 4946 11942 4956 11994
rect 4980 11942 5010 11994
rect 5010 11942 5022 11994
rect 5022 11942 5036 11994
rect 5060 11942 5074 11994
rect 5074 11942 5086 11994
rect 5086 11942 5116 11994
rect 5140 11942 5150 11994
rect 5150 11942 5196 11994
rect 4900 11940 4956 11942
rect 4980 11940 5036 11942
rect 5060 11940 5116 11942
rect 5140 11940 5196 11942
rect 6900 11994 6956 11996
rect 6980 11994 7036 11996
rect 7060 11994 7116 11996
rect 7140 11994 7196 11996
rect 6900 11942 6946 11994
rect 6946 11942 6956 11994
rect 6980 11942 7010 11994
rect 7010 11942 7022 11994
rect 7022 11942 7036 11994
rect 7060 11942 7074 11994
rect 7074 11942 7086 11994
rect 7086 11942 7116 11994
rect 7140 11942 7150 11994
rect 7150 11942 7196 11994
rect 6900 11940 6956 11942
rect 6980 11940 7036 11942
rect 7060 11940 7116 11942
rect 7140 11940 7196 11942
rect 6090 11600 6146 11656
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4618 10920 4674 10976
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4066 9560 4122 9616
rect 3882 8200 3938 8256
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3606 6160 3662 6216
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4900 10906 4956 10908
rect 4980 10906 5036 10908
rect 5060 10906 5116 10908
rect 5140 10906 5196 10908
rect 4900 10854 4946 10906
rect 4946 10854 4956 10906
rect 4980 10854 5010 10906
rect 5010 10854 5022 10906
rect 5022 10854 5036 10906
rect 5060 10854 5074 10906
rect 5074 10854 5086 10906
rect 5086 10854 5116 10906
rect 5140 10854 5150 10906
rect 5150 10854 5196 10906
rect 4900 10852 4956 10854
rect 4980 10852 5036 10854
rect 5060 10852 5116 10854
rect 5140 10852 5196 10854
rect 4900 9818 4956 9820
rect 4980 9818 5036 9820
rect 5060 9818 5116 9820
rect 5140 9818 5196 9820
rect 4900 9766 4946 9818
rect 4946 9766 4956 9818
rect 4980 9766 5010 9818
rect 5010 9766 5022 9818
rect 5022 9766 5036 9818
rect 5060 9766 5074 9818
rect 5074 9766 5086 9818
rect 5086 9766 5116 9818
rect 5140 9766 5150 9818
rect 5150 9766 5196 9818
rect 4900 9764 4956 9766
rect 4980 9764 5036 9766
rect 5060 9764 5116 9766
rect 5140 9764 5196 9766
rect 4900 8730 4956 8732
rect 4980 8730 5036 8732
rect 5060 8730 5116 8732
rect 5140 8730 5196 8732
rect 4900 8678 4946 8730
rect 4946 8678 4956 8730
rect 4980 8678 5010 8730
rect 5010 8678 5022 8730
rect 5022 8678 5036 8730
rect 5060 8678 5074 8730
rect 5074 8678 5086 8730
rect 5086 8678 5116 8730
rect 5140 8678 5150 8730
rect 5150 8678 5196 8730
rect 4900 8676 4956 8678
rect 4980 8676 5036 8678
rect 5060 8676 5116 8678
rect 5140 8676 5196 8678
rect 4900 7642 4956 7644
rect 4980 7642 5036 7644
rect 5060 7642 5116 7644
rect 5140 7642 5196 7644
rect 4900 7590 4946 7642
rect 4946 7590 4956 7642
rect 4980 7590 5010 7642
rect 5010 7590 5022 7642
rect 5022 7590 5036 7642
rect 5060 7590 5074 7642
rect 5074 7590 5086 7642
rect 5086 7590 5116 7642
rect 5140 7590 5150 7642
rect 5150 7590 5196 7642
rect 4900 7588 4956 7590
rect 4980 7588 5036 7590
rect 5060 7588 5116 7590
rect 5140 7588 5196 7590
rect 4900 6554 4956 6556
rect 4980 6554 5036 6556
rect 5060 6554 5116 6556
rect 5140 6554 5196 6556
rect 4900 6502 4946 6554
rect 4946 6502 4956 6554
rect 4980 6502 5010 6554
rect 5010 6502 5022 6554
rect 5022 6502 5036 6554
rect 5060 6502 5074 6554
rect 5074 6502 5086 6554
rect 5086 6502 5116 6554
rect 5140 6502 5150 6554
rect 5150 6502 5196 6554
rect 4900 6500 4956 6502
rect 4980 6500 5036 6502
rect 5060 6500 5116 6502
rect 5140 6500 5196 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4900 5466 4956 5468
rect 4980 5466 5036 5468
rect 5060 5466 5116 5468
rect 5140 5466 5196 5468
rect 4900 5414 4946 5466
rect 4946 5414 4956 5466
rect 4980 5414 5010 5466
rect 5010 5414 5022 5466
rect 5022 5414 5036 5466
rect 5060 5414 5074 5466
rect 5074 5414 5086 5466
rect 5086 5414 5116 5466
rect 5140 5414 5150 5466
rect 5150 5414 5196 5466
rect 4900 5412 4956 5414
rect 4980 5412 5036 5414
rect 5060 5412 5116 5414
rect 5140 5412 5196 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 2778 720 2834 776
rect 4900 4378 4956 4380
rect 4980 4378 5036 4380
rect 5060 4378 5116 4380
rect 5140 4378 5196 4380
rect 4900 4326 4946 4378
rect 4946 4326 4956 4378
rect 4980 4326 5010 4378
rect 5010 4326 5022 4378
rect 5022 4326 5036 4378
rect 5060 4326 5074 4378
rect 5074 4326 5086 4378
rect 5086 4326 5116 4378
rect 5140 4326 5150 4378
rect 5150 4326 5196 4378
rect 4900 4324 4956 4326
rect 4980 4324 5036 4326
rect 5060 4324 5116 4326
rect 5140 4324 5196 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4900 3290 4956 3292
rect 4980 3290 5036 3292
rect 5060 3290 5116 3292
rect 5140 3290 5196 3292
rect 4900 3238 4946 3290
rect 4946 3238 4956 3290
rect 4980 3238 5010 3290
rect 5010 3238 5022 3290
rect 5022 3238 5036 3290
rect 5060 3238 5074 3290
rect 5074 3238 5086 3290
rect 5086 3238 5116 3290
rect 5140 3238 5150 3290
rect 5150 3238 5196 3290
rect 4900 3236 4956 3238
rect 4980 3236 5036 3238
rect 5060 3236 5116 3238
rect 5140 3236 5196 3238
rect 4434 2896 4490 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6220 11450 6276 11452
rect 6300 11450 6356 11452
rect 6380 11450 6436 11452
rect 6460 11450 6516 11452
rect 6220 11398 6266 11450
rect 6266 11398 6276 11450
rect 6300 11398 6330 11450
rect 6330 11398 6342 11450
rect 6342 11398 6356 11450
rect 6380 11398 6394 11450
rect 6394 11398 6406 11450
rect 6406 11398 6436 11450
rect 6460 11398 6470 11450
rect 6470 11398 6516 11450
rect 6220 11396 6276 11398
rect 6300 11396 6356 11398
rect 6380 11396 6436 11398
rect 6460 11396 6516 11398
rect 6900 10906 6956 10908
rect 6980 10906 7036 10908
rect 7060 10906 7116 10908
rect 7140 10906 7196 10908
rect 6900 10854 6946 10906
rect 6946 10854 6956 10906
rect 6980 10854 7010 10906
rect 7010 10854 7022 10906
rect 7022 10854 7036 10906
rect 7060 10854 7074 10906
rect 7074 10854 7086 10906
rect 7086 10854 7116 10906
rect 7140 10854 7150 10906
rect 7150 10854 7196 10906
rect 6900 10852 6956 10854
rect 6980 10852 7036 10854
rect 7060 10852 7116 10854
rect 7140 10852 7196 10854
rect 6220 10362 6276 10364
rect 6300 10362 6356 10364
rect 6380 10362 6436 10364
rect 6460 10362 6516 10364
rect 6220 10310 6266 10362
rect 6266 10310 6276 10362
rect 6300 10310 6330 10362
rect 6330 10310 6342 10362
rect 6342 10310 6356 10362
rect 6380 10310 6394 10362
rect 6394 10310 6406 10362
rect 6406 10310 6436 10362
rect 6460 10310 6470 10362
rect 6470 10310 6516 10362
rect 6220 10308 6276 10310
rect 6300 10308 6356 10310
rect 6380 10308 6436 10310
rect 6460 10308 6516 10310
rect 6734 10104 6790 10160
rect 6220 9274 6276 9276
rect 6300 9274 6356 9276
rect 6380 9274 6436 9276
rect 6460 9274 6516 9276
rect 6220 9222 6266 9274
rect 6266 9222 6276 9274
rect 6300 9222 6330 9274
rect 6330 9222 6342 9274
rect 6342 9222 6356 9274
rect 6380 9222 6394 9274
rect 6394 9222 6406 9274
rect 6406 9222 6436 9274
rect 6460 9222 6470 9274
rect 6470 9222 6516 9274
rect 6220 9220 6276 9222
rect 6300 9220 6356 9222
rect 6380 9220 6436 9222
rect 6460 9220 6516 9222
rect 6900 9818 6956 9820
rect 6980 9818 7036 9820
rect 7060 9818 7116 9820
rect 7140 9818 7196 9820
rect 6900 9766 6946 9818
rect 6946 9766 6956 9818
rect 6980 9766 7010 9818
rect 7010 9766 7022 9818
rect 7022 9766 7036 9818
rect 7060 9766 7074 9818
rect 7074 9766 7086 9818
rect 7086 9766 7116 9818
rect 7140 9766 7150 9818
rect 7150 9766 7196 9818
rect 6900 9764 6956 9766
rect 6980 9764 7036 9766
rect 7060 9764 7116 9766
rect 7140 9764 7196 9766
rect 6220 8186 6276 8188
rect 6300 8186 6356 8188
rect 6380 8186 6436 8188
rect 6460 8186 6516 8188
rect 6220 8134 6266 8186
rect 6266 8134 6276 8186
rect 6300 8134 6330 8186
rect 6330 8134 6342 8186
rect 6342 8134 6356 8186
rect 6380 8134 6394 8186
rect 6394 8134 6406 8186
rect 6406 8134 6436 8186
rect 6460 8134 6470 8186
rect 6470 8134 6516 8186
rect 6220 8132 6276 8134
rect 6300 8132 6356 8134
rect 6380 8132 6436 8134
rect 6460 8132 6516 8134
rect 6900 8730 6956 8732
rect 6980 8730 7036 8732
rect 7060 8730 7116 8732
rect 7140 8730 7196 8732
rect 6900 8678 6946 8730
rect 6946 8678 6956 8730
rect 6980 8678 7010 8730
rect 7010 8678 7022 8730
rect 7022 8678 7036 8730
rect 7060 8678 7074 8730
rect 7074 8678 7086 8730
rect 7086 8678 7116 8730
rect 7140 8678 7150 8730
rect 7150 8678 7196 8730
rect 6900 8676 6956 8678
rect 6980 8676 7036 8678
rect 7060 8676 7116 8678
rect 7140 8676 7196 8678
rect 6900 7642 6956 7644
rect 6980 7642 7036 7644
rect 7060 7642 7116 7644
rect 7140 7642 7196 7644
rect 6900 7590 6946 7642
rect 6946 7590 6956 7642
rect 6980 7590 7010 7642
rect 7010 7590 7022 7642
rect 7022 7590 7036 7642
rect 7060 7590 7074 7642
rect 7074 7590 7086 7642
rect 7086 7590 7116 7642
rect 7140 7590 7150 7642
rect 7150 7590 7196 7642
rect 6900 7588 6956 7590
rect 6980 7588 7036 7590
rect 7060 7588 7116 7590
rect 7140 7588 7196 7590
rect 6220 7098 6276 7100
rect 6300 7098 6356 7100
rect 6380 7098 6436 7100
rect 6460 7098 6516 7100
rect 6220 7046 6266 7098
rect 6266 7046 6276 7098
rect 6300 7046 6330 7098
rect 6330 7046 6342 7098
rect 6342 7046 6356 7098
rect 6380 7046 6394 7098
rect 6394 7046 6406 7098
rect 6406 7046 6436 7098
rect 6460 7046 6470 7098
rect 6470 7046 6516 7098
rect 6220 7044 6276 7046
rect 6300 7044 6356 7046
rect 6380 7044 6436 7046
rect 6460 7044 6516 7046
rect 6900 6554 6956 6556
rect 6980 6554 7036 6556
rect 7060 6554 7116 6556
rect 7140 6554 7196 6556
rect 6900 6502 6946 6554
rect 6946 6502 6956 6554
rect 6980 6502 7010 6554
rect 7010 6502 7022 6554
rect 7022 6502 7036 6554
rect 7060 6502 7074 6554
rect 7074 6502 7086 6554
rect 7086 6502 7116 6554
rect 7140 6502 7150 6554
rect 7150 6502 7196 6554
rect 6900 6500 6956 6502
rect 6980 6500 7036 6502
rect 7060 6500 7116 6502
rect 7140 6500 7196 6502
rect 6220 6010 6276 6012
rect 6300 6010 6356 6012
rect 6380 6010 6436 6012
rect 6460 6010 6516 6012
rect 6220 5958 6266 6010
rect 6266 5958 6276 6010
rect 6300 5958 6330 6010
rect 6330 5958 6342 6010
rect 6342 5958 6356 6010
rect 6380 5958 6394 6010
rect 6394 5958 6406 6010
rect 6406 5958 6436 6010
rect 6460 5958 6470 6010
rect 6470 5958 6516 6010
rect 6220 5956 6276 5958
rect 6300 5956 6356 5958
rect 6380 5956 6436 5958
rect 6460 5956 6516 5958
rect 5814 2352 5870 2408
rect 4900 2202 4956 2204
rect 4980 2202 5036 2204
rect 5060 2202 5116 2204
rect 5140 2202 5196 2204
rect 4900 2150 4946 2202
rect 4946 2150 4956 2202
rect 4980 2150 5010 2202
rect 5010 2150 5022 2202
rect 5022 2150 5036 2202
rect 5060 2150 5074 2202
rect 5074 2150 5086 2202
rect 5086 2150 5116 2202
rect 5140 2150 5150 2202
rect 5150 2150 5196 2202
rect 4900 2148 4956 2150
rect 4980 2148 5036 2150
rect 5060 2148 5116 2150
rect 5140 2148 5196 2150
rect 3882 1400 3938 1456
rect 6220 4922 6276 4924
rect 6300 4922 6356 4924
rect 6380 4922 6436 4924
rect 6460 4922 6516 4924
rect 6220 4870 6266 4922
rect 6266 4870 6276 4922
rect 6300 4870 6330 4922
rect 6330 4870 6342 4922
rect 6342 4870 6356 4922
rect 6380 4870 6394 4922
rect 6394 4870 6406 4922
rect 6406 4870 6436 4922
rect 6460 4870 6470 4922
rect 6470 4870 6516 4922
rect 6220 4868 6276 4870
rect 6300 4868 6356 4870
rect 6380 4868 6436 4870
rect 6460 4868 6516 4870
rect 6900 5466 6956 5468
rect 6980 5466 7036 5468
rect 7060 5466 7116 5468
rect 7140 5466 7196 5468
rect 6900 5414 6946 5466
rect 6946 5414 6956 5466
rect 6980 5414 7010 5466
rect 7010 5414 7022 5466
rect 7022 5414 7036 5466
rect 7060 5414 7074 5466
rect 7074 5414 7086 5466
rect 7086 5414 7116 5466
rect 7140 5414 7150 5466
rect 7150 5414 7196 5466
rect 6900 5412 6956 5414
rect 6980 5412 7036 5414
rect 7060 5412 7116 5414
rect 7140 5412 7196 5414
rect 8220 12538 8276 12540
rect 8300 12538 8356 12540
rect 8380 12538 8436 12540
rect 8460 12538 8516 12540
rect 8220 12486 8266 12538
rect 8266 12486 8276 12538
rect 8300 12486 8330 12538
rect 8330 12486 8342 12538
rect 8342 12486 8356 12538
rect 8380 12486 8394 12538
rect 8394 12486 8406 12538
rect 8406 12486 8436 12538
rect 8460 12486 8470 12538
rect 8470 12486 8516 12538
rect 8220 12484 8276 12486
rect 8300 12484 8356 12486
rect 8380 12484 8436 12486
rect 8460 12484 8516 12486
rect 8900 11994 8956 11996
rect 8980 11994 9036 11996
rect 9060 11994 9116 11996
rect 9140 11994 9196 11996
rect 8900 11942 8946 11994
rect 8946 11942 8956 11994
rect 8980 11942 9010 11994
rect 9010 11942 9022 11994
rect 9022 11942 9036 11994
rect 9060 11942 9074 11994
rect 9074 11942 9086 11994
rect 9086 11942 9116 11994
rect 9140 11942 9150 11994
rect 9150 11942 9196 11994
rect 8900 11940 8956 11942
rect 8980 11940 9036 11942
rect 9060 11940 9116 11942
rect 9140 11940 9196 11942
rect 8220 11450 8276 11452
rect 8300 11450 8356 11452
rect 8380 11450 8436 11452
rect 8460 11450 8516 11452
rect 8220 11398 8266 11450
rect 8266 11398 8276 11450
rect 8300 11398 8330 11450
rect 8330 11398 8342 11450
rect 8342 11398 8356 11450
rect 8380 11398 8394 11450
rect 8394 11398 8406 11450
rect 8406 11398 8436 11450
rect 8460 11398 8470 11450
rect 8470 11398 8516 11450
rect 8220 11396 8276 11398
rect 8300 11396 8356 11398
rect 8380 11396 8436 11398
rect 8460 11396 8516 11398
rect 8900 10906 8956 10908
rect 8980 10906 9036 10908
rect 9060 10906 9116 10908
rect 9140 10906 9196 10908
rect 8900 10854 8946 10906
rect 8946 10854 8956 10906
rect 8980 10854 9010 10906
rect 9010 10854 9022 10906
rect 9022 10854 9036 10906
rect 9060 10854 9074 10906
rect 9074 10854 9086 10906
rect 9086 10854 9116 10906
rect 9140 10854 9150 10906
rect 9150 10854 9196 10906
rect 8900 10852 8956 10854
rect 8980 10852 9036 10854
rect 9060 10852 9116 10854
rect 9140 10852 9196 10854
rect 8220 10362 8276 10364
rect 8300 10362 8356 10364
rect 8380 10362 8436 10364
rect 8460 10362 8516 10364
rect 8220 10310 8266 10362
rect 8266 10310 8276 10362
rect 8300 10310 8330 10362
rect 8330 10310 8342 10362
rect 8342 10310 8356 10362
rect 8380 10310 8394 10362
rect 8394 10310 8406 10362
rect 8406 10310 8436 10362
rect 8460 10310 8470 10362
rect 8470 10310 8516 10362
rect 8220 10308 8276 10310
rect 8300 10308 8356 10310
rect 8380 10308 8436 10310
rect 8460 10308 8516 10310
rect 8900 9818 8956 9820
rect 8980 9818 9036 9820
rect 9060 9818 9116 9820
rect 9140 9818 9196 9820
rect 8900 9766 8946 9818
rect 8946 9766 8956 9818
rect 8980 9766 9010 9818
rect 9010 9766 9022 9818
rect 9022 9766 9036 9818
rect 9060 9766 9074 9818
rect 9074 9766 9086 9818
rect 9086 9766 9116 9818
rect 9140 9766 9150 9818
rect 9150 9766 9196 9818
rect 8900 9764 8956 9766
rect 8980 9764 9036 9766
rect 9060 9764 9116 9766
rect 9140 9764 9196 9766
rect 8206 9580 8262 9616
rect 8206 9560 8208 9580
rect 8208 9560 8260 9580
rect 8260 9560 8262 9580
rect 8220 9274 8276 9276
rect 8300 9274 8356 9276
rect 8380 9274 8436 9276
rect 8460 9274 8516 9276
rect 8220 9222 8266 9274
rect 8266 9222 8276 9274
rect 8300 9222 8330 9274
rect 8330 9222 8342 9274
rect 8342 9222 8356 9274
rect 8380 9222 8394 9274
rect 8394 9222 8406 9274
rect 8406 9222 8436 9274
rect 8460 9222 8470 9274
rect 8470 9222 8516 9274
rect 8220 9220 8276 9222
rect 8300 9220 8356 9222
rect 8380 9220 8436 9222
rect 8460 9220 8516 9222
rect 8220 8186 8276 8188
rect 8300 8186 8356 8188
rect 8380 8186 8436 8188
rect 8460 8186 8516 8188
rect 8220 8134 8266 8186
rect 8266 8134 8276 8186
rect 8300 8134 8330 8186
rect 8330 8134 8342 8186
rect 8342 8134 8356 8186
rect 8380 8134 8394 8186
rect 8394 8134 8406 8186
rect 8406 8134 8436 8186
rect 8460 8134 8470 8186
rect 8470 8134 8516 8186
rect 8220 8132 8276 8134
rect 8300 8132 8356 8134
rect 8380 8132 8436 8134
rect 8460 8132 8516 8134
rect 8220 7098 8276 7100
rect 8300 7098 8356 7100
rect 8380 7098 8436 7100
rect 8460 7098 8516 7100
rect 8220 7046 8266 7098
rect 8266 7046 8276 7098
rect 8300 7046 8330 7098
rect 8330 7046 8342 7098
rect 8342 7046 8356 7098
rect 8380 7046 8394 7098
rect 8394 7046 8406 7098
rect 8406 7046 8436 7098
rect 8460 7046 8470 7098
rect 8470 7046 8516 7098
rect 8220 7044 8276 7046
rect 8300 7044 8356 7046
rect 8380 7044 8436 7046
rect 8460 7044 8516 7046
rect 6220 3834 6276 3836
rect 6300 3834 6356 3836
rect 6380 3834 6436 3836
rect 6460 3834 6516 3836
rect 6220 3782 6266 3834
rect 6266 3782 6276 3834
rect 6300 3782 6330 3834
rect 6330 3782 6342 3834
rect 6342 3782 6356 3834
rect 6380 3782 6394 3834
rect 6394 3782 6406 3834
rect 6406 3782 6436 3834
rect 6460 3782 6470 3834
rect 6470 3782 6516 3834
rect 6220 3780 6276 3782
rect 6300 3780 6356 3782
rect 6380 3780 6436 3782
rect 6460 3780 6516 3782
rect 6900 4378 6956 4380
rect 6980 4378 7036 4380
rect 7060 4378 7116 4380
rect 7140 4378 7196 4380
rect 6900 4326 6946 4378
rect 6946 4326 6956 4378
rect 6980 4326 7010 4378
rect 7010 4326 7022 4378
rect 7022 4326 7036 4378
rect 7060 4326 7074 4378
rect 7074 4326 7086 4378
rect 7086 4326 7116 4378
rect 7140 4326 7150 4378
rect 7150 4326 7196 4378
rect 6900 4324 6956 4326
rect 6980 4324 7036 4326
rect 7060 4324 7116 4326
rect 7140 4324 7196 4326
rect 8220 6010 8276 6012
rect 8300 6010 8356 6012
rect 8380 6010 8436 6012
rect 8460 6010 8516 6012
rect 8220 5958 8266 6010
rect 8266 5958 8276 6010
rect 8300 5958 8330 6010
rect 8330 5958 8342 6010
rect 8342 5958 8356 6010
rect 8380 5958 8394 6010
rect 8394 5958 8406 6010
rect 8406 5958 8436 6010
rect 8460 5958 8470 6010
rect 8470 5958 8516 6010
rect 8220 5956 8276 5958
rect 8300 5956 8356 5958
rect 8380 5956 8436 5958
rect 8460 5956 8516 5958
rect 8574 5208 8630 5264
rect 8482 5072 8538 5128
rect 8220 4922 8276 4924
rect 8300 4922 8356 4924
rect 8380 4922 8436 4924
rect 8460 4922 8516 4924
rect 8220 4870 8266 4922
rect 8266 4870 8276 4922
rect 8300 4870 8330 4922
rect 8330 4870 8342 4922
rect 8342 4870 8356 4922
rect 8380 4870 8394 4922
rect 8394 4870 8406 4922
rect 8406 4870 8436 4922
rect 8460 4870 8470 4922
rect 8470 4870 8516 4922
rect 8220 4868 8276 4870
rect 8300 4868 8356 4870
rect 8380 4868 8436 4870
rect 8460 4868 8516 4870
rect 8482 4120 8538 4176
rect 8220 3834 8276 3836
rect 8300 3834 8356 3836
rect 8380 3834 8436 3836
rect 8460 3834 8516 3836
rect 8220 3782 8266 3834
rect 8266 3782 8276 3834
rect 8300 3782 8330 3834
rect 8330 3782 8342 3834
rect 8342 3782 8356 3834
rect 8380 3782 8394 3834
rect 8394 3782 8406 3834
rect 8406 3782 8436 3834
rect 8460 3782 8470 3834
rect 8470 3782 8516 3834
rect 8220 3780 8276 3782
rect 8300 3780 8356 3782
rect 8380 3780 8436 3782
rect 8460 3780 8516 3782
rect 6900 3290 6956 3292
rect 6980 3290 7036 3292
rect 7060 3290 7116 3292
rect 7140 3290 7196 3292
rect 6900 3238 6946 3290
rect 6946 3238 6956 3290
rect 6980 3238 7010 3290
rect 7010 3238 7022 3290
rect 7022 3238 7036 3290
rect 7060 3238 7074 3290
rect 7074 3238 7086 3290
rect 7086 3238 7116 3290
rect 7140 3238 7150 3290
rect 7150 3238 7196 3290
rect 6900 3236 6956 3238
rect 6980 3236 7036 3238
rect 7060 3236 7116 3238
rect 7140 3236 7196 3238
rect 6220 2746 6276 2748
rect 6300 2746 6356 2748
rect 6380 2746 6436 2748
rect 6460 2746 6516 2748
rect 6220 2694 6266 2746
rect 6266 2694 6276 2746
rect 6300 2694 6330 2746
rect 6330 2694 6342 2746
rect 6342 2694 6356 2746
rect 6380 2694 6394 2746
rect 6394 2694 6406 2746
rect 6406 2694 6436 2746
rect 6460 2694 6470 2746
rect 6470 2694 6516 2746
rect 6220 2692 6276 2694
rect 6300 2692 6356 2694
rect 6380 2692 6436 2694
rect 6460 2692 6516 2694
rect 8900 8730 8956 8732
rect 8980 8730 9036 8732
rect 9060 8730 9116 8732
rect 9140 8730 9196 8732
rect 8900 8678 8946 8730
rect 8946 8678 8956 8730
rect 8980 8678 9010 8730
rect 9010 8678 9022 8730
rect 9022 8678 9036 8730
rect 9060 8678 9074 8730
rect 9074 8678 9086 8730
rect 9086 8678 9116 8730
rect 9140 8678 9150 8730
rect 9150 8678 9196 8730
rect 8900 8676 8956 8678
rect 8980 8676 9036 8678
rect 9060 8676 9116 8678
rect 9140 8676 9196 8678
rect 10782 13640 10838 13696
rect 10598 12960 10654 13016
rect 10220 12538 10276 12540
rect 10300 12538 10356 12540
rect 10380 12538 10436 12540
rect 10460 12538 10516 12540
rect 10220 12486 10266 12538
rect 10266 12486 10276 12538
rect 10300 12486 10330 12538
rect 10330 12486 10342 12538
rect 10342 12486 10356 12538
rect 10380 12486 10394 12538
rect 10394 12486 10406 12538
rect 10406 12486 10436 12538
rect 10460 12486 10470 12538
rect 10470 12486 10516 12538
rect 10220 12484 10276 12486
rect 10300 12484 10356 12486
rect 10380 12484 10436 12486
rect 10460 12484 10516 12486
rect 10220 11450 10276 11452
rect 10300 11450 10356 11452
rect 10380 11450 10436 11452
rect 10460 11450 10516 11452
rect 10220 11398 10266 11450
rect 10266 11398 10276 11450
rect 10300 11398 10330 11450
rect 10330 11398 10342 11450
rect 10342 11398 10356 11450
rect 10380 11398 10394 11450
rect 10394 11398 10406 11450
rect 10406 11398 10436 11450
rect 10460 11398 10470 11450
rect 10470 11398 10516 11450
rect 10220 11396 10276 11398
rect 10300 11396 10356 11398
rect 10380 11396 10436 11398
rect 10460 11396 10516 11398
rect 9310 10104 9366 10160
rect 10220 10362 10276 10364
rect 10300 10362 10356 10364
rect 10380 10362 10436 10364
rect 10460 10362 10516 10364
rect 10220 10310 10266 10362
rect 10266 10310 10276 10362
rect 10300 10310 10330 10362
rect 10330 10310 10342 10362
rect 10342 10310 10356 10362
rect 10380 10310 10394 10362
rect 10394 10310 10406 10362
rect 10406 10310 10436 10362
rect 10460 10310 10470 10362
rect 10470 10310 10516 10362
rect 10220 10308 10276 10310
rect 10300 10308 10356 10310
rect 10380 10308 10436 10310
rect 10460 10308 10516 10310
rect 8900 7642 8956 7644
rect 8980 7642 9036 7644
rect 9060 7642 9116 7644
rect 9140 7642 9196 7644
rect 8900 7590 8946 7642
rect 8946 7590 8956 7642
rect 8980 7590 9010 7642
rect 9010 7590 9022 7642
rect 9022 7590 9036 7642
rect 9060 7590 9074 7642
rect 9074 7590 9086 7642
rect 9086 7590 9116 7642
rect 9140 7590 9150 7642
rect 9150 7590 9196 7642
rect 8900 7588 8956 7590
rect 8980 7588 9036 7590
rect 9060 7588 9116 7590
rect 9140 7588 9196 7590
rect 8942 6840 8998 6896
rect 8900 6554 8956 6556
rect 8980 6554 9036 6556
rect 9060 6554 9116 6556
rect 9140 6554 9196 6556
rect 8900 6502 8946 6554
rect 8946 6502 8956 6554
rect 8980 6502 9010 6554
rect 9010 6502 9022 6554
rect 9022 6502 9036 6554
rect 9060 6502 9074 6554
rect 9074 6502 9086 6554
rect 9086 6502 9116 6554
rect 9140 6502 9150 6554
rect 9150 6502 9196 6554
rect 8900 6500 8956 6502
rect 8980 6500 9036 6502
rect 9060 6500 9116 6502
rect 9140 6500 9196 6502
rect 8900 5466 8956 5468
rect 8980 5466 9036 5468
rect 9060 5466 9116 5468
rect 9140 5466 9196 5468
rect 8900 5414 8946 5466
rect 8946 5414 8956 5466
rect 8980 5414 9010 5466
rect 9010 5414 9022 5466
rect 9022 5414 9036 5466
rect 9060 5414 9074 5466
rect 9074 5414 9086 5466
rect 9086 5414 9116 5466
rect 9140 5414 9150 5466
rect 9150 5414 9196 5466
rect 8900 5412 8956 5414
rect 8980 5412 9036 5414
rect 9060 5412 9116 5414
rect 9140 5412 9196 5414
rect 8900 4378 8956 4380
rect 8980 4378 9036 4380
rect 9060 4378 9116 4380
rect 9140 4378 9196 4380
rect 8900 4326 8946 4378
rect 8946 4326 8956 4378
rect 8980 4326 9010 4378
rect 9010 4326 9022 4378
rect 9022 4326 9036 4378
rect 9060 4326 9074 4378
rect 9074 4326 9086 4378
rect 9086 4326 9116 4378
rect 9140 4326 9150 4378
rect 9150 4326 9196 4378
rect 8900 4324 8956 4326
rect 8980 4324 9036 4326
rect 9060 4324 9116 4326
rect 9140 4324 9196 4326
rect 10220 9274 10276 9276
rect 10300 9274 10356 9276
rect 10380 9274 10436 9276
rect 10460 9274 10516 9276
rect 10220 9222 10266 9274
rect 10266 9222 10276 9274
rect 10300 9222 10330 9274
rect 10330 9222 10342 9274
rect 10342 9222 10356 9274
rect 10380 9222 10394 9274
rect 10394 9222 10406 9274
rect 10406 9222 10436 9274
rect 10460 9222 10470 9274
rect 10470 9222 10516 9274
rect 10220 9220 10276 9222
rect 10300 9220 10356 9222
rect 10380 9220 10436 9222
rect 10460 9220 10516 9222
rect 10220 8186 10276 8188
rect 10300 8186 10356 8188
rect 10380 8186 10436 8188
rect 10460 8186 10516 8188
rect 10220 8134 10266 8186
rect 10266 8134 10276 8186
rect 10300 8134 10330 8186
rect 10330 8134 10342 8186
rect 10342 8134 10356 8186
rect 10380 8134 10394 8186
rect 10394 8134 10406 8186
rect 10406 8134 10436 8186
rect 10460 8134 10470 8186
rect 10470 8134 10516 8186
rect 10220 8132 10276 8134
rect 10300 8132 10356 8134
rect 10380 8132 10436 8134
rect 10460 8132 10516 8134
rect 10782 12280 10838 12336
rect 10900 11994 10956 11996
rect 10980 11994 11036 11996
rect 11060 11994 11116 11996
rect 11140 11994 11196 11996
rect 10900 11942 10946 11994
rect 10946 11942 10956 11994
rect 10980 11942 11010 11994
rect 11010 11942 11022 11994
rect 11022 11942 11036 11994
rect 11060 11942 11074 11994
rect 11074 11942 11086 11994
rect 11086 11942 11116 11994
rect 11140 11942 11150 11994
rect 11150 11942 11196 11994
rect 10900 11940 10956 11942
rect 10980 11940 11036 11942
rect 11060 11940 11116 11942
rect 11140 11940 11196 11942
rect 11242 11600 11298 11656
rect 10900 10906 10956 10908
rect 10980 10906 11036 10908
rect 11060 10906 11116 10908
rect 11140 10906 11196 10908
rect 10900 10854 10946 10906
rect 10946 10854 10956 10906
rect 10980 10854 11010 10906
rect 11010 10854 11022 10906
rect 11022 10854 11036 10906
rect 11060 10854 11074 10906
rect 11074 10854 11086 10906
rect 11086 10854 11116 10906
rect 11140 10854 11150 10906
rect 11150 10854 11196 10906
rect 10900 10852 10956 10854
rect 10980 10852 11036 10854
rect 11060 10852 11116 10854
rect 11140 10852 11196 10854
rect 11334 10920 11390 10976
rect 10900 9818 10956 9820
rect 10980 9818 11036 9820
rect 11060 9818 11116 9820
rect 11140 9818 11196 9820
rect 10900 9766 10946 9818
rect 10946 9766 10956 9818
rect 10980 9766 11010 9818
rect 11010 9766 11022 9818
rect 11022 9766 11036 9818
rect 11060 9766 11074 9818
rect 11074 9766 11086 9818
rect 11086 9766 11116 9818
rect 11140 9766 11150 9818
rect 11150 9766 11196 9818
rect 10900 9764 10956 9766
rect 10980 9764 11036 9766
rect 11060 9764 11116 9766
rect 11140 9764 11196 9766
rect 10966 8880 11022 8936
rect 10900 8730 10956 8732
rect 10980 8730 11036 8732
rect 11060 8730 11116 8732
rect 11140 8730 11196 8732
rect 10900 8678 10946 8730
rect 10946 8678 10956 8730
rect 10980 8678 11010 8730
rect 11010 8678 11022 8730
rect 11022 8678 11036 8730
rect 11060 8678 11074 8730
rect 11074 8678 11086 8730
rect 11086 8678 11116 8730
rect 11140 8678 11150 8730
rect 11150 8678 11196 8730
rect 10900 8676 10956 8678
rect 10980 8676 11036 8678
rect 11060 8676 11116 8678
rect 11140 8676 11196 8678
rect 10782 8200 10838 8256
rect 10220 7098 10276 7100
rect 10300 7098 10356 7100
rect 10380 7098 10436 7100
rect 10460 7098 10516 7100
rect 10220 7046 10266 7098
rect 10266 7046 10276 7098
rect 10300 7046 10330 7098
rect 10330 7046 10342 7098
rect 10342 7046 10356 7098
rect 10380 7046 10394 7098
rect 10394 7046 10406 7098
rect 10406 7046 10436 7098
rect 10460 7046 10470 7098
rect 10470 7046 10516 7098
rect 10220 7044 10276 7046
rect 10300 7044 10356 7046
rect 10380 7044 10436 7046
rect 10460 7044 10516 7046
rect 10900 7642 10956 7644
rect 10980 7642 11036 7644
rect 11060 7642 11116 7644
rect 11140 7642 11196 7644
rect 10900 7590 10946 7642
rect 10946 7590 10956 7642
rect 10980 7590 11010 7642
rect 11010 7590 11022 7642
rect 11022 7590 11036 7642
rect 11060 7590 11074 7642
rect 11074 7590 11086 7642
rect 11086 7590 11116 7642
rect 11140 7590 11150 7642
rect 11150 7590 11196 7642
rect 10900 7588 10956 7590
rect 10980 7588 11036 7590
rect 11060 7588 11116 7590
rect 11140 7588 11196 7590
rect 11334 7540 11390 7576
rect 11334 7520 11336 7540
rect 11336 7520 11388 7540
rect 11388 7520 11390 7540
rect 10900 6554 10956 6556
rect 10980 6554 11036 6556
rect 11060 6554 11116 6556
rect 11140 6554 11196 6556
rect 10900 6502 10946 6554
rect 10946 6502 10956 6554
rect 10980 6502 11010 6554
rect 11010 6502 11022 6554
rect 11022 6502 11036 6554
rect 11060 6502 11074 6554
rect 11074 6502 11086 6554
rect 11086 6502 11116 6554
rect 11140 6502 11150 6554
rect 11150 6502 11196 6554
rect 10900 6500 10956 6502
rect 10980 6500 11036 6502
rect 11060 6500 11116 6502
rect 11140 6500 11196 6502
rect 10220 6010 10276 6012
rect 10300 6010 10356 6012
rect 10380 6010 10436 6012
rect 10460 6010 10516 6012
rect 10220 5958 10266 6010
rect 10266 5958 10276 6010
rect 10300 5958 10330 6010
rect 10330 5958 10342 6010
rect 10342 5958 10356 6010
rect 10380 5958 10394 6010
rect 10394 5958 10406 6010
rect 10406 5958 10436 6010
rect 10460 5958 10470 6010
rect 10470 5958 10516 6010
rect 10220 5956 10276 5958
rect 10300 5956 10356 5958
rect 10380 5956 10436 5958
rect 10460 5956 10516 5958
rect 11426 6196 11428 6216
rect 11428 6196 11480 6216
rect 11480 6196 11482 6216
rect 11426 6160 11482 6196
rect 10900 5466 10956 5468
rect 10980 5466 11036 5468
rect 11060 5466 11116 5468
rect 11140 5466 11196 5468
rect 10900 5414 10946 5466
rect 10946 5414 10956 5466
rect 10980 5414 11010 5466
rect 11010 5414 11022 5466
rect 11022 5414 11036 5466
rect 11060 5414 11074 5466
rect 11074 5414 11086 5466
rect 11086 5414 11116 5466
rect 11140 5414 11150 5466
rect 11150 5414 11196 5466
rect 10900 5412 10956 5414
rect 10980 5412 11036 5414
rect 11060 5412 11116 5414
rect 11140 5412 11196 5414
rect 10220 4922 10276 4924
rect 10300 4922 10356 4924
rect 10380 4922 10436 4924
rect 10460 4922 10516 4924
rect 10220 4870 10266 4922
rect 10266 4870 10276 4922
rect 10300 4870 10330 4922
rect 10330 4870 10342 4922
rect 10342 4870 10356 4922
rect 10380 4870 10394 4922
rect 10394 4870 10406 4922
rect 10406 4870 10436 4922
rect 10460 4870 10470 4922
rect 10470 4870 10516 4922
rect 10220 4868 10276 4870
rect 10300 4868 10356 4870
rect 10380 4868 10436 4870
rect 10460 4868 10516 4870
rect 11426 5480 11482 5536
rect 10900 4378 10956 4380
rect 10980 4378 11036 4380
rect 11060 4378 11116 4380
rect 11140 4378 11196 4380
rect 10900 4326 10946 4378
rect 10946 4326 10956 4378
rect 10980 4326 11010 4378
rect 11010 4326 11022 4378
rect 11022 4326 11036 4378
rect 11060 4326 11074 4378
rect 11074 4326 11086 4378
rect 11086 4326 11116 4378
rect 11140 4326 11150 4378
rect 11150 4326 11196 4378
rect 10900 4324 10956 4326
rect 10980 4324 11036 4326
rect 11060 4324 11116 4326
rect 11140 4324 11196 4326
rect 11334 4800 11390 4856
rect 11242 4156 11244 4176
rect 11244 4156 11296 4176
rect 11296 4156 11298 4176
rect 11242 4120 11298 4156
rect 10220 3834 10276 3836
rect 10300 3834 10356 3836
rect 10380 3834 10436 3836
rect 10460 3834 10516 3836
rect 10220 3782 10266 3834
rect 10266 3782 10276 3834
rect 10300 3782 10330 3834
rect 10330 3782 10342 3834
rect 10342 3782 10356 3834
rect 10380 3782 10394 3834
rect 10394 3782 10406 3834
rect 10406 3782 10436 3834
rect 10460 3782 10470 3834
rect 10470 3782 10516 3834
rect 10220 3780 10276 3782
rect 10300 3780 10356 3782
rect 10380 3780 10436 3782
rect 10460 3780 10516 3782
rect 8942 3440 8998 3496
rect 11242 3440 11298 3496
rect 8900 3290 8956 3292
rect 8980 3290 9036 3292
rect 9060 3290 9116 3292
rect 9140 3290 9196 3292
rect 8900 3238 8946 3290
rect 8946 3238 8956 3290
rect 8980 3238 9010 3290
rect 9010 3238 9022 3290
rect 9022 3238 9036 3290
rect 9060 3238 9074 3290
rect 9074 3238 9086 3290
rect 9086 3238 9116 3290
rect 9140 3238 9150 3290
rect 9150 3238 9196 3290
rect 8900 3236 8956 3238
rect 8980 3236 9036 3238
rect 9060 3236 9116 3238
rect 9140 3236 9196 3238
rect 8220 2746 8276 2748
rect 8300 2746 8356 2748
rect 8380 2746 8436 2748
rect 8460 2746 8516 2748
rect 6900 2202 6956 2204
rect 6980 2202 7036 2204
rect 7060 2202 7116 2204
rect 7140 2202 7196 2204
rect 6900 2150 6946 2202
rect 6946 2150 6956 2202
rect 6980 2150 7010 2202
rect 7010 2150 7022 2202
rect 7022 2150 7036 2202
rect 7060 2150 7074 2202
rect 7074 2150 7086 2202
rect 7086 2150 7116 2202
rect 7140 2150 7150 2202
rect 7150 2150 7196 2202
rect 6900 2148 6956 2150
rect 6980 2148 7036 2150
rect 7060 2148 7116 2150
rect 7140 2148 7196 2150
rect 6734 1400 6790 1456
rect 2962 40 3018 96
rect 8220 2694 8266 2746
rect 8266 2694 8276 2746
rect 8300 2694 8330 2746
rect 8330 2694 8342 2746
rect 8342 2694 8356 2746
rect 8380 2694 8394 2746
rect 8394 2694 8406 2746
rect 8406 2694 8436 2746
rect 8460 2694 8470 2746
rect 8470 2694 8516 2746
rect 8220 2692 8276 2694
rect 8300 2692 8356 2694
rect 8380 2692 8436 2694
rect 8460 2692 8516 2694
rect 8900 2202 8956 2204
rect 8980 2202 9036 2204
rect 9060 2202 9116 2204
rect 9140 2202 9196 2204
rect 8900 2150 8946 2202
rect 8946 2150 8956 2202
rect 8980 2150 9010 2202
rect 9010 2150 9022 2202
rect 9022 2150 9036 2202
rect 9060 2150 9074 2202
rect 9074 2150 9086 2202
rect 9086 2150 9116 2202
rect 9140 2150 9150 2202
rect 9150 2150 9196 2202
rect 8900 2148 8956 2150
rect 8980 2148 9036 2150
rect 9060 2148 9116 2150
rect 9140 2148 9196 2150
rect 7286 720 7342 776
rect 10900 3290 10956 3292
rect 10980 3290 11036 3292
rect 11060 3290 11116 3292
rect 11140 3290 11196 3292
rect 10900 3238 10946 3290
rect 10946 3238 10956 3290
rect 10980 3238 11010 3290
rect 11010 3238 11022 3290
rect 11022 3238 11036 3290
rect 11060 3238 11074 3290
rect 11074 3238 11086 3290
rect 11086 3238 11116 3290
rect 11140 3238 11150 3290
rect 11150 3238 11196 3290
rect 10900 3236 10956 3238
rect 10980 3236 11036 3238
rect 11060 3236 11116 3238
rect 11140 3236 11196 3238
rect 11334 2760 11390 2816
rect 10220 2746 10276 2748
rect 10300 2746 10356 2748
rect 10380 2746 10436 2748
rect 10460 2746 10516 2748
rect 10220 2694 10266 2746
rect 10266 2694 10276 2746
rect 10300 2694 10330 2746
rect 10330 2694 10342 2746
rect 10342 2694 10356 2746
rect 10380 2694 10394 2746
rect 10394 2694 10406 2746
rect 10406 2694 10436 2746
rect 10460 2694 10470 2746
rect 10470 2694 10516 2746
rect 10220 2692 10276 2694
rect 10300 2692 10356 2694
rect 10380 2692 10436 2694
rect 10460 2692 10516 2694
rect 10900 2202 10956 2204
rect 10980 2202 11036 2204
rect 11060 2202 11116 2204
rect 11140 2202 11196 2204
rect 10900 2150 10946 2202
rect 10946 2150 10956 2202
rect 10980 2150 11010 2202
rect 11010 2150 11022 2202
rect 11022 2150 11036 2202
rect 11060 2150 11074 2202
rect 11074 2150 11086 2202
rect 11086 2150 11116 2202
rect 11140 2150 11150 2202
rect 11150 2150 11196 2202
rect 10900 2148 10956 2150
rect 10980 2148 11036 2150
rect 11060 2148 11116 2150
rect 11140 2148 11196 2150
rect 11426 2080 11482 2136
rect 9218 40 9274 96
<< metal3 >>
rect 0 15058 800 15088
rect 2957 15058 3023 15061
rect 0 15056 3023 15058
rect 0 15000 2962 15056
rect 3018 15000 3023 15056
rect 0 14998 3023 15000
rect 0 14968 800 14998
rect 2957 14995 3023 14998
rect 9213 15058 9279 15061
rect 12188 15058 12988 15088
rect 9213 15056 12988 15058
rect 9213 15000 9218 15056
rect 9274 15000 12988 15056
rect 9213 14998 12988 15000
rect 9213 14995 9279 14998
rect 12188 14968 12988 14998
rect 0 14378 800 14408
rect 2865 14378 2931 14381
rect 0 14376 2931 14378
rect 0 14320 2870 14376
rect 2926 14320 2931 14376
rect 0 14318 2931 14320
rect 0 14288 800 14318
rect 2865 14315 2931 14318
rect 8109 14378 8175 14381
rect 12188 14378 12988 14408
rect 8109 14376 12988 14378
rect 8109 14320 8114 14376
rect 8170 14320 12988 14376
rect 8109 14318 12988 14320
rect 8109 14315 8175 14318
rect 12188 14288 12988 14318
rect 0 13698 800 13728
rect 3141 13698 3207 13701
rect 0 13696 3207 13698
rect 0 13640 3146 13696
rect 3202 13640 3207 13696
rect 0 13638 3207 13640
rect 0 13608 800 13638
rect 3141 13635 3207 13638
rect 10777 13698 10843 13701
rect 12188 13698 12988 13728
rect 10777 13696 12988 13698
rect 10777 13640 10782 13696
rect 10838 13640 12988 13696
rect 10777 13638 12988 13640
rect 10777 13635 10843 13638
rect 12188 13608 12988 13638
rect 0 13018 800 13048
rect 2773 13018 2839 13021
rect 0 13016 2839 13018
rect 0 12960 2778 13016
rect 2834 12960 2839 13016
rect 0 12958 2839 12960
rect 0 12928 800 12958
rect 2773 12955 2839 12958
rect 10593 13018 10659 13021
rect 12188 13018 12988 13048
rect 10593 13016 12988 13018
rect 10593 12960 10598 13016
rect 10654 12960 12988 13016
rect 10593 12958 12988 12960
rect 10593 12955 10659 12958
rect 12188 12928 12988 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 6210 12544 6526 12545
rect 6210 12480 6216 12544
rect 6280 12480 6296 12544
rect 6360 12480 6376 12544
rect 6440 12480 6456 12544
rect 6520 12480 6526 12544
rect 6210 12479 6526 12480
rect 8210 12544 8526 12545
rect 8210 12480 8216 12544
rect 8280 12480 8296 12544
rect 8360 12480 8376 12544
rect 8440 12480 8456 12544
rect 8520 12480 8526 12544
rect 8210 12479 8526 12480
rect 10210 12544 10526 12545
rect 10210 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10526 12544
rect 10210 12479 10526 12480
rect 0 12338 800 12368
rect 3877 12338 3943 12341
rect 0 12336 3943 12338
rect 0 12280 3882 12336
rect 3938 12280 3943 12336
rect 0 12278 3943 12280
rect 0 12248 800 12278
rect 3877 12275 3943 12278
rect 10777 12338 10843 12341
rect 12188 12338 12988 12368
rect 10777 12336 12988 12338
rect 10777 12280 10782 12336
rect 10838 12280 12988 12336
rect 10777 12278 12988 12280
rect 10777 12275 10843 12278
rect 12188 12248 12988 12278
rect 4890 12000 5206 12001
rect 4890 11936 4896 12000
rect 4960 11936 4976 12000
rect 5040 11936 5056 12000
rect 5120 11936 5136 12000
rect 5200 11936 5206 12000
rect 4890 11935 5206 11936
rect 6890 12000 7206 12001
rect 6890 11936 6896 12000
rect 6960 11936 6976 12000
rect 7040 11936 7056 12000
rect 7120 11936 7136 12000
rect 7200 11936 7206 12000
rect 6890 11935 7206 11936
rect 8890 12000 9206 12001
rect 8890 11936 8896 12000
rect 8960 11936 8976 12000
rect 9040 11936 9056 12000
rect 9120 11936 9136 12000
rect 9200 11936 9206 12000
rect 8890 11935 9206 11936
rect 10890 12000 11206 12001
rect 10890 11936 10896 12000
rect 10960 11936 10976 12000
rect 11040 11936 11056 12000
rect 11120 11936 11136 12000
rect 11200 11936 11206 12000
rect 10890 11935 11206 11936
rect 0 11658 800 11688
rect 6085 11658 6151 11661
rect 0 11656 6151 11658
rect 0 11600 6090 11656
rect 6146 11600 6151 11656
rect 0 11598 6151 11600
rect 0 11568 800 11598
rect 6085 11595 6151 11598
rect 11237 11658 11303 11661
rect 12188 11658 12988 11688
rect 11237 11656 12988 11658
rect 11237 11600 11242 11656
rect 11298 11600 12988 11656
rect 11237 11598 12988 11600
rect 11237 11595 11303 11598
rect 12188 11568 12988 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 6210 11456 6526 11457
rect 6210 11392 6216 11456
rect 6280 11392 6296 11456
rect 6360 11392 6376 11456
rect 6440 11392 6456 11456
rect 6520 11392 6526 11456
rect 6210 11391 6526 11392
rect 8210 11456 8526 11457
rect 8210 11392 8216 11456
rect 8280 11392 8296 11456
rect 8360 11392 8376 11456
rect 8440 11392 8456 11456
rect 8520 11392 8526 11456
rect 8210 11391 8526 11392
rect 10210 11456 10526 11457
rect 10210 11392 10216 11456
rect 10280 11392 10296 11456
rect 10360 11392 10376 11456
rect 10440 11392 10456 11456
rect 10520 11392 10526 11456
rect 10210 11391 10526 11392
rect 0 10978 800 11008
rect 4613 10978 4679 10981
rect 0 10976 4679 10978
rect 0 10920 4618 10976
rect 4674 10920 4679 10976
rect 0 10918 4679 10920
rect 0 10888 800 10918
rect 4613 10915 4679 10918
rect 11329 10978 11395 10981
rect 12188 10978 12988 11008
rect 11329 10976 12988 10978
rect 11329 10920 11334 10976
rect 11390 10920 12988 10976
rect 11329 10918 12988 10920
rect 11329 10915 11395 10918
rect 4890 10912 5206 10913
rect 4890 10848 4896 10912
rect 4960 10848 4976 10912
rect 5040 10848 5056 10912
rect 5120 10848 5136 10912
rect 5200 10848 5206 10912
rect 4890 10847 5206 10848
rect 6890 10912 7206 10913
rect 6890 10848 6896 10912
rect 6960 10848 6976 10912
rect 7040 10848 7056 10912
rect 7120 10848 7136 10912
rect 7200 10848 7206 10912
rect 6890 10847 7206 10848
rect 8890 10912 9206 10913
rect 8890 10848 8896 10912
rect 8960 10848 8976 10912
rect 9040 10848 9056 10912
rect 9120 10848 9136 10912
rect 9200 10848 9206 10912
rect 8890 10847 9206 10848
rect 10890 10912 11206 10913
rect 10890 10848 10896 10912
rect 10960 10848 10976 10912
rect 11040 10848 11056 10912
rect 11120 10848 11136 10912
rect 11200 10848 11206 10912
rect 12188 10888 12988 10918
rect 10890 10847 11206 10848
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 6210 10368 6526 10369
rect 6210 10304 6216 10368
rect 6280 10304 6296 10368
rect 6360 10304 6376 10368
rect 6440 10304 6456 10368
rect 6520 10304 6526 10368
rect 6210 10303 6526 10304
rect 8210 10368 8526 10369
rect 8210 10304 8216 10368
rect 8280 10304 8296 10368
rect 8360 10304 8376 10368
rect 8440 10304 8456 10368
rect 8520 10304 8526 10368
rect 8210 10303 8526 10304
rect 10210 10368 10526 10369
rect 10210 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10526 10368
rect 10210 10303 10526 10304
rect 12188 10298 12988 10328
rect 0 10238 2790 10298
rect 0 10208 800 10238
rect 2730 10162 2790 10238
rect 10734 10238 12988 10298
rect 6729 10162 6795 10165
rect 2730 10160 6795 10162
rect 2730 10104 6734 10160
rect 6790 10104 6795 10160
rect 2730 10102 6795 10104
rect 6729 10099 6795 10102
rect 9305 10162 9371 10165
rect 10734 10162 10794 10238
rect 12188 10208 12988 10238
rect 9305 10160 10794 10162
rect 9305 10104 9310 10160
rect 9366 10104 10794 10160
rect 9305 10102 10794 10104
rect 9305 10099 9371 10102
rect 4890 9824 5206 9825
rect 4890 9760 4896 9824
rect 4960 9760 4976 9824
rect 5040 9760 5056 9824
rect 5120 9760 5136 9824
rect 5200 9760 5206 9824
rect 4890 9759 5206 9760
rect 6890 9824 7206 9825
rect 6890 9760 6896 9824
rect 6960 9760 6976 9824
rect 7040 9760 7056 9824
rect 7120 9760 7136 9824
rect 7200 9760 7206 9824
rect 6890 9759 7206 9760
rect 8890 9824 9206 9825
rect 8890 9760 8896 9824
rect 8960 9760 8976 9824
rect 9040 9760 9056 9824
rect 9120 9760 9136 9824
rect 9200 9760 9206 9824
rect 8890 9759 9206 9760
rect 10890 9824 11206 9825
rect 10890 9760 10896 9824
rect 10960 9760 10976 9824
rect 11040 9760 11056 9824
rect 11120 9760 11136 9824
rect 11200 9760 11206 9824
rect 10890 9759 11206 9760
rect 0 9618 800 9648
rect 4061 9618 4127 9621
rect 0 9616 4127 9618
rect 0 9560 4066 9616
rect 4122 9560 4127 9616
rect 0 9558 4127 9560
rect 0 9528 800 9558
rect 4061 9555 4127 9558
rect 8201 9618 8267 9621
rect 12188 9618 12988 9648
rect 8201 9616 12988 9618
rect 8201 9560 8206 9616
rect 8262 9560 12988 9616
rect 8201 9558 12988 9560
rect 8201 9555 8267 9558
rect 12188 9528 12988 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 6210 9280 6526 9281
rect 6210 9216 6216 9280
rect 6280 9216 6296 9280
rect 6360 9216 6376 9280
rect 6440 9216 6456 9280
rect 6520 9216 6526 9280
rect 6210 9215 6526 9216
rect 8210 9280 8526 9281
rect 8210 9216 8216 9280
rect 8280 9216 8296 9280
rect 8360 9216 8376 9280
rect 8440 9216 8456 9280
rect 8520 9216 8526 9280
rect 8210 9215 8526 9216
rect 10210 9280 10526 9281
rect 10210 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10526 9280
rect 10210 9215 10526 9216
rect 0 8938 800 8968
rect 1301 8938 1367 8941
rect 0 8936 1367 8938
rect 0 8880 1306 8936
rect 1362 8880 1367 8936
rect 0 8878 1367 8880
rect 0 8848 800 8878
rect 1301 8875 1367 8878
rect 10961 8938 11027 8941
rect 12188 8938 12988 8968
rect 10961 8936 12988 8938
rect 10961 8880 10966 8936
rect 11022 8880 12988 8936
rect 10961 8878 12988 8880
rect 10961 8875 11027 8878
rect 12188 8848 12988 8878
rect 4890 8736 5206 8737
rect 4890 8672 4896 8736
rect 4960 8672 4976 8736
rect 5040 8672 5056 8736
rect 5120 8672 5136 8736
rect 5200 8672 5206 8736
rect 4890 8671 5206 8672
rect 6890 8736 7206 8737
rect 6890 8672 6896 8736
rect 6960 8672 6976 8736
rect 7040 8672 7056 8736
rect 7120 8672 7136 8736
rect 7200 8672 7206 8736
rect 6890 8671 7206 8672
rect 8890 8736 9206 8737
rect 8890 8672 8896 8736
rect 8960 8672 8976 8736
rect 9040 8672 9056 8736
rect 9120 8672 9136 8736
rect 9200 8672 9206 8736
rect 8890 8671 9206 8672
rect 10890 8736 11206 8737
rect 10890 8672 10896 8736
rect 10960 8672 10976 8736
rect 11040 8672 11056 8736
rect 11120 8672 11136 8736
rect 11200 8672 11206 8736
rect 10890 8671 11206 8672
rect 0 8258 800 8288
rect 3877 8258 3943 8261
rect 0 8256 3943 8258
rect 0 8200 3882 8256
rect 3938 8200 3943 8256
rect 0 8198 3943 8200
rect 0 8168 800 8198
rect 3877 8195 3943 8198
rect 10777 8258 10843 8261
rect 12188 8258 12988 8288
rect 10777 8256 12988 8258
rect 10777 8200 10782 8256
rect 10838 8200 12988 8256
rect 10777 8198 12988 8200
rect 10777 8195 10843 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 6210 8192 6526 8193
rect 6210 8128 6216 8192
rect 6280 8128 6296 8192
rect 6360 8128 6376 8192
rect 6440 8128 6456 8192
rect 6520 8128 6526 8192
rect 6210 8127 6526 8128
rect 8210 8192 8526 8193
rect 8210 8128 8216 8192
rect 8280 8128 8296 8192
rect 8360 8128 8376 8192
rect 8440 8128 8456 8192
rect 8520 8128 8526 8192
rect 8210 8127 8526 8128
rect 10210 8192 10526 8193
rect 10210 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10526 8192
rect 12188 8168 12988 8198
rect 10210 8127 10526 8128
rect 4890 7648 5206 7649
rect 0 7578 800 7608
rect 4890 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5136 7648
rect 5200 7584 5206 7648
rect 4890 7583 5206 7584
rect 6890 7648 7206 7649
rect 6890 7584 6896 7648
rect 6960 7584 6976 7648
rect 7040 7584 7056 7648
rect 7120 7584 7136 7648
rect 7200 7584 7206 7648
rect 6890 7583 7206 7584
rect 8890 7648 9206 7649
rect 8890 7584 8896 7648
rect 8960 7584 8976 7648
rect 9040 7584 9056 7648
rect 9120 7584 9136 7648
rect 9200 7584 9206 7648
rect 8890 7583 9206 7584
rect 10890 7648 11206 7649
rect 10890 7584 10896 7648
rect 10960 7584 10976 7648
rect 11040 7584 11056 7648
rect 11120 7584 11136 7648
rect 11200 7584 11206 7648
rect 10890 7583 11206 7584
rect 2773 7578 2839 7581
rect 0 7576 2839 7578
rect 0 7520 2778 7576
rect 2834 7520 2839 7576
rect 0 7518 2839 7520
rect 0 7488 800 7518
rect 2773 7515 2839 7518
rect 11329 7578 11395 7581
rect 12188 7578 12988 7608
rect 11329 7576 12988 7578
rect 11329 7520 11334 7576
rect 11390 7520 12988 7576
rect 11329 7518 12988 7520
rect 11329 7515 11395 7518
rect 12188 7488 12988 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 6210 7104 6526 7105
rect 6210 7040 6216 7104
rect 6280 7040 6296 7104
rect 6360 7040 6376 7104
rect 6440 7040 6456 7104
rect 6520 7040 6526 7104
rect 6210 7039 6526 7040
rect 8210 7104 8526 7105
rect 8210 7040 8216 7104
rect 8280 7040 8296 7104
rect 8360 7040 8376 7104
rect 8440 7040 8456 7104
rect 8520 7040 8526 7104
rect 8210 7039 8526 7040
rect 10210 7104 10526 7105
rect 10210 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10526 7104
rect 10210 7039 10526 7040
rect 0 6898 800 6928
rect 1209 6898 1275 6901
rect 0 6896 1275 6898
rect 0 6840 1214 6896
rect 1270 6840 1275 6896
rect 0 6838 1275 6840
rect 0 6808 800 6838
rect 1209 6835 1275 6838
rect 8937 6898 9003 6901
rect 12188 6898 12988 6928
rect 8937 6896 12988 6898
rect 8937 6840 8942 6896
rect 8998 6840 12988 6896
rect 8937 6838 12988 6840
rect 8937 6835 9003 6838
rect 12188 6808 12988 6838
rect 4890 6560 5206 6561
rect 4890 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5136 6560
rect 5200 6496 5206 6560
rect 4890 6495 5206 6496
rect 6890 6560 7206 6561
rect 6890 6496 6896 6560
rect 6960 6496 6976 6560
rect 7040 6496 7056 6560
rect 7120 6496 7136 6560
rect 7200 6496 7206 6560
rect 6890 6495 7206 6496
rect 8890 6560 9206 6561
rect 8890 6496 8896 6560
rect 8960 6496 8976 6560
rect 9040 6496 9056 6560
rect 9120 6496 9136 6560
rect 9200 6496 9206 6560
rect 8890 6495 9206 6496
rect 10890 6560 11206 6561
rect 10890 6496 10896 6560
rect 10960 6496 10976 6560
rect 11040 6496 11056 6560
rect 11120 6496 11136 6560
rect 11200 6496 11206 6560
rect 10890 6495 11206 6496
rect 0 6218 800 6248
rect 3601 6218 3667 6221
rect 0 6216 3667 6218
rect 0 6160 3606 6216
rect 3662 6160 3667 6216
rect 0 6158 3667 6160
rect 0 6128 800 6158
rect 3601 6155 3667 6158
rect 11421 6218 11487 6221
rect 12188 6218 12988 6248
rect 11421 6216 12988 6218
rect 11421 6160 11426 6216
rect 11482 6160 12988 6216
rect 11421 6158 12988 6160
rect 11421 6155 11487 6158
rect 12188 6128 12988 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 6210 6016 6526 6017
rect 6210 5952 6216 6016
rect 6280 5952 6296 6016
rect 6360 5952 6376 6016
rect 6440 5952 6456 6016
rect 6520 5952 6526 6016
rect 6210 5951 6526 5952
rect 8210 6016 8526 6017
rect 8210 5952 8216 6016
rect 8280 5952 8296 6016
rect 8360 5952 8376 6016
rect 8440 5952 8456 6016
rect 8520 5952 8526 6016
rect 8210 5951 8526 5952
rect 10210 6016 10526 6017
rect 10210 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10526 6016
rect 10210 5951 10526 5952
rect 0 5538 800 5568
rect 11421 5538 11487 5541
rect 12188 5538 12988 5568
rect 0 5478 2790 5538
rect 0 5448 800 5478
rect 2730 5266 2790 5478
rect 11421 5536 12988 5538
rect 11421 5480 11426 5536
rect 11482 5480 12988 5536
rect 11421 5478 12988 5480
rect 11421 5475 11487 5478
rect 4890 5472 5206 5473
rect 4890 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5136 5472
rect 5200 5408 5206 5472
rect 4890 5407 5206 5408
rect 6890 5472 7206 5473
rect 6890 5408 6896 5472
rect 6960 5408 6976 5472
rect 7040 5408 7056 5472
rect 7120 5408 7136 5472
rect 7200 5408 7206 5472
rect 6890 5407 7206 5408
rect 8890 5472 9206 5473
rect 8890 5408 8896 5472
rect 8960 5408 8976 5472
rect 9040 5408 9056 5472
rect 9120 5408 9136 5472
rect 9200 5408 9206 5472
rect 8890 5407 9206 5408
rect 10890 5472 11206 5473
rect 10890 5408 10896 5472
rect 10960 5408 10976 5472
rect 11040 5408 11056 5472
rect 11120 5408 11136 5472
rect 11200 5408 11206 5472
rect 12188 5448 12988 5478
rect 10890 5407 11206 5408
rect 8569 5266 8635 5269
rect 2730 5264 8635 5266
rect 2730 5208 8574 5264
rect 8630 5208 8635 5264
rect 2730 5206 8635 5208
rect 8569 5203 8635 5206
rect 8477 5130 8543 5133
rect 2730 5128 8543 5130
rect 2730 5072 8482 5128
rect 8538 5072 8543 5128
rect 2730 5070 8543 5072
rect 0 4858 800 4888
rect 2730 4858 2790 5070
rect 8477 5067 8543 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 6210 4928 6526 4929
rect 6210 4864 6216 4928
rect 6280 4864 6296 4928
rect 6360 4864 6376 4928
rect 6440 4864 6456 4928
rect 6520 4864 6526 4928
rect 6210 4863 6526 4864
rect 8210 4928 8526 4929
rect 8210 4864 8216 4928
rect 8280 4864 8296 4928
rect 8360 4864 8376 4928
rect 8440 4864 8456 4928
rect 8520 4864 8526 4928
rect 8210 4863 8526 4864
rect 10210 4928 10526 4929
rect 10210 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10526 4928
rect 10210 4863 10526 4864
rect 0 4798 2790 4858
rect 11329 4858 11395 4861
rect 12188 4858 12988 4888
rect 11329 4856 12988 4858
rect 11329 4800 11334 4856
rect 11390 4800 12988 4856
rect 11329 4798 12988 4800
rect 0 4768 800 4798
rect 11329 4795 11395 4798
rect 12188 4768 12988 4798
rect 4890 4384 5206 4385
rect 4890 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5136 4384
rect 5200 4320 5206 4384
rect 4890 4319 5206 4320
rect 6890 4384 7206 4385
rect 6890 4320 6896 4384
rect 6960 4320 6976 4384
rect 7040 4320 7056 4384
rect 7120 4320 7136 4384
rect 7200 4320 7206 4384
rect 6890 4319 7206 4320
rect 8890 4384 9206 4385
rect 8890 4320 8896 4384
rect 8960 4320 8976 4384
rect 9040 4320 9056 4384
rect 9120 4320 9136 4384
rect 9200 4320 9206 4384
rect 8890 4319 9206 4320
rect 10890 4384 11206 4385
rect 10890 4320 10896 4384
rect 10960 4320 10976 4384
rect 11040 4320 11056 4384
rect 11120 4320 11136 4384
rect 11200 4320 11206 4384
rect 10890 4319 11206 4320
rect 0 4178 800 4208
rect 8477 4178 8543 4181
rect 0 4176 8543 4178
rect 0 4120 8482 4176
rect 8538 4120 8543 4176
rect 0 4118 8543 4120
rect 0 4088 800 4118
rect 8477 4115 8543 4118
rect 11237 4178 11303 4181
rect 12188 4178 12988 4208
rect 11237 4176 12988 4178
rect 11237 4120 11242 4176
rect 11298 4120 12988 4176
rect 11237 4118 12988 4120
rect 11237 4115 11303 4118
rect 12188 4088 12988 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 6210 3840 6526 3841
rect 6210 3776 6216 3840
rect 6280 3776 6296 3840
rect 6360 3776 6376 3840
rect 6440 3776 6456 3840
rect 6520 3776 6526 3840
rect 6210 3775 6526 3776
rect 8210 3840 8526 3841
rect 8210 3776 8216 3840
rect 8280 3776 8296 3840
rect 8360 3776 8376 3840
rect 8440 3776 8456 3840
rect 8520 3776 8526 3840
rect 8210 3775 8526 3776
rect 10210 3840 10526 3841
rect 10210 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10526 3840
rect 10210 3775 10526 3776
rect 0 3498 800 3528
rect 8937 3498 9003 3501
rect 0 3496 9003 3498
rect 0 3440 8942 3496
rect 8998 3440 9003 3496
rect 0 3438 9003 3440
rect 0 3408 800 3438
rect 8937 3435 9003 3438
rect 11237 3498 11303 3501
rect 12188 3498 12988 3528
rect 11237 3496 12988 3498
rect 11237 3440 11242 3496
rect 11298 3440 12988 3496
rect 11237 3438 12988 3440
rect 11237 3435 11303 3438
rect 12188 3408 12988 3438
rect 4890 3296 5206 3297
rect 4890 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5136 3296
rect 5200 3232 5206 3296
rect 4890 3231 5206 3232
rect 6890 3296 7206 3297
rect 6890 3232 6896 3296
rect 6960 3232 6976 3296
rect 7040 3232 7056 3296
rect 7120 3232 7136 3296
rect 7200 3232 7206 3296
rect 6890 3231 7206 3232
rect 8890 3296 9206 3297
rect 8890 3232 8896 3296
rect 8960 3232 8976 3296
rect 9040 3232 9056 3296
rect 9120 3232 9136 3296
rect 9200 3232 9206 3296
rect 8890 3231 9206 3232
rect 10890 3296 11206 3297
rect 10890 3232 10896 3296
rect 10960 3232 10976 3296
rect 11040 3232 11056 3296
rect 11120 3232 11136 3296
rect 11200 3232 11206 3296
rect 10890 3231 11206 3232
rect 4429 2954 4495 2957
rect 2730 2952 4495 2954
rect 2730 2896 4434 2952
rect 4490 2896 4495 2952
rect 2730 2894 4495 2896
rect 0 2818 800 2848
rect 2730 2818 2790 2894
rect 4429 2891 4495 2894
rect 0 2758 2790 2818
rect 11329 2818 11395 2821
rect 12188 2818 12988 2848
rect 11329 2816 12988 2818
rect 11329 2760 11334 2816
rect 11390 2760 12988 2816
rect 11329 2758 12988 2760
rect 0 2728 800 2758
rect 11329 2755 11395 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 6210 2752 6526 2753
rect 6210 2688 6216 2752
rect 6280 2688 6296 2752
rect 6360 2688 6376 2752
rect 6440 2688 6456 2752
rect 6520 2688 6526 2752
rect 6210 2687 6526 2688
rect 8210 2752 8526 2753
rect 8210 2688 8216 2752
rect 8280 2688 8296 2752
rect 8360 2688 8376 2752
rect 8440 2688 8456 2752
rect 8520 2688 8526 2752
rect 8210 2687 8526 2688
rect 10210 2752 10526 2753
rect 10210 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10526 2752
rect 12188 2728 12988 2758
rect 10210 2687 10526 2688
rect 5809 2410 5875 2413
rect 4294 2408 5875 2410
rect 4294 2352 5814 2408
rect 5870 2352 5875 2408
rect 4294 2350 5875 2352
rect 0 2138 800 2168
rect 4294 2138 4354 2350
rect 5809 2347 5875 2350
rect 4890 2208 5206 2209
rect 4890 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5136 2208
rect 5200 2144 5206 2208
rect 4890 2143 5206 2144
rect 6890 2208 7206 2209
rect 6890 2144 6896 2208
rect 6960 2144 6976 2208
rect 7040 2144 7056 2208
rect 7120 2144 7136 2208
rect 7200 2144 7206 2208
rect 6890 2143 7206 2144
rect 8890 2208 9206 2209
rect 8890 2144 8896 2208
rect 8960 2144 8976 2208
rect 9040 2144 9056 2208
rect 9120 2144 9136 2208
rect 9200 2144 9206 2208
rect 8890 2143 9206 2144
rect 10890 2208 11206 2209
rect 10890 2144 10896 2208
rect 10960 2144 10976 2208
rect 11040 2144 11056 2208
rect 11120 2144 11136 2208
rect 11200 2144 11206 2208
rect 10890 2143 11206 2144
rect 0 2078 4354 2138
rect 11421 2138 11487 2141
rect 12188 2138 12988 2168
rect 11421 2136 12988 2138
rect 11421 2080 11426 2136
rect 11482 2080 12988 2136
rect 11421 2078 12988 2080
rect 0 2048 800 2078
rect 11421 2075 11487 2078
rect 12188 2048 12988 2078
rect 0 1458 800 1488
rect 3877 1458 3943 1461
rect 0 1456 3943 1458
rect 0 1400 3882 1456
rect 3938 1400 3943 1456
rect 0 1398 3943 1400
rect 0 1368 800 1398
rect 3877 1395 3943 1398
rect 6729 1458 6795 1461
rect 12188 1458 12988 1488
rect 6729 1456 12988 1458
rect 6729 1400 6734 1456
rect 6790 1400 12988 1456
rect 6729 1398 12988 1400
rect 6729 1395 6795 1398
rect 12188 1368 12988 1398
rect 0 778 800 808
rect 2773 778 2839 781
rect 0 776 2839 778
rect 0 720 2778 776
rect 2834 720 2839 776
rect 0 718 2839 720
rect 0 688 800 718
rect 2773 715 2839 718
rect 7281 778 7347 781
rect 12188 778 12988 808
rect 7281 776 12988 778
rect 7281 720 7286 776
rect 7342 720 12988 776
rect 7281 718 12988 720
rect 7281 715 7347 718
rect 12188 688 12988 718
rect 0 98 800 128
rect 2957 98 3023 101
rect 0 96 3023 98
rect 0 40 2962 96
rect 3018 40 3023 96
rect 0 38 3023 40
rect 0 8 800 38
rect 2957 35 3023 38
rect 9213 98 9279 101
rect 12188 98 12988 128
rect 9213 96 12988 98
rect 9213 40 9218 96
rect 9274 40 12988 96
rect 9213 38 12988 40
rect 9213 35 9279 38
rect 12188 8 12988 38
<< via3 >>
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 6216 12540 6280 12544
rect 6216 12484 6220 12540
rect 6220 12484 6276 12540
rect 6276 12484 6280 12540
rect 6216 12480 6280 12484
rect 6296 12540 6360 12544
rect 6296 12484 6300 12540
rect 6300 12484 6356 12540
rect 6356 12484 6360 12540
rect 6296 12480 6360 12484
rect 6376 12540 6440 12544
rect 6376 12484 6380 12540
rect 6380 12484 6436 12540
rect 6436 12484 6440 12540
rect 6376 12480 6440 12484
rect 6456 12540 6520 12544
rect 6456 12484 6460 12540
rect 6460 12484 6516 12540
rect 6516 12484 6520 12540
rect 6456 12480 6520 12484
rect 8216 12540 8280 12544
rect 8216 12484 8220 12540
rect 8220 12484 8276 12540
rect 8276 12484 8280 12540
rect 8216 12480 8280 12484
rect 8296 12540 8360 12544
rect 8296 12484 8300 12540
rect 8300 12484 8356 12540
rect 8356 12484 8360 12540
rect 8296 12480 8360 12484
rect 8376 12540 8440 12544
rect 8376 12484 8380 12540
rect 8380 12484 8436 12540
rect 8436 12484 8440 12540
rect 8376 12480 8440 12484
rect 8456 12540 8520 12544
rect 8456 12484 8460 12540
rect 8460 12484 8516 12540
rect 8516 12484 8520 12540
rect 8456 12480 8520 12484
rect 10216 12540 10280 12544
rect 10216 12484 10220 12540
rect 10220 12484 10276 12540
rect 10276 12484 10280 12540
rect 10216 12480 10280 12484
rect 10296 12540 10360 12544
rect 10296 12484 10300 12540
rect 10300 12484 10356 12540
rect 10356 12484 10360 12540
rect 10296 12480 10360 12484
rect 10376 12540 10440 12544
rect 10376 12484 10380 12540
rect 10380 12484 10436 12540
rect 10436 12484 10440 12540
rect 10376 12480 10440 12484
rect 10456 12540 10520 12544
rect 10456 12484 10460 12540
rect 10460 12484 10516 12540
rect 10516 12484 10520 12540
rect 10456 12480 10520 12484
rect 4896 11996 4960 12000
rect 4896 11940 4900 11996
rect 4900 11940 4956 11996
rect 4956 11940 4960 11996
rect 4896 11936 4960 11940
rect 4976 11996 5040 12000
rect 4976 11940 4980 11996
rect 4980 11940 5036 11996
rect 5036 11940 5040 11996
rect 4976 11936 5040 11940
rect 5056 11996 5120 12000
rect 5056 11940 5060 11996
rect 5060 11940 5116 11996
rect 5116 11940 5120 11996
rect 5056 11936 5120 11940
rect 5136 11996 5200 12000
rect 5136 11940 5140 11996
rect 5140 11940 5196 11996
rect 5196 11940 5200 11996
rect 5136 11936 5200 11940
rect 6896 11996 6960 12000
rect 6896 11940 6900 11996
rect 6900 11940 6956 11996
rect 6956 11940 6960 11996
rect 6896 11936 6960 11940
rect 6976 11996 7040 12000
rect 6976 11940 6980 11996
rect 6980 11940 7036 11996
rect 7036 11940 7040 11996
rect 6976 11936 7040 11940
rect 7056 11996 7120 12000
rect 7056 11940 7060 11996
rect 7060 11940 7116 11996
rect 7116 11940 7120 11996
rect 7056 11936 7120 11940
rect 7136 11996 7200 12000
rect 7136 11940 7140 11996
rect 7140 11940 7196 11996
rect 7196 11940 7200 11996
rect 7136 11936 7200 11940
rect 8896 11996 8960 12000
rect 8896 11940 8900 11996
rect 8900 11940 8956 11996
rect 8956 11940 8960 11996
rect 8896 11936 8960 11940
rect 8976 11996 9040 12000
rect 8976 11940 8980 11996
rect 8980 11940 9036 11996
rect 9036 11940 9040 11996
rect 8976 11936 9040 11940
rect 9056 11996 9120 12000
rect 9056 11940 9060 11996
rect 9060 11940 9116 11996
rect 9116 11940 9120 11996
rect 9056 11936 9120 11940
rect 9136 11996 9200 12000
rect 9136 11940 9140 11996
rect 9140 11940 9196 11996
rect 9196 11940 9200 11996
rect 9136 11936 9200 11940
rect 10896 11996 10960 12000
rect 10896 11940 10900 11996
rect 10900 11940 10956 11996
rect 10956 11940 10960 11996
rect 10896 11936 10960 11940
rect 10976 11996 11040 12000
rect 10976 11940 10980 11996
rect 10980 11940 11036 11996
rect 11036 11940 11040 11996
rect 10976 11936 11040 11940
rect 11056 11996 11120 12000
rect 11056 11940 11060 11996
rect 11060 11940 11116 11996
rect 11116 11940 11120 11996
rect 11056 11936 11120 11940
rect 11136 11996 11200 12000
rect 11136 11940 11140 11996
rect 11140 11940 11196 11996
rect 11196 11940 11200 11996
rect 11136 11936 11200 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 6216 11452 6280 11456
rect 6216 11396 6220 11452
rect 6220 11396 6276 11452
rect 6276 11396 6280 11452
rect 6216 11392 6280 11396
rect 6296 11452 6360 11456
rect 6296 11396 6300 11452
rect 6300 11396 6356 11452
rect 6356 11396 6360 11452
rect 6296 11392 6360 11396
rect 6376 11452 6440 11456
rect 6376 11396 6380 11452
rect 6380 11396 6436 11452
rect 6436 11396 6440 11452
rect 6376 11392 6440 11396
rect 6456 11452 6520 11456
rect 6456 11396 6460 11452
rect 6460 11396 6516 11452
rect 6516 11396 6520 11452
rect 6456 11392 6520 11396
rect 8216 11452 8280 11456
rect 8216 11396 8220 11452
rect 8220 11396 8276 11452
rect 8276 11396 8280 11452
rect 8216 11392 8280 11396
rect 8296 11452 8360 11456
rect 8296 11396 8300 11452
rect 8300 11396 8356 11452
rect 8356 11396 8360 11452
rect 8296 11392 8360 11396
rect 8376 11452 8440 11456
rect 8376 11396 8380 11452
rect 8380 11396 8436 11452
rect 8436 11396 8440 11452
rect 8376 11392 8440 11396
rect 8456 11452 8520 11456
rect 8456 11396 8460 11452
rect 8460 11396 8516 11452
rect 8516 11396 8520 11452
rect 8456 11392 8520 11396
rect 10216 11452 10280 11456
rect 10216 11396 10220 11452
rect 10220 11396 10276 11452
rect 10276 11396 10280 11452
rect 10216 11392 10280 11396
rect 10296 11452 10360 11456
rect 10296 11396 10300 11452
rect 10300 11396 10356 11452
rect 10356 11396 10360 11452
rect 10296 11392 10360 11396
rect 10376 11452 10440 11456
rect 10376 11396 10380 11452
rect 10380 11396 10436 11452
rect 10436 11396 10440 11452
rect 10376 11392 10440 11396
rect 10456 11452 10520 11456
rect 10456 11396 10460 11452
rect 10460 11396 10516 11452
rect 10516 11396 10520 11452
rect 10456 11392 10520 11396
rect 4896 10908 4960 10912
rect 4896 10852 4900 10908
rect 4900 10852 4956 10908
rect 4956 10852 4960 10908
rect 4896 10848 4960 10852
rect 4976 10908 5040 10912
rect 4976 10852 4980 10908
rect 4980 10852 5036 10908
rect 5036 10852 5040 10908
rect 4976 10848 5040 10852
rect 5056 10908 5120 10912
rect 5056 10852 5060 10908
rect 5060 10852 5116 10908
rect 5116 10852 5120 10908
rect 5056 10848 5120 10852
rect 5136 10908 5200 10912
rect 5136 10852 5140 10908
rect 5140 10852 5196 10908
rect 5196 10852 5200 10908
rect 5136 10848 5200 10852
rect 6896 10908 6960 10912
rect 6896 10852 6900 10908
rect 6900 10852 6956 10908
rect 6956 10852 6960 10908
rect 6896 10848 6960 10852
rect 6976 10908 7040 10912
rect 6976 10852 6980 10908
rect 6980 10852 7036 10908
rect 7036 10852 7040 10908
rect 6976 10848 7040 10852
rect 7056 10908 7120 10912
rect 7056 10852 7060 10908
rect 7060 10852 7116 10908
rect 7116 10852 7120 10908
rect 7056 10848 7120 10852
rect 7136 10908 7200 10912
rect 7136 10852 7140 10908
rect 7140 10852 7196 10908
rect 7196 10852 7200 10908
rect 7136 10848 7200 10852
rect 8896 10908 8960 10912
rect 8896 10852 8900 10908
rect 8900 10852 8956 10908
rect 8956 10852 8960 10908
rect 8896 10848 8960 10852
rect 8976 10908 9040 10912
rect 8976 10852 8980 10908
rect 8980 10852 9036 10908
rect 9036 10852 9040 10908
rect 8976 10848 9040 10852
rect 9056 10908 9120 10912
rect 9056 10852 9060 10908
rect 9060 10852 9116 10908
rect 9116 10852 9120 10908
rect 9056 10848 9120 10852
rect 9136 10908 9200 10912
rect 9136 10852 9140 10908
rect 9140 10852 9196 10908
rect 9196 10852 9200 10908
rect 9136 10848 9200 10852
rect 10896 10908 10960 10912
rect 10896 10852 10900 10908
rect 10900 10852 10956 10908
rect 10956 10852 10960 10908
rect 10896 10848 10960 10852
rect 10976 10908 11040 10912
rect 10976 10852 10980 10908
rect 10980 10852 11036 10908
rect 11036 10852 11040 10908
rect 10976 10848 11040 10852
rect 11056 10908 11120 10912
rect 11056 10852 11060 10908
rect 11060 10852 11116 10908
rect 11116 10852 11120 10908
rect 11056 10848 11120 10852
rect 11136 10908 11200 10912
rect 11136 10852 11140 10908
rect 11140 10852 11196 10908
rect 11196 10852 11200 10908
rect 11136 10848 11200 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 6216 10364 6280 10368
rect 6216 10308 6220 10364
rect 6220 10308 6276 10364
rect 6276 10308 6280 10364
rect 6216 10304 6280 10308
rect 6296 10364 6360 10368
rect 6296 10308 6300 10364
rect 6300 10308 6356 10364
rect 6356 10308 6360 10364
rect 6296 10304 6360 10308
rect 6376 10364 6440 10368
rect 6376 10308 6380 10364
rect 6380 10308 6436 10364
rect 6436 10308 6440 10364
rect 6376 10304 6440 10308
rect 6456 10364 6520 10368
rect 6456 10308 6460 10364
rect 6460 10308 6516 10364
rect 6516 10308 6520 10364
rect 6456 10304 6520 10308
rect 8216 10364 8280 10368
rect 8216 10308 8220 10364
rect 8220 10308 8276 10364
rect 8276 10308 8280 10364
rect 8216 10304 8280 10308
rect 8296 10364 8360 10368
rect 8296 10308 8300 10364
rect 8300 10308 8356 10364
rect 8356 10308 8360 10364
rect 8296 10304 8360 10308
rect 8376 10364 8440 10368
rect 8376 10308 8380 10364
rect 8380 10308 8436 10364
rect 8436 10308 8440 10364
rect 8376 10304 8440 10308
rect 8456 10364 8520 10368
rect 8456 10308 8460 10364
rect 8460 10308 8516 10364
rect 8516 10308 8520 10364
rect 8456 10304 8520 10308
rect 10216 10364 10280 10368
rect 10216 10308 10220 10364
rect 10220 10308 10276 10364
rect 10276 10308 10280 10364
rect 10216 10304 10280 10308
rect 10296 10364 10360 10368
rect 10296 10308 10300 10364
rect 10300 10308 10356 10364
rect 10356 10308 10360 10364
rect 10296 10304 10360 10308
rect 10376 10364 10440 10368
rect 10376 10308 10380 10364
rect 10380 10308 10436 10364
rect 10436 10308 10440 10364
rect 10376 10304 10440 10308
rect 10456 10364 10520 10368
rect 10456 10308 10460 10364
rect 10460 10308 10516 10364
rect 10516 10308 10520 10364
rect 10456 10304 10520 10308
rect 4896 9820 4960 9824
rect 4896 9764 4900 9820
rect 4900 9764 4956 9820
rect 4956 9764 4960 9820
rect 4896 9760 4960 9764
rect 4976 9820 5040 9824
rect 4976 9764 4980 9820
rect 4980 9764 5036 9820
rect 5036 9764 5040 9820
rect 4976 9760 5040 9764
rect 5056 9820 5120 9824
rect 5056 9764 5060 9820
rect 5060 9764 5116 9820
rect 5116 9764 5120 9820
rect 5056 9760 5120 9764
rect 5136 9820 5200 9824
rect 5136 9764 5140 9820
rect 5140 9764 5196 9820
rect 5196 9764 5200 9820
rect 5136 9760 5200 9764
rect 6896 9820 6960 9824
rect 6896 9764 6900 9820
rect 6900 9764 6956 9820
rect 6956 9764 6960 9820
rect 6896 9760 6960 9764
rect 6976 9820 7040 9824
rect 6976 9764 6980 9820
rect 6980 9764 7036 9820
rect 7036 9764 7040 9820
rect 6976 9760 7040 9764
rect 7056 9820 7120 9824
rect 7056 9764 7060 9820
rect 7060 9764 7116 9820
rect 7116 9764 7120 9820
rect 7056 9760 7120 9764
rect 7136 9820 7200 9824
rect 7136 9764 7140 9820
rect 7140 9764 7196 9820
rect 7196 9764 7200 9820
rect 7136 9760 7200 9764
rect 8896 9820 8960 9824
rect 8896 9764 8900 9820
rect 8900 9764 8956 9820
rect 8956 9764 8960 9820
rect 8896 9760 8960 9764
rect 8976 9820 9040 9824
rect 8976 9764 8980 9820
rect 8980 9764 9036 9820
rect 9036 9764 9040 9820
rect 8976 9760 9040 9764
rect 9056 9820 9120 9824
rect 9056 9764 9060 9820
rect 9060 9764 9116 9820
rect 9116 9764 9120 9820
rect 9056 9760 9120 9764
rect 9136 9820 9200 9824
rect 9136 9764 9140 9820
rect 9140 9764 9196 9820
rect 9196 9764 9200 9820
rect 9136 9760 9200 9764
rect 10896 9820 10960 9824
rect 10896 9764 10900 9820
rect 10900 9764 10956 9820
rect 10956 9764 10960 9820
rect 10896 9760 10960 9764
rect 10976 9820 11040 9824
rect 10976 9764 10980 9820
rect 10980 9764 11036 9820
rect 11036 9764 11040 9820
rect 10976 9760 11040 9764
rect 11056 9820 11120 9824
rect 11056 9764 11060 9820
rect 11060 9764 11116 9820
rect 11116 9764 11120 9820
rect 11056 9760 11120 9764
rect 11136 9820 11200 9824
rect 11136 9764 11140 9820
rect 11140 9764 11196 9820
rect 11196 9764 11200 9820
rect 11136 9760 11200 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 6216 9276 6280 9280
rect 6216 9220 6220 9276
rect 6220 9220 6276 9276
rect 6276 9220 6280 9276
rect 6216 9216 6280 9220
rect 6296 9276 6360 9280
rect 6296 9220 6300 9276
rect 6300 9220 6356 9276
rect 6356 9220 6360 9276
rect 6296 9216 6360 9220
rect 6376 9276 6440 9280
rect 6376 9220 6380 9276
rect 6380 9220 6436 9276
rect 6436 9220 6440 9276
rect 6376 9216 6440 9220
rect 6456 9276 6520 9280
rect 6456 9220 6460 9276
rect 6460 9220 6516 9276
rect 6516 9220 6520 9276
rect 6456 9216 6520 9220
rect 8216 9276 8280 9280
rect 8216 9220 8220 9276
rect 8220 9220 8276 9276
rect 8276 9220 8280 9276
rect 8216 9216 8280 9220
rect 8296 9276 8360 9280
rect 8296 9220 8300 9276
rect 8300 9220 8356 9276
rect 8356 9220 8360 9276
rect 8296 9216 8360 9220
rect 8376 9276 8440 9280
rect 8376 9220 8380 9276
rect 8380 9220 8436 9276
rect 8436 9220 8440 9276
rect 8376 9216 8440 9220
rect 8456 9276 8520 9280
rect 8456 9220 8460 9276
rect 8460 9220 8516 9276
rect 8516 9220 8520 9276
rect 8456 9216 8520 9220
rect 10216 9276 10280 9280
rect 10216 9220 10220 9276
rect 10220 9220 10276 9276
rect 10276 9220 10280 9276
rect 10216 9216 10280 9220
rect 10296 9276 10360 9280
rect 10296 9220 10300 9276
rect 10300 9220 10356 9276
rect 10356 9220 10360 9276
rect 10296 9216 10360 9220
rect 10376 9276 10440 9280
rect 10376 9220 10380 9276
rect 10380 9220 10436 9276
rect 10436 9220 10440 9276
rect 10376 9216 10440 9220
rect 10456 9276 10520 9280
rect 10456 9220 10460 9276
rect 10460 9220 10516 9276
rect 10516 9220 10520 9276
rect 10456 9216 10520 9220
rect 4896 8732 4960 8736
rect 4896 8676 4900 8732
rect 4900 8676 4956 8732
rect 4956 8676 4960 8732
rect 4896 8672 4960 8676
rect 4976 8732 5040 8736
rect 4976 8676 4980 8732
rect 4980 8676 5036 8732
rect 5036 8676 5040 8732
rect 4976 8672 5040 8676
rect 5056 8732 5120 8736
rect 5056 8676 5060 8732
rect 5060 8676 5116 8732
rect 5116 8676 5120 8732
rect 5056 8672 5120 8676
rect 5136 8732 5200 8736
rect 5136 8676 5140 8732
rect 5140 8676 5196 8732
rect 5196 8676 5200 8732
rect 5136 8672 5200 8676
rect 6896 8732 6960 8736
rect 6896 8676 6900 8732
rect 6900 8676 6956 8732
rect 6956 8676 6960 8732
rect 6896 8672 6960 8676
rect 6976 8732 7040 8736
rect 6976 8676 6980 8732
rect 6980 8676 7036 8732
rect 7036 8676 7040 8732
rect 6976 8672 7040 8676
rect 7056 8732 7120 8736
rect 7056 8676 7060 8732
rect 7060 8676 7116 8732
rect 7116 8676 7120 8732
rect 7056 8672 7120 8676
rect 7136 8732 7200 8736
rect 7136 8676 7140 8732
rect 7140 8676 7196 8732
rect 7196 8676 7200 8732
rect 7136 8672 7200 8676
rect 8896 8732 8960 8736
rect 8896 8676 8900 8732
rect 8900 8676 8956 8732
rect 8956 8676 8960 8732
rect 8896 8672 8960 8676
rect 8976 8732 9040 8736
rect 8976 8676 8980 8732
rect 8980 8676 9036 8732
rect 9036 8676 9040 8732
rect 8976 8672 9040 8676
rect 9056 8732 9120 8736
rect 9056 8676 9060 8732
rect 9060 8676 9116 8732
rect 9116 8676 9120 8732
rect 9056 8672 9120 8676
rect 9136 8732 9200 8736
rect 9136 8676 9140 8732
rect 9140 8676 9196 8732
rect 9196 8676 9200 8732
rect 9136 8672 9200 8676
rect 10896 8732 10960 8736
rect 10896 8676 10900 8732
rect 10900 8676 10956 8732
rect 10956 8676 10960 8732
rect 10896 8672 10960 8676
rect 10976 8732 11040 8736
rect 10976 8676 10980 8732
rect 10980 8676 11036 8732
rect 11036 8676 11040 8732
rect 10976 8672 11040 8676
rect 11056 8732 11120 8736
rect 11056 8676 11060 8732
rect 11060 8676 11116 8732
rect 11116 8676 11120 8732
rect 11056 8672 11120 8676
rect 11136 8732 11200 8736
rect 11136 8676 11140 8732
rect 11140 8676 11196 8732
rect 11196 8676 11200 8732
rect 11136 8672 11200 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 6216 8188 6280 8192
rect 6216 8132 6220 8188
rect 6220 8132 6276 8188
rect 6276 8132 6280 8188
rect 6216 8128 6280 8132
rect 6296 8188 6360 8192
rect 6296 8132 6300 8188
rect 6300 8132 6356 8188
rect 6356 8132 6360 8188
rect 6296 8128 6360 8132
rect 6376 8188 6440 8192
rect 6376 8132 6380 8188
rect 6380 8132 6436 8188
rect 6436 8132 6440 8188
rect 6376 8128 6440 8132
rect 6456 8188 6520 8192
rect 6456 8132 6460 8188
rect 6460 8132 6516 8188
rect 6516 8132 6520 8188
rect 6456 8128 6520 8132
rect 8216 8188 8280 8192
rect 8216 8132 8220 8188
rect 8220 8132 8276 8188
rect 8276 8132 8280 8188
rect 8216 8128 8280 8132
rect 8296 8188 8360 8192
rect 8296 8132 8300 8188
rect 8300 8132 8356 8188
rect 8356 8132 8360 8188
rect 8296 8128 8360 8132
rect 8376 8188 8440 8192
rect 8376 8132 8380 8188
rect 8380 8132 8436 8188
rect 8436 8132 8440 8188
rect 8376 8128 8440 8132
rect 8456 8188 8520 8192
rect 8456 8132 8460 8188
rect 8460 8132 8516 8188
rect 8516 8132 8520 8188
rect 8456 8128 8520 8132
rect 10216 8188 10280 8192
rect 10216 8132 10220 8188
rect 10220 8132 10276 8188
rect 10276 8132 10280 8188
rect 10216 8128 10280 8132
rect 10296 8188 10360 8192
rect 10296 8132 10300 8188
rect 10300 8132 10356 8188
rect 10356 8132 10360 8188
rect 10296 8128 10360 8132
rect 10376 8188 10440 8192
rect 10376 8132 10380 8188
rect 10380 8132 10436 8188
rect 10436 8132 10440 8188
rect 10376 8128 10440 8132
rect 10456 8188 10520 8192
rect 10456 8132 10460 8188
rect 10460 8132 10516 8188
rect 10516 8132 10520 8188
rect 10456 8128 10520 8132
rect 4896 7644 4960 7648
rect 4896 7588 4900 7644
rect 4900 7588 4956 7644
rect 4956 7588 4960 7644
rect 4896 7584 4960 7588
rect 4976 7644 5040 7648
rect 4976 7588 4980 7644
rect 4980 7588 5036 7644
rect 5036 7588 5040 7644
rect 4976 7584 5040 7588
rect 5056 7644 5120 7648
rect 5056 7588 5060 7644
rect 5060 7588 5116 7644
rect 5116 7588 5120 7644
rect 5056 7584 5120 7588
rect 5136 7644 5200 7648
rect 5136 7588 5140 7644
rect 5140 7588 5196 7644
rect 5196 7588 5200 7644
rect 5136 7584 5200 7588
rect 6896 7644 6960 7648
rect 6896 7588 6900 7644
rect 6900 7588 6956 7644
rect 6956 7588 6960 7644
rect 6896 7584 6960 7588
rect 6976 7644 7040 7648
rect 6976 7588 6980 7644
rect 6980 7588 7036 7644
rect 7036 7588 7040 7644
rect 6976 7584 7040 7588
rect 7056 7644 7120 7648
rect 7056 7588 7060 7644
rect 7060 7588 7116 7644
rect 7116 7588 7120 7644
rect 7056 7584 7120 7588
rect 7136 7644 7200 7648
rect 7136 7588 7140 7644
rect 7140 7588 7196 7644
rect 7196 7588 7200 7644
rect 7136 7584 7200 7588
rect 8896 7644 8960 7648
rect 8896 7588 8900 7644
rect 8900 7588 8956 7644
rect 8956 7588 8960 7644
rect 8896 7584 8960 7588
rect 8976 7644 9040 7648
rect 8976 7588 8980 7644
rect 8980 7588 9036 7644
rect 9036 7588 9040 7644
rect 8976 7584 9040 7588
rect 9056 7644 9120 7648
rect 9056 7588 9060 7644
rect 9060 7588 9116 7644
rect 9116 7588 9120 7644
rect 9056 7584 9120 7588
rect 9136 7644 9200 7648
rect 9136 7588 9140 7644
rect 9140 7588 9196 7644
rect 9196 7588 9200 7644
rect 9136 7584 9200 7588
rect 10896 7644 10960 7648
rect 10896 7588 10900 7644
rect 10900 7588 10956 7644
rect 10956 7588 10960 7644
rect 10896 7584 10960 7588
rect 10976 7644 11040 7648
rect 10976 7588 10980 7644
rect 10980 7588 11036 7644
rect 11036 7588 11040 7644
rect 10976 7584 11040 7588
rect 11056 7644 11120 7648
rect 11056 7588 11060 7644
rect 11060 7588 11116 7644
rect 11116 7588 11120 7644
rect 11056 7584 11120 7588
rect 11136 7644 11200 7648
rect 11136 7588 11140 7644
rect 11140 7588 11196 7644
rect 11196 7588 11200 7644
rect 11136 7584 11200 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 6216 7100 6280 7104
rect 6216 7044 6220 7100
rect 6220 7044 6276 7100
rect 6276 7044 6280 7100
rect 6216 7040 6280 7044
rect 6296 7100 6360 7104
rect 6296 7044 6300 7100
rect 6300 7044 6356 7100
rect 6356 7044 6360 7100
rect 6296 7040 6360 7044
rect 6376 7100 6440 7104
rect 6376 7044 6380 7100
rect 6380 7044 6436 7100
rect 6436 7044 6440 7100
rect 6376 7040 6440 7044
rect 6456 7100 6520 7104
rect 6456 7044 6460 7100
rect 6460 7044 6516 7100
rect 6516 7044 6520 7100
rect 6456 7040 6520 7044
rect 8216 7100 8280 7104
rect 8216 7044 8220 7100
rect 8220 7044 8276 7100
rect 8276 7044 8280 7100
rect 8216 7040 8280 7044
rect 8296 7100 8360 7104
rect 8296 7044 8300 7100
rect 8300 7044 8356 7100
rect 8356 7044 8360 7100
rect 8296 7040 8360 7044
rect 8376 7100 8440 7104
rect 8376 7044 8380 7100
rect 8380 7044 8436 7100
rect 8436 7044 8440 7100
rect 8376 7040 8440 7044
rect 8456 7100 8520 7104
rect 8456 7044 8460 7100
rect 8460 7044 8516 7100
rect 8516 7044 8520 7100
rect 8456 7040 8520 7044
rect 10216 7100 10280 7104
rect 10216 7044 10220 7100
rect 10220 7044 10276 7100
rect 10276 7044 10280 7100
rect 10216 7040 10280 7044
rect 10296 7100 10360 7104
rect 10296 7044 10300 7100
rect 10300 7044 10356 7100
rect 10356 7044 10360 7100
rect 10296 7040 10360 7044
rect 10376 7100 10440 7104
rect 10376 7044 10380 7100
rect 10380 7044 10436 7100
rect 10436 7044 10440 7100
rect 10376 7040 10440 7044
rect 10456 7100 10520 7104
rect 10456 7044 10460 7100
rect 10460 7044 10516 7100
rect 10516 7044 10520 7100
rect 10456 7040 10520 7044
rect 4896 6556 4960 6560
rect 4896 6500 4900 6556
rect 4900 6500 4956 6556
rect 4956 6500 4960 6556
rect 4896 6496 4960 6500
rect 4976 6556 5040 6560
rect 4976 6500 4980 6556
rect 4980 6500 5036 6556
rect 5036 6500 5040 6556
rect 4976 6496 5040 6500
rect 5056 6556 5120 6560
rect 5056 6500 5060 6556
rect 5060 6500 5116 6556
rect 5116 6500 5120 6556
rect 5056 6496 5120 6500
rect 5136 6556 5200 6560
rect 5136 6500 5140 6556
rect 5140 6500 5196 6556
rect 5196 6500 5200 6556
rect 5136 6496 5200 6500
rect 6896 6556 6960 6560
rect 6896 6500 6900 6556
rect 6900 6500 6956 6556
rect 6956 6500 6960 6556
rect 6896 6496 6960 6500
rect 6976 6556 7040 6560
rect 6976 6500 6980 6556
rect 6980 6500 7036 6556
rect 7036 6500 7040 6556
rect 6976 6496 7040 6500
rect 7056 6556 7120 6560
rect 7056 6500 7060 6556
rect 7060 6500 7116 6556
rect 7116 6500 7120 6556
rect 7056 6496 7120 6500
rect 7136 6556 7200 6560
rect 7136 6500 7140 6556
rect 7140 6500 7196 6556
rect 7196 6500 7200 6556
rect 7136 6496 7200 6500
rect 8896 6556 8960 6560
rect 8896 6500 8900 6556
rect 8900 6500 8956 6556
rect 8956 6500 8960 6556
rect 8896 6496 8960 6500
rect 8976 6556 9040 6560
rect 8976 6500 8980 6556
rect 8980 6500 9036 6556
rect 9036 6500 9040 6556
rect 8976 6496 9040 6500
rect 9056 6556 9120 6560
rect 9056 6500 9060 6556
rect 9060 6500 9116 6556
rect 9116 6500 9120 6556
rect 9056 6496 9120 6500
rect 9136 6556 9200 6560
rect 9136 6500 9140 6556
rect 9140 6500 9196 6556
rect 9196 6500 9200 6556
rect 9136 6496 9200 6500
rect 10896 6556 10960 6560
rect 10896 6500 10900 6556
rect 10900 6500 10956 6556
rect 10956 6500 10960 6556
rect 10896 6496 10960 6500
rect 10976 6556 11040 6560
rect 10976 6500 10980 6556
rect 10980 6500 11036 6556
rect 11036 6500 11040 6556
rect 10976 6496 11040 6500
rect 11056 6556 11120 6560
rect 11056 6500 11060 6556
rect 11060 6500 11116 6556
rect 11116 6500 11120 6556
rect 11056 6496 11120 6500
rect 11136 6556 11200 6560
rect 11136 6500 11140 6556
rect 11140 6500 11196 6556
rect 11196 6500 11200 6556
rect 11136 6496 11200 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 6216 6012 6280 6016
rect 6216 5956 6220 6012
rect 6220 5956 6276 6012
rect 6276 5956 6280 6012
rect 6216 5952 6280 5956
rect 6296 6012 6360 6016
rect 6296 5956 6300 6012
rect 6300 5956 6356 6012
rect 6356 5956 6360 6012
rect 6296 5952 6360 5956
rect 6376 6012 6440 6016
rect 6376 5956 6380 6012
rect 6380 5956 6436 6012
rect 6436 5956 6440 6012
rect 6376 5952 6440 5956
rect 6456 6012 6520 6016
rect 6456 5956 6460 6012
rect 6460 5956 6516 6012
rect 6516 5956 6520 6012
rect 6456 5952 6520 5956
rect 8216 6012 8280 6016
rect 8216 5956 8220 6012
rect 8220 5956 8276 6012
rect 8276 5956 8280 6012
rect 8216 5952 8280 5956
rect 8296 6012 8360 6016
rect 8296 5956 8300 6012
rect 8300 5956 8356 6012
rect 8356 5956 8360 6012
rect 8296 5952 8360 5956
rect 8376 6012 8440 6016
rect 8376 5956 8380 6012
rect 8380 5956 8436 6012
rect 8436 5956 8440 6012
rect 8376 5952 8440 5956
rect 8456 6012 8520 6016
rect 8456 5956 8460 6012
rect 8460 5956 8516 6012
rect 8516 5956 8520 6012
rect 8456 5952 8520 5956
rect 10216 6012 10280 6016
rect 10216 5956 10220 6012
rect 10220 5956 10276 6012
rect 10276 5956 10280 6012
rect 10216 5952 10280 5956
rect 10296 6012 10360 6016
rect 10296 5956 10300 6012
rect 10300 5956 10356 6012
rect 10356 5956 10360 6012
rect 10296 5952 10360 5956
rect 10376 6012 10440 6016
rect 10376 5956 10380 6012
rect 10380 5956 10436 6012
rect 10436 5956 10440 6012
rect 10376 5952 10440 5956
rect 10456 6012 10520 6016
rect 10456 5956 10460 6012
rect 10460 5956 10516 6012
rect 10516 5956 10520 6012
rect 10456 5952 10520 5956
rect 4896 5468 4960 5472
rect 4896 5412 4900 5468
rect 4900 5412 4956 5468
rect 4956 5412 4960 5468
rect 4896 5408 4960 5412
rect 4976 5468 5040 5472
rect 4976 5412 4980 5468
rect 4980 5412 5036 5468
rect 5036 5412 5040 5468
rect 4976 5408 5040 5412
rect 5056 5468 5120 5472
rect 5056 5412 5060 5468
rect 5060 5412 5116 5468
rect 5116 5412 5120 5468
rect 5056 5408 5120 5412
rect 5136 5468 5200 5472
rect 5136 5412 5140 5468
rect 5140 5412 5196 5468
rect 5196 5412 5200 5468
rect 5136 5408 5200 5412
rect 6896 5468 6960 5472
rect 6896 5412 6900 5468
rect 6900 5412 6956 5468
rect 6956 5412 6960 5468
rect 6896 5408 6960 5412
rect 6976 5468 7040 5472
rect 6976 5412 6980 5468
rect 6980 5412 7036 5468
rect 7036 5412 7040 5468
rect 6976 5408 7040 5412
rect 7056 5468 7120 5472
rect 7056 5412 7060 5468
rect 7060 5412 7116 5468
rect 7116 5412 7120 5468
rect 7056 5408 7120 5412
rect 7136 5468 7200 5472
rect 7136 5412 7140 5468
rect 7140 5412 7196 5468
rect 7196 5412 7200 5468
rect 7136 5408 7200 5412
rect 8896 5468 8960 5472
rect 8896 5412 8900 5468
rect 8900 5412 8956 5468
rect 8956 5412 8960 5468
rect 8896 5408 8960 5412
rect 8976 5468 9040 5472
rect 8976 5412 8980 5468
rect 8980 5412 9036 5468
rect 9036 5412 9040 5468
rect 8976 5408 9040 5412
rect 9056 5468 9120 5472
rect 9056 5412 9060 5468
rect 9060 5412 9116 5468
rect 9116 5412 9120 5468
rect 9056 5408 9120 5412
rect 9136 5468 9200 5472
rect 9136 5412 9140 5468
rect 9140 5412 9196 5468
rect 9196 5412 9200 5468
rect 9136 5408 9200 5412
rect 10896 5468 10960 5472
rect 10896 5412 10900 5468
rect 10900 5412 10956 5468
rect 10956 5412 10960 5468
rect 10896 5408 10960 5412
rect 10976 5468 11040 5472
rect 10976 5412 10980 5468
rect 10980 5412 11036 5468
rect 11036 5412 11040 5468
rect 10976 5408 11040 5412
rect 11056 5468 11120 5472
rect 11056 5412 11060 5468
rect 11060 5412 11116 5468
rect 11116 5412 11120 5468
rect 11056 5408 11120 5412
rect 11136 5468 11200 5472
rect 11136 5412 11140 5468
rect 11140 5412 11196 5468
rect 11196 5412 11200 5468
rect 11136 5408 11200 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 6216 4924 6280 4928
rect 6216 4868 6220 4924
rect 6220 4868 6276 4924
rect 6276 4868 6280 4924
rect 6216 4864 6280 4868
rect 6296 4924 6360 4928
rect 6296 4868 6300 4924
rect 6300 4868 6356 4924
rect 6356 4868 6360 4924
rect 6296 4864 6360 4868
rect 6376 4924 6440 4928
rect 6376 4868 6380 4924
rect 6380 4868 6436 4924
rect 6436 4868 6440 4924
rect 6376 4864 6440 4868
rect 6456 4924 6520 4928
rect 6456 4868 6460 4924
rect 6460 4868 6516 4924
rect 6516 4868 6520 4924
rect 6456 4864 6520 4868
rect 8216 4924 8280 4928
rect 8216 4868 8220 4924
rect 8220 4868 8276 4924
rect 8276 4868 8280 4924
rect 8216 4864 8280 4868
rect 8296 4924 8360 4928
rect 8296 4868 8300 4924
rect 8300 4868 8356 4924
rect 8356 4868 8360 4924
rect 8296 4864 8360 4868
rect 8376 4924 8440 4928
rect 8376 4868 8380 4924
rect 8380 4868 8436 4924
rect 8436 4868 8440 4924
rect 8376 4864 8440 4868
rect 8456 4924 8520 4928
rect 8456 4868 8460 4924
rect 8460 4868 8516 4924
rect 8516 4868 8520 4924
rect 8456 4864 8520 4868
rect 10216 4924 10280 4928
rect 10216 4868 10220 4924
rect 10220 4868 10276 4924
rect 10276 4868 10280 4924
rect 10216 4864 10280 4868
rect 10296 4924 10360 4928
rect 10296 4868 10300 4924
rect 10300 4868 10356 4924
rect 10356 4868 10360 4924
rect 10296 4864 10360 4868
rect 10376 4924 10440 4928
rect 10376 4868 10380 4924
rect 10380 4868 10436 4924
rect 10436 4868 10440 4924
rect 10376 4864 10440 4868
rect 10456 4924 10520 4928
rect 10456 4868 10460 4924
rect 10460 4868 10516 4924
rect 10516 4868 10520 4924
rect 10456 4864 10520 4868
rect 4896 4380 4960 4384
rect 4896 4324 4900 4380
rect 4900 4324 4956 4380
rect 4956 4324 4960 4380
rect 4896 4320 4960 4324
rect 4976 4380 5040 4384
rect 4976 4324 4980 4380
rect 4980 4324 5036 4380
rect 5036 4324 5040 4380
rect 4976 4320 5040 4324
rect 5056 4380 5120 4384
rect 5056 4324 5060 4380
rect 5060 4324 5116 4380
rect 5116 4324 5120 4380
rect 5056 4320 5120 4324
rect 5136 4380 5200 4384
rect 5136 4324 5140 4380
rect 5140 4324 5196 4380
rect 5196 4324 5200 4380
rect 5136 4320 5200 4324
rect 6896 4380 6960 4384
rect 6896 4324 6900 4380
rect 6900 4324 6956 4380
rect 6956 4324 6960 4380
rect 6896 4320 6960 4324
rect 6976 4380 7040 4384
rect 6976 4324 6980 4380
rect 6980 4324 7036 4380
rect 7036 4324 7040 4380
rect 6976 4320 7040 4324
rect 7056 4380 7120 4384
rect 7056 4324 7060 4380
rect 7060 4324 7116 4380
rect 7116 4324 7120 4380
rect 7056 4320 7120 4324
rect 7136 4380 7200 4384
rect 7136 4324 7140 4380
rect 7140 4324 7196 4380
rect 7196 4324 7200 4380
rect 7136 4320 7200 4324
rect 8896 4380 8960 4384
rect 8896 4324 8900 4380
rect 8900 4324 8956 4380
rect 8956 4324 8960 4380
rect 8896 4320 8960 4324
rect 8976 4380 9040 4384
rect 8976 4324 8980 4380
rect 8980 4324 9036 4380
rect 9036 4324 9040 4380
rect 8976 4320 9040 4324
rect 9056 4380 9120 4384
rect 9056 4324 9060 4380
rect 9060 4324 9116 4380
rect 9116 4324 9120 4380
rect 9056 4320 9120 4324
rect 9136 4380 9200 4384
rect 9136 4324 9140 4380
rect 9140 4324 9196 4380
rect 9196 4324 9200 4380
rect 9136 4320 9200 4324
rect 10896 4380 10960 4384
rect 10896 4324 10900 4380
rect 10900 4324 10956 4380
rect 10956 4324 10960 4380
rect 10896 4320 10960 4324
rect 10976 4380 11040 4384
rect 10976 4324 10980 4380
rect 10980 4324 11036 4380
rect 11036 4324 11040 4380
rect 10976 4320 11040 4324
rect 11056 4380 11120 4384
rect 11056 4324 11060 4380
rect 11060 4324 11116 4380
rect 11116 4324 11120 4380
rect 11056 4320 11120 4324
rect 11136 4380 11200 4384
rect 11136 4324 11140 4380
rect 11140 4324 11196 4380
rect 11196 4324 11200 4380
rect 11136 4320 11200 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 6216 3836 6280 3840
rect 6216 3780 6220 3836
rect 6220 3780 6276 3836
rect 6276 3780 6280 3836
rect 6216 3776 6280 3780
rect 6296 3836 6360 3840
rect 6296 3780 6300 3836
rect 6300 3780 6356 3836
rect 6356 3780 6360 3836
rect 6296 3776 6360 3780
rect 6376 3836 6440 3840
rect 6376 3780 6380 3836
rect 6380 3780 6436 3836
rect 6436 3780 6440 3836
rect 6376 3776 6440 3780
rect 6456 3836 6520 3840
rect 6456 3780 6460 3836
rect 6460 3780 6516 3836
rect 6516 3780 6520 3836
rect 6456 3776 6520 3780
rect 8216 3836 8280 3840
rect 8216 3780 8220 3836
rect 8220 3780 8276 3836
rect 8276 3780 8280 3836
rect 8216 3776 8280 3780
rect 8296 3836 8360 3840
rect 8296 3780 8300 3836
rect 8300 3780 8356 3836
rect 8356 3780 8360 3836
rect 8296 3776 8360 3780
rect 8376 3836 8440 3840
rect 8376 3780 8380 3836
rect 8380 3780 8436 3836
rect 8436 3780 8440 3836
rect 8376 3776 8440 3780
rect 8456 3836 8520 3840
rect 8456 3780 8460 3836
rect 8460 3780 8516 3836
rect 8516 3780 8520 3836
rect 8456 3776 8520 3780
rect 10216 3836 10280 3840
rect 10216 3780 10220 3836
rect 10220 3780 10276 3836
rect 10276 3780 10280 3836
rect 10216 3776 10280 3780
rect 10296 3836 10360 3840
rect 10296 3780 10300 3836
rect 10300 3780 10356 3836
rect 10356 3780 10360 3836
rect 10296 3776 10360 3780
rect 10376 3836 10440 3840
rect 10376 3780 10380 3836
rect 10380 3780 10436 3836
rect 10436 3780 10440 3836
rect 10376 3776 10440 3780
rect 10456 3836 10520 3840
rect 10456 3780 10460 3836
rect 10460 3780 10516 3836
rect 10516 3780 10520 3836
rect 10456 3776 10520 3780
rect 4896 3292 4960 3296
rect 4896 3236 4900 3292
rect 4900 3236 4956 3292
rect 4956 3236 4960 3292
rect 4896 3232 4960 3236
rect 4976 3292 5040 3296
rect 4976 3236 4980 3292
rect 4980 3236 5036 3292
rect 5036 3236 5040 3292
rect 4976 3232 5040 3236
rect 5056 3292 5120 3296
rect 5056 3236 5060 3292
rect 5060 3236 5116 3292
rect 5116 3236 5120 3292
rect 5056 3232 5120 3236
rect 5136 3292 5200 3296
rect 5136 3236 5140 3292
rect 5140 3236 5196 3292
rect 5196 3236 5200 3292
rect 5136 3232 5200 3236
rect 6896 3292 6960 3296
rect 6896 3236 6900 3292
rect 6900 3236 6956 3292
rect 6956 3236 6960 3292
rect 6896 3232 6960 3236
rect 6976 3292 7040 3296
rect 6976 3236 6980 3292
rect 6980 3236 7036 3292
rect 7036 3236 7040 3292
rect 6976 3232 7040 3236
rect 7056 3292 7120 3296
rect 7056 3236 7060 3292
rect 7060 3236 7116 3292
rect 7116 3236 7120 3292
rect 7056 3232 7120 3236
rect 7136 3292 7200 3296
rect 7136 3236 7140 3292
rect 7140 3236 7196 3292
rect 7196 3236 7200 3292
rect 7136 3232 7200 3236
rect 8896 3292 8960 3296
rect 8896 3236 8900 3292
rect 8900 3236 8956 3292
rect 8956 3236 8960 3292
rect 8896 3232 8960 3236
rect 8976 3292 9040 3296
rect 8976 3236 8980 3292
rect 8980 3236 9036 3292
rect 9036 3236 9040 3292
rect 8976 3232 9040 3236
rect 9056 3292 9120 3296
rect 9056 3236 9060 3292
rect 9060 3236 9116 3292
rect 9116 3236 9120 3292
rect 9056 3232 9120 3236
rect 9136 3292 9200 3296
rect 9136 3236 9140 3292
rect 9140 3236 9196 3292
rect 9196 3236 9200 3292
rect 9136 3232 9200 3236
rect 10896 3292 10960 3296
rect 10896 3236 10900 3292
rect 10900 3236 10956 3292
rect 10956 3236 10960 3292
rect 10896 3232 10960 3236
rect 10976 3292 11040 3296
rect 10976 3236 10980 3292
rect 10980 3236 11036 3292
rect 11036 3236 11040 3292
rect 10976 3232 11040 3236
rect 11056 3292 11120 3296
rect 11056 3236 11060 3292
rect 11060 3236 11116 3292
rect 11116 3236 11120 3292
rect 11056 3232 11120 3236
rect 11136 3292 11200 3296
rect 11136 3236 11140 3292
rect 11140 3236 11196 3292
rect 11196 3236 11200 3292
rect 11136 3232 11200 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 6216 2748 6280 2752
rect 6216 2692 6220 2748
rect 6220 2692 6276 2748
rect 6276 2692 6280 2748
rect 6216 2688 6280 2692
rect 6296 2748 6360 2752
rect 6296 2692 6300 2748
rect 6300 2692 6356 2748
rect 6356 2692 6360 2748
rect 6296 2688 6360 2692
rect 6376 2748 6440 2752
rect 6376 2692 6380 2748
rect 6380 2692 6436 2748
rect 6436 2692 6440 2748
rect 6376 2688 6440 2692
rect 6456 2748 6520 2752
rect 6456 2692 6460 2748
rect 6460 2692 6516 2748
rect 6516 2692 6520 2748
rect 6456 2688 6520 2692
rect 8216 2748 8280 2752
rect 8216 2692 8220 2748
rect 8220 2692 8276 2748
rect 8276 2692 8280 2748
rect 8216 2688 8280 2692
rect 8296 2748 8360 2752
rect 8296 2692 8300 2748
rect 8300 2692 8356 2748
rect 8356 2692 8360 2748
rect 8296 2688 8360 2692
rect 8376 2748 8440 2752
rect 8376 2692 8380 2748
rect 8380 2692 8436 2748
rect 8436 2692 8440 2748
rect 8376 2688 8440 2692
rect 8456 2748 8520 2752
rect 8456 2692 8460 2748
rect 8460 2692 8516 2748
rect 8516 2692 8520 2748
rect 8456 2688 8520 2692
rect 10216 2748 10280 2752
rect 10216 2692 10220 2748
rect 10220 2692 10276 2748
rect 10276 2692 10280 2748
rect 10216 2688 10280 2692
rect 10296 2748 10360 2752
rect 10296 2692 10300 2748
rect 10300 2692 10356 2748
rect 10356 2692 10360 2748
rect 10296 2688 10360 2692
rect 10376 2748 10440 2752
rect 10376 2692 10380 2748
rect 10380 2692 10436 2748
rect 10436 2692 10440 2748
rect 10376 2688 10440 2692
rect 10456 2748 10520 2752
rect 10456 2692 10460 2748
rect 10460 2692 10516 2748
rect 10516 2692 10520 2748
rect 10456 2688 10520 2692
rect 4896 2204 4960 2208
rect 4896 2148 4900 2204
rect 4900 2148 4956 2204
rect 4956 2148 4960 2204
rect 4896 2144 4960 2148
rect 4976 2204 5040 2208
rect 4976 2148 4980 2204
rect 4980 2148 5036 2204
rect 5036 2148 5040 2204
rect 4976 2144 5040 2148
rect 5056 2204 5120 2208
rect 5056 2148 5060 2204
rect 5060 2148 5116 2204
rect 5116 2148 5120 2204
rect 5056 2144 5120 2148
rect 5136 2204 5200 2208
rect 5136 2148 5140 2204
rect 5140 2148 5196 2204
rect 5196 2148 5200 2204
rect 5136 2144 5200 2148
rect 6896 2204 6960 2208
rect 6896 2148 6900 2204
rect 6900 2148 6956 2204
rect 6956 2148 6960 2204
rect 6896 2144 6960 2148
rect 6976 2204 7040 2208
rect 6976 2148 6980 2204
rect 6980 2148 7036 2204
rect 7036 2148 7040 2204
rect 6976 2144 7040 2148
rect 7056 2204 7120 2208
rect 7056 2148 7060 2204
rect 7060 2148 7116 2204
rect 7116 2148 7120 2204
rect 7056 2144 7120 2148
rect 7136 2204 7200 2208
rect 7136 2148 7140 2204
rect 7140 2148 7196 2204
rect 7196 2148 7200 2204
rect 7136 2144 7200 2148
rect 8896 2204 8960 2208
rect 8896 2148 8900 2204
rect 8900 2148 8956 2204
rect 8956 2148 8960 2204
rect 8896 2144 8960 2148
rect 8976 2204 9040 2208
rect 8976 2148 8980 2204
rect 8980 2148 9036 2204
rect 9036 2148 9040 2204
rect 8976 2144 9040 2148
rect 9056 2204 9120 2208
rect 9056 2148 9060 2204
rect 9060 2148 9116 2204
rect 9116 2148 9120 2204
rect 9056 2144 9120 2148
rect 9136 2204 9200 2208
rect 9136 2148 9140 2204
rect 9140 2148 9196 2204
rect 9196 2148 9200 2204
rect 9136 2144 9200 2148
rect 10896 2204 10960 2208
rect 10896 2148 10900 2204
rect 10900 2148 10956 2204
rect 10956 2148 10960 2204
rect 10896 2144 10960 2148
rect 10976 2204 11040 2208
rect 10976 2148 10980 2204
rect 10980 2148 11036 2204
rect 11036 2148 11040 2204
rect 10976 2144 11040 2148
rect 11056 2204 11120 2208
rect 11056 2148 11060 2204
rect 11060 2148 11116 2204
rect 11116 2148 11120 2204
rect 11056 2144 11120 2148
rect 11136 2204 11200 2208
rect 11136 2148 11140 2204
rect 11140 2148 11196 2204
rect 11196 2148 11200 2204
rect 11136 2144 11200 2148
<< metal4 >>
rect 4198 12544 4538 12560
rect 4198 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4538 12544
rect 4198 11624 4538 12480
rect 4198 11456 4250 11624
rect 4486 11456 4538 11624
rect 4198 11392 4216 11456
rect 4520 11392 4538 11456
rect 4198 11388 4250 11392
rect 4486 11388 4538 11392
rect 4198 10368 4538 11388
rect 4198 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4538 10368
rect 4198 9624 4538 10304
rect 4198 9388 4250 9624
rect 4486 9388 4538 9624
rect 4198 9280 4538 9388
rect 4198 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4538 9280
rect 4198 8192 4538 9216
rect 4198 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4538 8192
rect 4198 7624 4538 8128
rect 4198 7388 4250 7624
rect 4486 7388 4538 7624
rect 4198 7104 4538 7388
rect 4198 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4538 7104
rect 4198 6016 4538 7040
rect 4198 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4538 6016
rect 4198 5624 4538 5952
rect 4198 5388 4250 5624
rect 4486 5388 4538 5624
rect 4198 4928 4538 5388
rect 4198 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4538 4928
rect 4198 3840 4538 4864
rect 4198 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4538 3840
rect 4198 2752 4538 3776
rect 4198 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4538 2752
rect 4198 2128 4538 2688
rect 4878 12304 5218 12560
rect 4878 12068 4930 12304
rect 5166 12068 5218 12304
rect 4878 12000 5218 12068
rect 4878 11936 4896 12000
rect 4960 11936 4976 12000
rect 5040 11936 5056 12000
rect 5120 11936 5136 12000
rect 5200 11936 5218 12000
rect 4878 10912 5218 11936
rect 4878 10848 4896 10912
rect 4960 10848 4976 10912
rect 5040 10848 5056 10912
rect 5120 10848 5136 10912
rect 5200 10848 5218 10912
rect 4878 10304 5218 10848
rect 4878 10068 4930 10304
rect 5166 10068 5218 10304
rect 4878 9824 5218 10068
rect 4878 9760 4896 9824
rect 4960 9760 4976 9824
rect 5040 9760 5056 9824
rect 5120 9760 5136 9824
rect 5200 9760 5218 9824
rect 4878 8736 5218 9760
rect 4878 8672 4896 8736
rect 4960 8672 4976 8736
rect 5040 8672 5056 8736
rect 5120 8672 5136 8736
rect 5200 8672 5218 8736
rect 4878 8304 5218 8672
rect 4878 8068 4930 8304
rect 5166 8068 5218 8304
rect 4878 7648 5218 8068
rect 4878 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5136 7648
rect 5200 7584 5218 7648
rect 4878 6560 5218 7584
rect 4878 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5136 6560
rect 5200 6496 5218 6560
rect 4878 6304 5218 6496
rect 4878 6068 4930 6304
rect 5166 6068 5218 6304
rect 4878 5472 5218 6068
rect 4878 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5136 5472
rect 5200 5408 5218 5472
rect 4878 4384 5218 5408
rect 4878 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5136 4384
rect 5200 4320 5218 4384
rect 4878 3296 5218 4320
rect 4878 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5136 3296
rect 5200 3232 5218 3296
rect 4878 2208 5218 3232
rect 4878 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5136 2208
rect 5200 2144 5218 2208
rect 4878 2128 5218 2144
rect 6198 12544 6538 12560
rect 6198 12480 6216 12544
rect 6280 12480 6296 12544
rect 6360 12480 6376 12544
rect 6440 12480 6456 12544
rect 6520 12480 6538 12544
rect 6198 11624 6538 12480
rect 6198 11456 6250 11624
rect 6486 11456 6538 11624
rect 6198 11392 6216 11456
rect 6520 11392 6538 11456
rect 6198 11388 6250 11392
rect 6486 11388 6538 11392
rect 6198 10368 6538 11388
rect 6198 10304 6216 10368
rect 6280 10304 6296 10368
rect 6360 10304 6376 10368
rect 6440 10304 6456 10368
rect 6520 10304 6538 10368
rect 6198 9624 6538 10304
rect 6198 9388 6250 9624
rect 6486 9388 6538 9624
rect 6198 9280 6538 9388
rect 6198 9216 6216 9280
rect 6280 9216 6296 9280
rect 6360 9216 6376 9280
rect 6440 9216 6456 9280
rect 6520 9216 6538 9280
rect 6198 8192 6538 9216
rect 6198 8128 6216 8192
rect 6280 8128 6296 8192
rect 6360 8128 6376 8192
rect 6440 8128 6456 8192
rect 6520 8128 6538 8192
rect 6198 7624 6538 8128
rect 6198 7388 6250 7624
rect 6486 7388 6538 7624
rect 6198 7104 6538 7388
rect 6198 7040 6216 7104
rect 6280 7040 6296 7104
rect 6360 7040 6376 7104
rect 6440 7040 6456 7104
rect 6520 7040 6538 7104
rect 6198 6016 6538 7040
rect 6198 5952 6216 6016
rect 6280 5952 6296 6016
rect 6360 5952 6376 6016
rect 6440 5952 6456 6016
rect 6520 5952 6538 6016
rect 6198 5624 6538 5952
rect 6198 5388 6250 5624
rect 6486 5388 6538 5624
rect 6198 4928 6538 5388
rect 6198 4864 6216 4928
rect 6280 4864 6296 4928
rect 6360 4864 6376 4928
rect 6440 4864 6456 4928
rect 6520 4864 6538 4928
rect 6198 3840 6538 4864
rect 6198 3776 6216 3840
rect 6280 3776 6296 3840
rect 6360 3776 6376 3840
rect 6440 3776 6456 3840
rect 6520 3776 6538 3840
rect 6198 2752 6538 3776
rect 6198 2688 6216 2752
rect 6280 2688 6296 2752
rect 6360 2688 6376 2752
rect 6440 2688 6456 2752
rect 6520 2688 6538 2752
rect 6198 2128 6538 2688
rect 6878 12304 7218 12560
rect 6878 12068 6930 12304
rect 7166 12068 7218 12304
rect 6878 12000 7218 12068
rect 6878 11936 6896 12000
rect 6960 11936 6976 12000
rect 7040 11936 7056 12000
rect 7120 11936 7136 12000
rect 7200 11936 7218 12000
rect 6878 10912 7218 11936
rect 6878 10848 6896 10912
rect 6960 10848 6976 10912
rect 7040 10848 7056 10912
rect 7120 10848 7136 10912
rect 7200 10848 7218 10912
rect 6878 10304 7218 10848
rect 6878 10068 6930 10304
rect 7166 10068 7218 10304
rect 6878 9824 7218 10068
rect 6878 9760 6896 9824
rect 6960 9760 6976 9824
rect 7040 9760 7056 9824
rect 7120 9760 7136 9824
rect 7200 9760 7218 9824
rect 6878 8736 7218 9760
rect 6878 8672 6896 8736
rect 6960 8672 6976 8736
rect 7040 8672 7056 8736
rect 7120 8672 7136 8736
rect 7200 8672 7218 8736
rect 6878 8304 7218 8672
rect 6878 8068 6930 8304
rect 7166 8068 7218 8304
rect 6878 7648 7218 8068
rect 6878 7584 6896 7648
rect 6960 7584 6976 7648
rect 7040 7584 7056 7648
rect 7120 7584 7136 7648
rect 7200 7584 7218 7648
rect 6878 6560 7218 7584
rect 6878 6496 6896 6560
rect 6960 6496 6976 6560
rect 7040 6496 7056 6560
rect 7120 6496 7136 6560
rect 7200 6496 7218 6560
rect 6878 6304 7218 6496
rect 6878 6068 6930 6304
rect 7166 6068 7218 6304
rect 6878 5472 7218 6068
rect 6878 5408 6896 5472
rect 6960 5408 6976 5472
rect 7040 5408 7056 5472
rect 7120 5408 7136 5472
rect 7200 5408 7218 5472
rect 6878 4384 7218 5408
rect 6878 4320 6896 4384
rect 6960 4320 6976 4384
rect 7040 4320 7056 4384
rect 7120 4320 7136 4384
rect 7200 4320 7218 4384
rect 6878 3296 7218 4320
rect 6878 3232 6896 3296
rect 6960 3232 6976 3296
rect 7040 3232 7056 3296
rect 7120 3232 7136 3296
rect 7200 3232 7218 3296
rect 6878 2208 7218 3232
rect 6878 2144 6896 2208
rect 6960 2144 6976 2208
rect 7040 2144 7056 2208
rect 7120 2144 7136 2208
rect 7200 2144 7218 2208
rect 6878 2128 7218 2144
rect 8198 12544 8538 12560
rect 8198 12480 8216 12544
rect 8280 12480 8296 12544
rect 8360 12480 8376 12544
rect 8440 12480 8456 12544
rect 8520 12480 8538 12544
rect 8198 11624 8538 12480
rect 8198 11456 8250 11624
rect 8486 11456 8538 11624
rect 8198 11392 8216 11456
rect 8520 11392 8538 11456
rect 8198 11388 8250 11392
rect 8486 11388 8538 11392
rect 8198 10368 8538 11388
rect 8198 10304 8216 10368
rect 8280 10304 8296 10368
rect 8360 10304 8376 10368
rect 8440 10304 8456 10368
rect 8520 10304 8538 10368
rect 8198 9624 8538 10304
rect 8198 9388 8250 9624
rect 8486 9388 8538 9624
rect 8198 9280 8538 9388
rect 8198 9216 8216 9280
rect 8280 9216 8296 9280
rect 8360 9216 8376 9280
rect 8440 9216 8456 9280
rect 8520 9216 8538 9280
rect 8198 8192 8538 9216
rect 8198 8128 8216 8192
rect 8280 8128 8296 8192
rect 8360 8128 8376 8192
rect 8440 8128 8456 8192
rect 8520 8128 8538 8192
rect 8198 7624 8538 8128
rect 8198 7388 8250 7624
rect 8486 7388 8538 7624
rect 8198 7104 8538 7388
rect 8198 7040 8216 7104
rect 8280 7040 8296 7104
rect 8360 7040 8376 7104
rect 8440 7040 8456 7104
rect 8520 7040 8538 7104
rect 8198 6016 8538 7040
rect 8198 5952 8216 6016
rect 8280 5952 8296 6016
rect 8360 5952 8376 6016
rect 8440 5952 8456 6016
rect 8520 5952 8538 6016
rect 8198 5624 8538 5952
rect 8198 5388 8250 5624
rect 8486 5388 8538 5624
rect 8198 4928 8538 5388
rect 8198 4864 8216 4928
rect 8280 4864 8296 4928
rect 8360 4864 8376 4928
rect 8440 4864 8456 4928
rect 8520 4864 8538 4928
rect 8198 3840 8538 4864
rect 8198 3776 8216 3840
rect 8280 3776 8296 3840
rect 8360 3776 8376 3840
rect 8440 3776 8456 3840
rect 8520 3776 8538 3840
rect 8198 2752 8538 3776
rect 8198 2688 8216 2752
rect 8280 2688 8296 2752
rect 8360 2688 8376 2752
rect 8440 2688 8456 2752
rect 8520 2688 8538 2752
rect 8198 2128 8538 2688
rect 8878 12304 9218 12560
rect 8878 12068 8930 12304
rect 9166 12068 9218 12304
rect 8878 12000 9218 12068
rect 8878 11936 8896 12000
rect 8960 11936 8976 12000
rect 9040 11936 9056 12000
rect 9120 11936 9136 12000
rect 9200 11936 9218 12000
rect 8878 10912 9218 11936
rect 8878 10848 8896 10912
rect 8960 10848 8976 10912
rect 9040 10848 9056 10912
rect 9120 10848 9136 10912
rect 9200 10848 9218 10912
rect 8878 10304 9218 10848
rect 8878 10068 8930 10304
rect 9166 10068 9218 10304
rect 8878 9824 9218 10068
rect 8878 9760 8896 9824
rect 8960 9760 8976 9824
rect 9040 9760 9056 9824
rect 9120 9760 9136 9824
rect 9200 9760 9218 9824
rect 8878 8736 9218 9760
rect 8878 8672 8896 8736
rect 8960 8672 8976 8736
rect 9040 8672 9056 8736
rect 9120 8672 9136 8736
rect 9200 8672 9218 8736
rect 8878 8304 9218 8672
rect 8878 8068 8930 8304
rect 9166 8068 9218 8304
rect 8878 7648 9218 8068
rect 8878 7584 8896 7648
rect 8960 7584 8976 7648
rect 9040 7584 9056 7648
rect 9120 7584 9136 7648
rect 9200 7584 9218 7648
rect 8878 6560 9218 7584
rect 8878 6496 8896 6560
rect 8960 6496 8976 6560
rect 9040 6496 9056 6560
rect 9120 6496 9136 6560
rect 9200 6496 9218 6560
rect 8878 6304 9218 6496
rect 8878 6068 8930 6304
rect 9166 6068 9218 6304
rect 8878 5472 9218 6068
rect 8878 5408 8896 5472
rect 8960 5408 8976 5472
rect 9040 5408 9056 5472
rect 9120 5408 9136 5472
rect 9200 5408 9218 5472
rect 8878 4384 9218 5408
rect 8878 4320 8896 4384
rect 8960 4320 8976 4384
rect 9040 4320 9056 4384
rect 9120 4320 9136 4384
rect 9200 4320 9218 4384
rect 8878 3296 9218 4320
rect 8878 3232 8896 3296
rect 8960 3232 8976 3296
rect 9040 3232 9056 3296
rect 9120 3232 9136 3296
rect 9200 3232 9218 3296
rect 8878 2208 9218 3232
rect 8878 2144 8896 2208
rect 8960 2144 8976 2208
rect 9040 2144 9056 2208
rect 9120 2144 9136 2208
rect 9200 2144 9218 2208
rect 8878 2128 9218 2144
rect 10198 12544 10538 12560
rect 10198 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10538 12544
rect 10198 11624 10538 12480
rect 10198 11456 10250 11624
rect 10486 11456 10538 11624
rect 10198 11392 10216 11456
rect 10520 11392 10538 11456
rect 10198 11388 10250 11392
rect 10486 11388 10538 11392
rect 10198 10368 10538 11388
rect 10198 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10538 10368
rect 10198 9624 10538 10304
rect 10198 9388 10250 9624
rect 10486 9388 10538 9624
rect 10198 9280 10538 9388
rect 10198 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10538 9280
rect 10198 8192 10538 9216
rect 10198 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10538 8192
rect 10198 7624 10538 8128
rect 10198 7388 10250 7624
rect 10486 7388 10538 7624
rect 10198 7104 10538 7388
rect 10198 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10538 7104
rect 10198 6016 10538 7040
rect 10198 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10538 6016
rect 10198 5624 10538 5952
rect 10198 5388 10250 5624
rect 10486 5388 10538 5624
rect 10198 4928 10538 5388
rect 10198 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10538 4928
rect 10198 3840 10538 4864
rect 10198 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10538 3840
rect 10198 2752 10538 3776
rect 10198 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10538 2752
rect 10198 2128 10538 2688
rect 10878 12304 11218 12560
rect 10878 12068 10930 12304
rect 11166 12068 11218 12304
rect 10878 12000 11218 12068
rect 10878 11936 10896 12000
rect 10960 11936 10976 12000
rect 11040 11936 11056 12000
rect 11120 11936 11136 12000
rect 11200 11936 11218 12000
rect 10878 10912 11218 11936
rect 10878 10848 10896 10912
rect 10960 10848 10976 10912
rect 11040 10848 11056 10912
rect 11120 10848 11136 10912
rect 11200 10848 11218 10912
rect 10878 10304 11218 10848
rect 10878 10068 10930 10304
rect 11166 10068 11218 10304
rect 10878 9824 11218 10068
rect 10878 9760 10896 9824
rect 10960 9760 10976 9824
rect 11040 9760 11056 9824
rect 11120 9760 11136 9824
rect 11200 9760 11218 9824
rect 10878 8736 11218 9760
rect 10878 8672 10896 8736
rect 10960 8672 10976 8736
rect 11040 8672 11056 8736
rect 11120 8672 11136 8736
rect 11200 8672 11218 8736
rect 10878 8304 11218 8672
rect 10878 8068 10930 8304
rect 11166 8068 11218 8304
rect 10878 7648 11218 8068
rect 10878 7584 10896 7648
rect 10960 7584 10976 7648
rect 11040 7584 11056 7648
rect 11120 7584 11136 7648
rect 11200 7584 11218 7648
rect 10878 6560 11218 7584
rect 10878 6496 10896 6560
rect 10960 6496 10976 6560
rect 11040 6496 11056 6560
rect 11120 6496 11136 6560
rect 11200 6496 11218 6560
rect 10878 6304 11218 6496
rect 10878 6068 10930 6304
rect 11166 6068 11218 6304
rect 10878 5472 11218 6068
rect 10878 5408 10896 5472
rect 10960 5408 10976 5472
rect 11040 5408 11056 5472
rect 11120 5408 11136 5472
rect 11200 5408 11218 5472
rect 10878 4384 11218 5408
rect 10878 4320 10896 4384
rect 10960 4320 10976 4384
rect 11040 4320 11056 4384
rect 11120 4320 11136 4384
rect 11200 4320 11218 4384
rect 10878 3296 11218 4320
rect 10878 3232 10896 3296
rect 10960 3232 10976 3296
rect 11040 3232 11056 3296
rect 11120 3232 11136 3296
rect 11200 3232 11218 3296
rect 10878 2208 11218 3232
rect 10878 2144 10896 2208
rect 10960 2144 10976 2208
rect 11040 2144 11056 2208
rect 11120 2144 11136 2208
rect 11200 2144 11218 2208
rect 10878 2128 11218 2144
<< via4 >>
rect 4250 11456 4486 11624
rect 4250 11392 4280 11456
rect 4280 11392 4296 11456
rect 4296 11392 4360 11456
rect 4360 11392 4376 11456
rect 4376 11392 4440 11456
rect 4440 11392 4456 11456
rect 4456 11392 4486 11456
rect 4250 11388 4486 11392
rect 4250 9388 4486 9624
rect 4250 7388 4486 7624
rect 4250 5388 4486 5624
rect 4930 12068 5166 12304
rect 4930 10068 5166 10304
rect 4930 8068 5166 8304
rect 4930 6068 5166 6304
rect 6250 11456 6486 11624
rect 6250 11392 6280 11456
rect 6280 11392 6296 11456
rect 6296 11392 6360 11456
rect 6360 11392 6376 11456
rect 6376 11392 6440 11456
rect 6440 11392 6456 11456
rect 6456 11392 6486 11456
rect 6250 11388 6486 11392
rect 6250 9388 6486 9624
rect 6250 7388 6486 7624
rect 6250 5388 6486 5624
rect 6930 12068 7166 12304
rect 6930 10068 7166 10304
rect 6930 8068 7166 8304
rect 6930 6068 7166 6304
rect 8250 11456 8486 11624
rect 8250 11392 8280 11456
rect 8280 11392 8296 11456
rect 8296 11392 8360 11456
rect 8360 11392 8376 11456
rect 8376 11392 8440 11456
rect 8440 11392 8456 11456
rect 8456 11392 8486 11456
rect 8250 11388 8486 11392
rect 8250 9388 8486 9624
rect 8250 7388 8486 7624
rect 8250 5388 8486 5624
rect 8930 12068 9166 12304
rect 8930 10068 9166 10304
rect 8930 8068 9166 8304
rect 8930 6068 9166 6304
rect 10250 11456 10486 11624
rect 10250 11392 10280 11456
rect 10280 11392 10296 11456
rect 10296 11392 10360 11456
rect 10360 11392 10376 11456
rect 10376 11392 10440 11456
rect 10440 11392 10456 11456
rect 10456 11392 10486 11456
rect 10250 11388 10486 11392
rect 10250 9388 10486 9624
rect 10250 7388 10486 7624
rect 10250 5388 10486 5624
rect 10930 12068 11166 12304
rect 10930 10068 11166 10304
rect 10930 8068 11166 8304
rect 10930 6068 11166 6304
<< metal5 >>
rect 1056 12304 11916 12356
rect 1056 12068 4930 12304
rect 5166 12068 6930 12304
rect 7166 12068 8930 12304
rect 9166 12068 10930 12304
rect 11166 12068 11916 12304
rect 1056 12016 11916 12068
rect 1056 11624 11916 11676
rect 1056 11388 4250 11624
rect 4486 11388 6250 11624
rect 6486 11388 8250 11624
rect 8486 11388 10250 11624
rect 10486 11388 11916 11624
rect 1056 11336 11916 11388
rect 1056 10304 11916 10356
rect 1056 10068 4930 10304
rect 5166 10068 6930 10304
rect 7166 10068 8930 10304
rect 9166 10068 10930 10304
rect 11166 10068 11916 10304
rect 1056 10016 11916 10068
rect 1056 9624 11916 9676
rect 1056 9388 4250 9624
rect 4486 9388 6250 9624
rect 6486 9388 8250 9624
rect 8486 9388 10250 9624
rect 10486 9388 11916 9624
rect 1056 9336 11916 9388
rect 1056 8304 11916 8356
rect 1056 8068 4930 8304
rect 5166 8068 6930 8304
rect 7166 8068 8930 8304
rect 9166 8068 10930 8304
rect 11166 8068 11916 8304
rect 1056 8016 11916 8068
rect 1056 7624 11916 7676
rect 1056 7388 4250 7624
rect 4486 7388 6250 7624
rect 6486 7388 8250 7624
rect 8486 7388 10250 7624
rect 10486 7388 11916 7624
rect 1056 7336 11916 7388
rect 1056 6304 11916 6356
rect 1056 6068 4930 6304
rect 5166 6068 6930 6304
rect 7166 6068 8930 6304
rect 9166 6068 10930 6304
rect 11166 6068 11916 6304
rect 1056 6016 11916 6068
rect 1056 5624 11916 5676
rect 1056 5388 4250 5624
rect 4486 5388 6250 5624
rect 6486 5388 8250 5624
rect 8486 5388 10250 5624
rect 10486 5388 11916 5624
rect 1056 5336 11916 5388
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK
timestamp 1
transform -1 0 8556 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CLK
timestamp 1
transform 1 0 7544 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CLK
timestamp 1
transform -1 0 7820 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 1
transform -1 0 8832 0 1 7616
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 1
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_27
timestamp 1
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_82
timestamp 1
transform 1 0 8648 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_90
timestamp 1
transform 1 0 9384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_41
timestamp 1
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_85
timestamp 1
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_91
timestamp 1
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_113
timestamp 1
transform 1 0 11500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_27
timestamp 1
transform 1 0 3588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_33
timestamp 1
transform 1 0 4140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_57
timestamp 1
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_65
timestamp 1
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_87
timestamp 1
transform 1 0 9108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_3
timestamp 1
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_50
timestamp 1
transform 1 0 5704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_58
timestamp 1
transform 1 0 6440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_109
timestamp 1
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_113
timestamp 1
transform 1 0 11500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_47
timestamp 1
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_69
timestamp 1
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_37
timestamp 1
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_60
timestamp 1
transform 1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_85
timestamp 1
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_91
timestamp 1
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_113
timestamp 1
transform 1 0 11500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_3
timestamp 1
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_30
timestamp 1
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_34
timestamp 1
transform 1 0 4232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_57
timestamp 1
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_63
timestamp 1
transform 1 0 6900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_85
timestamp 1
transform 1 0 8924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_50
timestamp 1
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_54
timestamp 1
transform 1 0 6072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_76
timestamp 1
transform 1 0 8096 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1636968456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_39
timestamp 1
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_43
timestamp 1
transform 1 0 5060 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_107
timestamp 1
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 1
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 1
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_106
timestamp 1
transform 1 0 10856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_24
timestamp 1
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49
timestamp 1
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_90
timestamp 1636968456
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_102
timestamp 1
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_24
timestamp 1
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_50
timestamp 1
transform 1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_58
timestamp 1
transform 1 0 6440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_109
timestamp 1
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_113
timestamp 1
transform 1 0 11500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_27
timestamp 1
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_35
timestamp 1
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_46
timestamp 1
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_65
timestamp 1
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_78
timestamp 1636968456
transform 1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_29
timestamp 1
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_35
timestamp 1
transform 1 0 4324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_44
timestamp 1
transform 1 0 5152 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_52
timestamp 1
transform 1 0 5888 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_73
timestamp 1
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_89
timestamp 1
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_111
timestamp 1
transform 1 0 11316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_64
timestamp 1
transform 1 0 6992 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_72
timestamp 1
transform 1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_96
timestamp 1636968456
transform 1 0 9936 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 1
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1636968456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_41
timestamp 1
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_106
timestamp 1
transform 1 0 10856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_11
timestamp 1
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_79
timestamp 1636968456
transform 1 0 8372 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_91
timestamp 1636968456
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_103
timestamp 1
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1636968456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_29
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_51
timestamp 1
transform 1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_55
timestamp 1
transform 1 0 6164 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_57
timestamp 1636968456
transform 1 0 6348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_69
timestamp 1636968456
transform 1 0 7452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 1
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1636968456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1636968456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_109
timestamp 1
transform 1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_113
timestamp 1
transform 1 0 11500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_19
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_20
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_21
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_22
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_23
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_24
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 11868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_25
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_26
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 11868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_27
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_28
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_29
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_30
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 11868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_31
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_32
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 11868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_33
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 11868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_34
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_35
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_36
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 11868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_37
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_40
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_41
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_44
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_46
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_47
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_48
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_49
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_50
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_51
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_52
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_53
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_54
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_55
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_56
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_57
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_58
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_59
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_60
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_61
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_62
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_63
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_64
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_65
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_66
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_67
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_68
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_69
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_70
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_71
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_72
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_73
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_74
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_75
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_76
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_77
timestamp 1
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_78
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_79
timestamp 1
transform 1 0 11408 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  x1_x1
timestamp 1
transform 1 0 9660 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1_x2
timestamp 1
transform 1 0 9476 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1_x3
timestamp 1
transform 1 0 9568 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1_x4
timestamp 1
transform 1 0 9384 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_8  x1_x5
timestamp 1
transform -1 0 6256 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  x1_x6
timestamp 1
transform 1 0 9476 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1_x7
timestamp 1
transform 1 0 9568 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1_x8
timestamp 1
transform 1 0 9476 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1_x9
timestamp 1
transform -1 0 8648 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1_x10
timestamp 1
transform -1 0 6900 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x1_x11
timestamp 1
transform 1 0 6900 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x1
timestamp 1
transform 1 0 4968 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x2
timestamp 1
transform 1 0 6440 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x3
timestamp 1
transform 1 0 6900 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  x2_x4
timestamp 1
transform -1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  x2_x5
timestamp 1
transform 1 0 8004 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x7
timestamp 1
transform -1 0 6256 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x11
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x12
timestamp 1
transform 1 0 2116 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x13
timestamp 1
transform -1 0 5980 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x14
timestamp 1
transform -1 0 3680 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x15
timestamp 1
transform 1 0 1748 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x16
timestamp 1
transform 1 0 2392 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x2_x21
timestamp 1
transform 1 0 3864 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  x2_x22
timestamp 1
transform -1 0 5152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x2_x23
timestamp 1
transform 1 0 4416 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_8  x2_x24
timestamp 1
transform -1 0 5336 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  x2_x25
timestamp 1
transform 1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  x3_x1
timestamp 1
transform -1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_0
timestamp 1
transform 1 0 6992 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_1
timestamp 1
transform 1 0 6900 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_2
timestamp 1
transform 1 0 6716 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_3
timestamp 1
transform 1 0 7176 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_4
timestamp 1
transform -1 0 6256 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_5
timestamp 1
transform 1 0 4232 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_6
timestamp 1
transform -1 0 5704 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_7
timestamp 1
transform -1 0 3680 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_8
timestamp 1
transform -1 0 3496 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x1_9
timestamp 1
transform -1 0 6624 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_8  x3_x2
timestamp 1
transform -1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_0
timestamp 1
transform -1 0 5704 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_1
timestamp 1
transform -1 0 8096 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_2
timestamp 1
transform -1 0 6256 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_3
timestamp 1
transform -1 0 8648 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_4
timestamp 1
transform -1 0 5888 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_5
timestamp 1
transform -1 0 5612 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_6
timestamp 1
transform -1 0 5704 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_7
timestamp 1
transform -1 0 3680 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_8
timestamp 1
transform -1 0 3864 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x3_x2_9
timestamp 1
transform -1 0 5428 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_0
timestamp 1
transform 1 0 9384 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_1
timestamp 1
transform 1 0 9384 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_2
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_3
timestamp 1
transform 1 0 9016 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_4
timestamp 1
transform 1 0 8924 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_5
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_6
timestamp 1
transform 1 0 5888 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_7
timestamp 1
transform -1 0 3312 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_8
timestamp 1
transform -1 0 3312 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  x4_x1_9
timestamp 1
transform -1 0 3680 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  x4_x1
timestamp 1
transform 1 0 8280 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x4_x2
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 498 592
<< labels >>
flabel metal3 s 12188 8 12988 128 0 FreeSans 480 0 0 0 CF[0]
port 0 nsew signal output
flabel metal3 s 12188 688 12988 808 0 FreeSans 480 0 0 0 CF[1]
port 1 nsew signal output
flabel metal3 s 12188 1368 12988 1488 0 FreeSans 480 0 0 0 CF[2]
port 2 nsew signal output
flabel metal3 s 12188 2048 12988 2168 0 FreeSans 480 0 0 0 CF[3]
port 3 nsew signal output
flabel metal3 s 12188 2728 12988 2848 0 FreeSans 480 0 0 0 CF[4]
port 4 nsew signal output
flabel metal3 s 12188 3408 12988 3528 0 FreeSans 480 0 0 0 CF[5]
port 5 nsew signal output
flabel metal3 s 12188 4088 12988 4208 0 FreeSans 480 0 0 0 CF[6]
port 6 nsew signal output
flabel metal3 s 12188 4768 12988 4888 0 FreeSans 480 0 0 0 CF[7]
port 7 nsew signal output
flabel metal3 s 12188 5448 12988 5568 0 FreeSans 480 0 0 0 CF[8]
port 8 nsew signal output
flabel metal3 s 12188 6128 12988 6248 0 FreeSans 480 0 0 0 CF[9]
port 9 nsew signal output
flabel metal3 s 12188 6808 12988 6928 0 FreeSans 480 0 0 0 CKO
port 10 nsew signal output
flabel metal3 s 12188 7488 12988 7608 0 FreeSans 480 0 0 0 CLK
port 11 nsew signal input
flabel metal3 s 12188 8168 12988 8288 0 FreeSans 480 0 0 0 CLKS
port 12 nsew signal output
flabel metal3 s 12188 8848 12988 8968 0 FreeSans 480 0 0 0 CLKSB
port 13 nsew signal output
flabel metal3 s 12188 9528 12988 9648 0 FreeSans 480 0 0 0 COMP_N
port 14 nsew signal input
flabel metal3 s 12188 10208 12988 10328 0 FreeSans 480 0 0 0 COMP_P
port 15 nsew signal input
flabel metal3 s 12188 10888 12988 11008 0 FreeSans 480 0 0 0 DOUT[0]
port 16 nsew signal output
flabel metal3 s 12188 11568 12988 11688 0 FreeSans 480 0 0 0 DOUT[1]
port 17 nsew signal output
flabel metal3 s 12188 12248 12988 12368 0 FreeSans 480 0 0 0 DOUT[2]
port 18 nsew signal output
flabel metal3 s 12188 12928 12988 13048 0 FreeSans 480 0 0 0 DOUT[3]
port 19 nsew signal output
flabel metal3 s 12188 13608 12988 13728 0 FreeSans 480 0 0 0 DOUT[4]
port 20 nsew signal output
flabel metal3 s 12188 14288 12988 14408 0 FreeSans 480 0 0 0 DOUT[5]
port 21 nsew signal output
flabel metal3 s 12188 14968 12988 15088 0 FreeSans 480 0 0 0 DOUT[6]
port 22 nsew signal output
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 DOUT[7]
port 23 nsew signal output
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 DOUT[8]
port 24 nsew signal output
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 DOUT[9]
port 25 nsew signal output
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 EN
port 26 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 SWN[0]
port 27 nsew signal output
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 SWN[1]
port 28 nsew signal output
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 SWN[2]
port 29 nsew signal output
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 SWN[3]
port 30 nsew signal output
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 SWN[4]
port 31 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 SWN[5]
port 32 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 SWN[6]
port 33 nsew signal output
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 SWN[7]
port 34 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 SWN[8]
port 35 nsew signal output
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 SWN[9]
port 36 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 SWP[0]
port 37 nsew signal output
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 SWP[1]
port 38 nsew signal output
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 SWP[2]
port 39 nsew signal output
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 SWP[3]
port 40 nsew signal output
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 SWP[4]
port 41 nsew signal output
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 SWP[5]
port 42 nsew signal output
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 SWP[6]
port 43 nsew signal output
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 SWP[7]
port 44 nsew signal output
flabel metal3 s 0 8 800 128 0 FreeSans 480 0 0 0 SWP[8]
port 45 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 SWP[9]
port 46 nsew signal output
flabel metal4 s 4198 2128 4538 12560 0 FreeSans 1920 90 0 0 VDDD
port 47 nsew power input
flabel metal4 s 6198 2128 6538 12560 0 FreeSans 1920 90 0 0 VDDD
port 47 nsew power input
flabel metal4 s 8198 2128 8538 12560 0 FreeSans 1920 90 0 0 VDDD
port 47 nsew power input
flabel metal4 s 10198 2128 10538 12560 0 FreeSans 1920 90 0 0 VDDD
port 47 nsew power input
flabel metal5 s 1056 5336 11916 5676 0 FreeSans 2560 0 0 0 VDDD
port 47 nsew power input
flabel metal5 s 1056 7336 11916 7676 0 FreeSans 2560 0 0 0 VDDD
port 47 nsew power input
flabel metal5 s 1056 9336 11916 9676 0 FreeSans 2560 0 0 0 VDDD
port 47 nsew power input
flabel metal5 s 1056 11336 11916 11676 0 FreeSans 2560 0 0 0 VDDD
port 47 nsew power input
flabel metal4 s 4878 2128 5218 12560 0 FreeSans 1920 90 0 0 VSSD
port 48 nsew ground input
flabel metal4 s 6878 2128 7218 12560 0 FreeSans 1920 90 0 0 VSSD
port 48 nsew ground input
flabel metal4 s 8878 2128 9218 12560 0 FreeSans 1920 90 0 0 VSSD
port 48 nsew ground input
flabel metal4 s 10878 2128 11218 12560 0 FreeSans 1920 90 0 0 VSSD
port 48 nsew ground input
flabel metal5 s 1056 6016 11916 6356 0 FreeSans 2560 0 0 0 VSSD
port 48 nsew ground input
flabel metal5 s 1056 8016 11916 8356 0 FreeSans 2560 0 0 0 VSSD
port 48 nsew ground input
flabel metal5 s 1056 10016 11916 10356 0 FreeSans 2560 0 0 0 VSSD
port 48 nsew ground input
flabel metal5 s 1056 12016 11916 12356 0 FreeSans 2560 0 0 0 VSSD
port 48 nsew ground input
rlabel via1 6486 12512 6486 12512 0 VDDD
rlabel metal1 6486 11968 6486 11968 0 VSSD
rlabel metal3 10726 68 10726 68 0 CF[0]
rlabel metal3 9760 748 9760 748 0 CF[1]
rlabel metal3 9484 1428 9484 1428 0 CF[2]
rlabel metal3 11830 2108 11830 2108 0 CF[3]
rlabel metal1 6210 3060 6210 3060 0 CF[4]
rlabel metal1 4922 4046 4922 4046 0 CF[5]
rlabel metal1 11224 4998 11224 4998 0 CF[6]
rlabel metal2 11362 5185 11362 5185 0 CF[7]
rlabel metal1 11362 6086 11362 6086 0 CF[8]
rlabel metal2 11454 6409 11454 6409 0 CF[9]
rlabel metal2 8970 7021 8970 7021 0 CKO
rlabel metal1 8510 7480 8510 7480 0 CLK
rlabel metal2 2622 4896 2622 4896 0 CLKS
rlabel via1 11017 8806 11017 8806 0 CLKSB
rlabel via2 8234 9571 8234 9571 0 COMP_N
rlabel metal2 9338 9299 9338 9299 0 COMP_P
rlabel metal1 11270 9486 11270 9486 0 DOUT[0]
rlabel metal1 11224 10234 11224 10234 0 DOUT[1]
rlabel metal1 10764 9146 10764 9146 0 DOUT[2]
rlabel metal3 11416 12988 11416 12988 0 DOUT[3]
rlabel metal3 11508 13668 11508 13668 0 DOUT[4]
rlabel metal3 10174 14348 10174 14348 0 DOUT[5]
rlabel metal3 10726 15028 10726 15028 0 DOUT[6]
rlabel metal1 2070 8398 2070 8398 0 DOUT[7]
rlabel metal3 1786 14348 1786 14348 0 DOUT[8]
rlabel metal3 1924 13668 1924 13668 0 DOUT[9]
rlabel metal3 1740 12988 1740 12988 0 EN
rlabel metal1 7222 7310 7222 7310 0 FINAL
rlabel metal2 3910 10727 3910 10727 0 SWN[0]
rlabel metal1 6210 6834 6210 6834 0 SWN[1]
rlabel metal1 4554 6426 4554 6426 0 SWN[2]
rlabel metal3 1717 10268 1717 10268 0 SWN[3]
rlabel metal2 4094 8823 4094 8823 0 SWN[4]
rlabel metal2 1334 8755 1334 8755 0 SWN[5]
rlabel metal2 3910 7531 3910 7531 0 SWN[6]
rlabel metal2 2806 6715 2806 6715 0 SWN[7]
rlabel metal1 1656 6426 1656 6426 0 SWN[8]
rlabel metal2 3634 5763 3634 5763 0 SWN[9]
rlabel metal3 1717 5508 1717 5508 0 SWP[0]
rlabel metal3 1717 4828 1717 4828 0 SWP[1]
rlabel metal2 8510 4301 8510 4301 0 SWP[2]
rlabel metal2 8970 3689 8970 3689 0 SWP[3]
rlabel metal3 1717 2788 1717 2788 0 SWP[4]
rlabel metal3 5083 2380 5083 2380 0 SWP[5]
rlabel metal3 2292 1428 2292 1428 0 SWP[6]
rlabel metal1 2300 4454 2300 4454 0 SWP[7]
rlabel metal3 1832 68 1832 68 0 SWP[8]
rlabel metal2 6256 748 6256 748 0 SWP[9]
rlabel metal1 7268 7514 7268 7514 0 clknet_0_CLK
rlabel metal1 6900 3570 6900 3570 0 clknet_1_0__leaf_CLK
rlabel metal1 2438 11798 2438 11798 0 clknet_1_1__leaf_CLK
rlabel metal2 5934 11934 5934 11934 0 x2/TRIG1
rlabel metal1 2438 10744 2438 10744 0 x2/TRIG2
rlabel metal1 5096 11322 5096 11322 0 x2/net1
rlabel metal2 4186 12002 4186 12002 0 x2/net10
rlabel metal1 7107 10642 7107 10642 0 x2/net11
rlabel metal1 4876 10030 4876 10030 0 x2/net12
rlabel metal2 4738 9724 4738 9724 0 x2/net13
rlabel metal2 6762 11492 6762 11492 0 x2/net2
rlabel metal2 7222 11288 7222 11288 0 x2/net3
rlabel metal1 8464 10710 8464 10710 0 x2/net4
rlabel metal2 9798 10982 9798 10982 0 x2/net5
rlabel metal1 4784 10574 4784 10574 0 x2/net6
rlabel metal1 3450 10098 3450 10098 0 x2/net7
rlabel metal1 1978 10234 1978 10234 0 x2/net8
rlabel metal2 2714 11492 2714 11492 0 x2/net9
rlabel metal2 7866 9248 7866 9248 0 x3/COMP_BUF_N
rlabel metal1 7360 6358 7360 6358 0 x3/COMP_BUF_P
<< properties >>
string FIXED_BBOX 0 0 12988 15132
<< end >>