* PEX produced on Min 03 Nov 2024 04:00:20  CST using ./iic-pex.sh with m=1 and s=1
* NGSPICE file created from auto_sampling.ext - technology: sky130A

X0 VDDD a_869_n2275# a_856_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_8421_n3089# a_7340_n3089# a_8074_n2847# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2 VDDD a_10528_n3115# x21.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_10007_n2007# a_9789_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4 VDDD a_8421_n3089# a_8596_n3115# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VDDD x23.Y CLKS VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 x3.Q a_6665_n2275# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X7 VDDD a_8074_n2847# a_7964_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X8 a_4210_n2847# a_3992_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X9 a_7762_n2249# x3.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 a_2979_n3089# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X11 a_4732_n3115# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X12 a_6143_n2007# a_5925_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X13 a_8118_n3089# a_8074_n2847# a_7952_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X14 a_10528_n3115# a_10353_n3089# a_10707_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X15 a_10050_n3089# a_10006_n2847# a_9884_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X16 a_8075_n2007# a_7857_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X17 a_1710_n3089# a_1544_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_10007_n2007# a_9789_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X19 VSSD a_10528_n3115# x21.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VSSD x23.Y CLKS VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_868_n3115# a_693_n3089# a_1047_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X22 a_1710_n3089# a_1544_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 a_856_n1883# a_n221_n2249# a_694_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 VSSD a_868_n3115# a_802_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_2735_n2249# a_1545_n2249# a_2626_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X26 VDDD a_2800_n3115# a_2787_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X27 VSSD x23.Y CLKS VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 VSSD CKC a_n387_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 a_803_n2249# a_n387_n2249# a_694_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X30 VDDD CKC a_n387_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X31 a_9896_n2723# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X32 a_7762_n2249# x3.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X33 VSSD RST a_10051_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X34 a_6664_n3115# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X35 a_2626_n2249# a_1545_n2249# a_2279_n2007# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X36 VSSD CKC a_1544_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X37 CLKS x23.Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 a_3642_n3089# a_3476_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X39 VDDD CKC a_1544_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X40 a_694_n2249# a_n221_n2249# a_347_n2007# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X41 a_2787_n2723# a_1710_n3089# a_2625_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X42 a_3642_n3089# a_3476_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X43 a_34_n2249# x21.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X44 a_693_n3089# a_n388_n3089# a_346_n2847# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X45 CLKS x23.Y VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X46 a_2980_n2249# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X47 a_8596_n3115# a_8421_n3089# a_8775_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X48 VSSD CKC a_n388_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X49 x23.Y x22.Y VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X50 VSSD a_2801_n2275# a_2735_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X51 VDDD a_868_n3115# x12.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X52 VDDD a_346_n2847# a_236_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X53 VDDD CKC a_n388_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X54 a_9788_n3089# a_9272_n3089# a_9693_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X55 VDDD a_8597_n2275# a_8584_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X56 a_6598_n3089# a_5408_n3089# a_6489_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X57 x16.Q a_8596_n3115# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X58 a_4558_n2249# a_3477_n2249# a_4211_n2007# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X59 a_9693_n3089# x16.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X60 VSSD CKC a_3476_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X61 VDDD x23.Y CLKS VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X62 a_2061_n2249# a_1545_n2249# a_1966_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X63 VDDD a_4733_n2275# x2.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X64 VDDD CKC a_3476_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X65 a_4720_n1883# a_3643_n2249# a_4558_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X66 a_2278_n2847# a_2060_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X67 VDDD x12.Q x22.Y VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X68 a_2156_n3089# a_1710_n3089# a_2060_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X69 a_5575_n2249# a_5409_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X70 VSSD a_868_n3115# x12.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X71 VDDD a_4211_n2007# a_4101_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X72 a_2169_n1883# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X73 a_5575_n2249# a_5409_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X74 x21.Q a_10528_n3115# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X75 VSSD RST a_8119_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X76 a_6489_n3089# a_5574_n3089# a_6142_n2847# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X77 VDDD x22.Y x23.Y VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 x16.Q a_8596_n3115# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X79 x12.Q a_868_n3115# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X80 a_224_n3089# a_n222_n3089# a_128_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X81 a_10707_n3089# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X82 a_1965_n3089# x12.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X83 VSSD a_10528_n3115# a_10462_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X84 a_7964_n2723# a_7340_n3089# a_7856_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X85 a_1047_n3089# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X86 a_236_n2723# a_n388_n3089# a_128_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X87 a_3897_n3089# x13.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X88 a_3992_n3089# a_3642_n3089# a_3897_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X89 a_10463_n2249# a_9273_n2249# a_10354_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X90 x21.Q a_10528_n3115# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X91 a_6652_n1883# a_5575_n2249# a_6490_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X92 VSSD a_6664_n3115# a_6598_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X93 x22.Y x12.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X94 a_4210_n2847# a_3992_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X95 x12.Q a_868_n3115# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X96 a_4101_n1883# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X97 a_4089_n2249# a_3643_n2249# a_3993_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X98 VDDD a_4557_n3089# a_4732_n3115# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X99 VSSD a_2801_n2275# x1.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X100 a_9884_n3089# a_9438_n3089# a_9788_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X101 a_3898_n2249# x1.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X102 a_10354_n2249# a_9439_n2249# a_10007_n2007# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X103 a_391_n2249# a_347_n2007# a_225_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X104 CLKSB CLKS VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X105 VDDD a_10354_n2249# a_10529_n2275# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X106 a_10515_n2723# a_9438_n3089# a_10353_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X107 a_5924_n3089# a_5574_n3089# a_5829_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X108 VDDD a_694_n2249# a_869_n2275# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X109 VDDD a_10006_n2847# a_9896_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X110 a_8775_n3089# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X111 a_6490_n2249# a_5575_n2249# a_6143_n2007# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X112 a_6489_n3089# a_5408_n3089# a_6142_n2847# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X113 VSSD a_8597_n2275# a_8531_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X114 VDDD a_6664_n3115# x15.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X115 x1.Q a_2801_n2275# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X116 VSSD RST a_391_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X117 a_9789_n2249# a_9439_n2249# a_9694_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X118 a_8531_n2249# a_7341_n2249# a_8422_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X119 VDDD a_6142_n2847# a_6032_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X120 VDDD x23.Y CLKS VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X121 VSSD RST a_4254_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X122 a_5830_n2249# x2.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X123 a_4100_n2723# a_3476_n3089# a_3992_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X124 a_10529_n2275# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X125 VDDD x23.Y CLKS VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X126 a_346_n2847# a_128_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X127 a_6186_n3089# a_6142_n2847# a_6020_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X128 a_6143_n2007# a_5925_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X129 a_869_n2275# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X130 VSSD a_6664_n3115# x15.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X131 VSSD CKC a_7340_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X132 VDDD a_8596_n3115# x16.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X133 VDDD CKC a_7340_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X134 VDDD a_8422_n2249# a_8597_n2275# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X135 a_4732_n3115# a_4557_n3089# a_4911_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X136 a_8583_n2723# a_7506_n3089# a_8421_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X137 CLKS x23.Y VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X138 a_6032_n2723# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X139 VDDD a_4733_n2275# a_4720_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X140 VSSD RST a_6186_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X141 a_5924_n3089# a_5408_n3089# a_5829_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X142 a_5830_n2249# x2.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X143 VDDD a_2279_n2007# a_2169_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X144 a_6032_n2723# a_5408_n3089# a_5924_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X145 x14.Q a_4732_n3115# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X146 VSSD a_8596_n3115# x16.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X147 a_10529_n2275# a_10354_n2249# a_10708_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X148 a_8119_n2249# a_8075_n2007# a_7953_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X149 a_34_n2249# x21.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X150 x12.D x11.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X151 a_10051_n2249# a_10007_n2007# a_9885_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X152 a_1711_n2249# a_1545_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X153 VSSD a_10529_n2275# x11.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X154 a_869_n2275# a_694_n2249# a_1048_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X155 VSSD CKC a_9272_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X156 a_1711_n2249# a_1545_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X157 a_8597_n2275# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X158 VSSD a_869_n2275# a_803_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X159 a_2625_n3089# a_1710_n3089# a_2278_n2847# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X160 VDDD a_2625_n3089# a_2800_n3115# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X161 a_6664_n3115# a_6489_n3089# a_6843_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X162 VDDD CKC a_9272_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X163 a_8074_n2847# a_7856_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X164 x14.Q a_4732_n3115# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X165 a_7965_n1883# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X166 a_7856_n3089# a_7340_n3089# a_7761_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X167 VDDD a_6665_n2275# a_6652_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X168 a_4666_n3089# a_3476_n3089# a_4557_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X169 a_2169_n1883# a_1545_n2249# a_2061_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X170 x15.Q a_6664_n3115# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X171 a_7761_n3089# x15.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X172 VDDD a_2801_n2275# x1.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X173 VSSD CKC a_1545_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X174 a_128_n3089# a_n388_n3089# a_33_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X175 a_3643_n2249# a_3477_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X176 VDDD CKC a_1545_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X177 a_694_n2249# a_n387_n2249# a_347_n2007# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X178 a_9693_n3089# x16.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X179 a_3643_n2249# a_3477_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X180 a_8074_n2847# a_7856_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X181 a_10006_n2847# a_9788_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X182 a_4557_n3089# a_3642_n3089# a_4210_n2847# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X183 VDDD a_10528_n3115# a_10515_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X184 a_855_n2723# a_n222_n3089# a_693_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X185 x15.Q a_6664_n3115# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X186 a_6020_n3089# a_5574_n3089# a_5924_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X187 a_8597_n2275# a_8422_n2249# a_8776_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X188 a_9789_n2249# a_9273_n2249# a_9694_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X189 a_1965_n3089# x12.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X190 a_6599_n2249# a_5409_n2249# a_6490_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X191 x1.Q a_2801_n2275# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X192 a_4911_n3089# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X193 VSSD a_4732_n3115# a_4666_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X194 a_9897_n1883# a_9273_n2249# a_9789_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X195 VSSD CKC a_3477_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X196 CLKSB CLKS VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X197 a_2625_n3089# a_1544_n3089# a_2278_n2847# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X198 VDDD CKC a_3477_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X199 a_2279_n2007# a_2061_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X200 a_2157_n2249# a_1711_n2249# a_2061_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X201 a_2800_n3115# a_2625_n3089# a_2979_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X202 VSSD a_869_n2275# x1.D VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X203 a_7952_n3089# a_7506_n3089# a_7856_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X204 a_346_n2847# a_128_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X205 a_237_n1883# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X206 a_10708_n2249# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X207 x5.Q a_8597_n2275# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X208 a_225_n2249# a_n221_n2249# a_129_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X209 a_7506_n3089# a_7340_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X210 VSSD a_10529_n2275# a_10463_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X211 VDDD a_6490_n2249# a_6665_n2275# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X212 a_1048_n2249# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X213 a_2322_n3089# a_2278_n2847# a_2156_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X214 a_7506_n3089# a_7340_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X215 VDDD a_8596_n3115# a_8583_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X216 a_2279_n2007# a_2061_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X217 a_6843_n3089# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X218 a_3898_n2249# x1.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X219 x11.Q a_10529_n2275# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X220 a_4557_n3089# a_3476_n3089# a_4210_n2847# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X221 a_2800_n3115# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X222 VSSD a_6665_n2275# a_6599_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X223 VDDD a_4732_n3115# x14.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X224 a_4211_n2007# a_3993_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X225 x1.D a_869_n2275# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X226 a_129_n2249# a_n221_n2249# a_34_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X227 a_7857_n2249# a_7507_n2249# a_7762_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X228 VDDD a_4210_n2847# a_4100_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X229 a_2168_n2723# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X230 VSSD RST a_2322_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X231 a_8422_n2249# a_7341_n2249# a_8075_n2007# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X232 a_9885_n2249# a_9439_n2249# a_9789_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X233 x12.D x11.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X234 a_10354_n2249# a_9273_n2249# a_10007_n2007# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X235 a_9438_n3089# a_9272_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X236 VDDD a_10529_n2275# x11.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X237 a_4254_n3089# a_4210_n2847# a_4088_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X238 a_9438_n3089# a_9272_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X239 a_4211_n2007# a_3993_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X240 VSSD a_4732_n3115# x14.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X241 VDDD a_8075_n2007# a_7965_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X242 a_8776_n2249# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X243 VSSD CKC a_5408_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X244 a_4733_n2275# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X245 VDDD CKC a_5408_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X246 a_2060_n3089# a_1710_n3089# a_1965_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X247 a_6651_n2723# a_5574_n3089# a_6489_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X248 a_4100_n2723# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X249 VDDD a_2801_n2275# a_2788_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X250 a_3992_n3089# a_3476_n3089# a_3897_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X251 a_8421_n3089# a_7506_n3089# a_8074_n2847# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X252 VSSD RST a_4255_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X253 VDDD a_868_n3115# a_855_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X254 a_10006_n2847# a_9788_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X255 a_9897_n1883# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X256 a_6187_n2249# a_6143_n2007# a_6021_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X257 CLKS x23.Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X258 VSSD a_6665_n2275# x3.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X259 VDDD a_10353_n3089# a_10528_n3115# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X260 a_6665_n2275# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X261 VDDD a_693_n3089# a_868_n3115# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X262 VSSD CKC a_7341_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X263 a_6142_n2847# a_5924_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X264 a_2788_n1883# a_1711_n2249# a_2626_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X265 VDDD CKC a_7341_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X266 a_4733_n2275# a_4558_n2249# a_4912_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X267 a_6033_n1883# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X268 CLKS x23.Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X269 a_2734_n3089# a_1544_n3089# a_2625_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X270 a_9788_n3089# a_9438_n3089# a_9693_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X271 VSSD RST a_6187_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X272 a_5925_n2249# a_5409_n2249# a_5830_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X273 a_5829_n3089# x14.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X274 VDDD a_347_n2007# a_237_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X275 VDDD a_869_n2275# x1.D VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X276 a_802_n3089# a_n388_n3089# a_693_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X277 a_10528_n3115# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X278 VSSD a_8597_n2275# x5.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X279 x23.Y x22.Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X280 a_7761_n3089# x15.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X281 VSSD x22.Y x23.Y VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X282 x5.Q a_8597_n2275# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X283 a_6142_n2847# a_5924_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X284 a_868_n3115# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X285 a_9694_n2249# x5.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X286 VSSD RST a_10050_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X287 VSSD CKC a_9273_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X288 a_2626_n2249# a_1711_n2249# a_2279_n2007# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X289 VDDD CKC a_9273_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X290 a_6665_n2275# a_6490_n2249# a_6844_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X291 a_8075_n2007# a_7857_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X292 x2.Q a_4733_n2275# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X293 VSSD x23.Y CLKS VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X294 a_693_n3089# a_n222_n3089# a_346_n2847# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X295 x11.Q a_10529_n2275# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X296 a_33_n3089# x12.D VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X297 a_7857_n2249# a_7341_n2249# a_7762_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X298 a_4667_n2249# a_3477_n2249# a_4558_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X299 VDDD a_4732_n3115# a_4719_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X300 x1.D a_869_n2275# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X301 VDDD a_2278_n2847# a_2168_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X302 a_1966_n2249# x1.D VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X303 a_237_n1883# a_n387_n2249# a_129_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X304 VSSD a_2800_n3115# a_2734_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X305 a_7965_n1883# a_7341_n2249# a_7857_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X306 a_129_n2249# a_n387_n2249# a_34_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X307 VDDD a_10529_n2275# a_10516_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X308 a_3993_n2249# a_3643_n2249# a_3898_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X309 a_33_n3089# x12.D VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X310 a_9694_n2249# x5.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X311 a_4558_n2249# a_3643_n2249# a_4211_n2007# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X312 a_2060_n3089# a_1544_n3089# a_1965_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X313 a_8596_n3115# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X314 a_6021_n2249# a_5575_n2249# a_5925_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X315 x3.Q a_6665_n2275# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X316 a_5574_n3089# a_5408_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X317 VDDD a_4558_n2249# a_4733_n2275# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X318 a_7964_n2723# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X319 a_4719_n2723# a_3642_n3089# a_4557_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X320 VSSD RST a_8118_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X321 a_5574_n3089# a_5408_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X322 VDDD a_6664_n3115# a_6651_n2723# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X323 a_1966_n2249# x1.D VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X324 a_2168_n2723# a_1544_n3089# a_2060_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X325 a_4912_n2249# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X326 VSSD a_4733_n2275# a_4667_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X327 VDDD a_2800_n3115# x13.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X328 a_10516_n1883# a_9439_n2249# a_10354_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X329 a_5925_n2249# a_5575_n2249# a_5830_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X330 VDDD a_10007_n2007# a_9897_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X331 a_2801_n2275# a_2626_n2249# a_2980_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X332 a_10462_n3089# a_9272_n3089# a_10353_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X333 CLKS x23.Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X334 a_6490_n2249# a_5409_n2249# a_6143_n2007# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X335 a_347_n2007# a_129_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X336 a_7953_n2249# a_7507_n2249# a_7857_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X337 a_n221_n2249# a_n387_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X338 VDDD a_6665_n2275# x3.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X339 a_n221_n2249# a_n387_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X340 x23.Y x22.Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X341 a_4088_n3089# a_3642_n3089# a_3992_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X342 a_7507_n2249# a_7341_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X343 VSSD a_2800_n3115# x13.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X344 VDDD a_6143_n2007# a_6033_n1883# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X345 a_2323_n2249# a_2279_n2007# a_2157_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X346 a_7507_n2249# a_7341_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X347 a_4101_n1883# a_3477_n2249# a_3993_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X348 a_10353_n3089# a_9438_n3089# a_10006_n2847# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X349 a_6844_n2249# RST VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X350 a_390_n3089# a_346_n2847# a_224_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X351 VSSD x23.Y CLKS VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X352 x13.Q a_2800_n3115# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X353 a_2801_n2275# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X354 a_347_n2007# a_129_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X355 a_3897_n3089# x13.Q VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X356 a_9896_n2723# a_9272_n3089# a_9788_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X357 VSSD x12.Q x22.Y VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X358 a_10353_n3089# a_9272_n3089# a_10006_n2847# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X359 CLKS x23.Y VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X360 a_5829_n3089# x14.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X361 a_n222_n3089# a_n388_n3089# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X362 VSSD x22.Y x23.Y VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X363 VSSD RST a_2323_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X364 a_n222_n3089# a_n388_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X365 VDDD a_8597_n2275# x5.Q VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X366 a_8584_n1883# a_7507_n2249# a_8422_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X367 VSSD a_8596_n3115# a_8530_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X368 a_236_n2723# RST VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X369 x13.Q a_2800_n3115# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X370 VSSD RST a_390_n3089# VSSD sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X371 a_9439_n2249# a_9273_n2249# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X372 a_8530_n3089# a_7340_n3089# a_8421_n3089# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X373 a_4255_n2249# a_4211_n2007# a_4089_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X374 a_9439_n2249# a_9273_n2249# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X375 a_6033_n1883# a_5409_n2249# a_5925_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X376 VDDD a_6489_n3089# a_6664_n3115# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X377 VSSD a_4733_n2275# x2.Q VSSD sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X378 CLKS x23.Y VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X379 x2.Q a_4733_n2275# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X380 a_2278_n2847# a_2060_n3089# VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X381 x22.Y x12.Q VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X382 a_2061_n2249# a_1711_n2249# a_1966_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X383 VSSD CKC a_5409_n2249# VSSD sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X384 VDDD CKC a_5409_n2249# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X385 x23.Y x22.Y VDDD VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X386 a_7856_n3089# a_7506_n3089# a_7761_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X387 a_128_n3089# a_n222_n3089# a_33_n3089# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X388 a_3993_n2249# a_3477_n2249# a_3898_n2249# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X389 VDDD x22.Y x23.Y VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X390 VDDD a_2626_n2249# a_2801_n2275# VDDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X391 a_8422_n2249# a_7507_n2249# a_8075_n2007# VSSD sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
C0 CLKSB VSSD 0.47924f
C1 CLKS VSSD 1.91823f
C2 RST VSSD 23.174099f
C3 CKC VSSD 13.7939f
C4 VDDD VSSD 61.2144f
C5 x23.Y VSSD 2.31504f $ **FLOATING
C6 x22.Y VSSD 1.2196f $ **FLOATING
C7 a_9896_n2723# VSSD 0.167731f $ **FLOATING
C8 a_9693_n3089# VSSD 0.258962f $ **FLOATING
C9 a_10353_n3089# VSSD 0.736061f $ **FLOATING
C10 a_10528_n3115# VSSD 1.13276f $ **FLOATING
C11 a_9788_n3089# VSSD 0.714373f $ **FLOATING
C12 a_10006_n2847# VSSD 0.652907f $ **FLOATING
C13 a_9438_n3089# VSSD 1.56815f $ **FLOATING
C14 a_9272_n3089# VSSD 1.91526f $ **FLOATING
C15 x16.Q VSSD 1.00558f $ **FLOATING
C16 a_7964_n2723# VSSD 0.167731f $ **FLOATING
C17 a_7761_n3089# VSSD 0.258962f $ **FLOATING
C18 a_8421_n3089# VSSD 0.736061f $ **FLOATING
C19 a_8596_n3115# VSSD 1.13276f $ **FLOATING
C20 a_7856_n3089# VSSD 0.714373f $ **FLOATING
C21 a_8074_n2847# VSSD 0.652907f $ **FLOATING
C22 a_7506_n3089# VSSD 1.56815f $ **FLOATING
C23 a_7340_n3089# VSSD 1.91526f $ **FLOATING
C24 x15.Q VSSD 1.00558f $ **FLOATING
C25 a_6032_n2723# VSSD 0.167731f $ **FLOATING
C26 a_5829_n3089# VSSD 0.258962f $ **FLOATING
C27 a_6489_n3089# VSSD 0.736061f $ **FLOATING
C28 a_6664_n3115# VSSD 1.13276f $ **FLOATING
C29 a_5924_n3089# VSSD 0.714373f $ **FLOATING
C30 a_6142_n2847# VSSD 0.652907f $ **FLOATING
C31 a_5574_n3089# VSSD 1.56815f $ **FLOATING
C32 a_5408_n3089# VSSD 1.91526f $ **FLOATING
C33 x14.Q VSSD 1.00558f $ **FLOATING
C34 a_4100_n2723# VSSD 0.167731f $ **FLOATING
C35 a_3897_n3089# VSSD 0.258962f $ **FLOATING
C36 a_4557_n3089# VSSD 0.736061f $ **FLOATING
C37 a_4732_n3115# VSSD 1.13276f $ **FLOATING
C38 a_3992_n3089# VSSD 0.714373f $ **FLOATING
C39 a_4210_n2847# VSSD 0.652907f $ **FLOATING
C40 a_3642_n3089# VSSD 1.56815f $ **FLOATING
C41 a_3476_n3089# VSSD 1.91526f $ **FLOATING
C42 x13.Q VSSD 1.00558f $ **FLOATING
C43 a_2168_n2723# VSSD 0.167731f $ **FLOATING
C44 a_1965_n3089# VSSD 0.258962f $ **FLOATING
C45 a_2625_n3089# VSSD 0.736061f $ **FLOATING
C46 a_2800_n3115# VSSD 1.13276f $ **FLOATING
C47 a_2060_n3089# VSSD 0.714373f $ **FLOATING
C48 a_2278_n2847# VSSD 0.652907f $ **FLOATING
C49 a_1710_n3089# VSSD 1.56815f $ **FLOATING
C50 a_1544_n3089# VSSD 1.91526f $ **FLOATING
C51 x12.Q VSSD 2.4147f $ **FLOATING
C52 a_236_n2723# VSSD 0.167731f $ **FLOATING
C53 a_33_n3089# VSSD 0.258962f $ **FLOATING
C54 a_693_n3089# VSSD 0.736061f $ **FLOATING
C55 a_868_n3115# VSSD 1.13276f $ **FLOATING
C56 a_128_n3089# VSSD 0.714373f $ **FLOATING
C57 a_346_n2847# VSSD 0.652907f $ **FLOATING
C58 a_n222_n3089# VSSD 1.56815f $ **FLOATING
C59 a_n388_n3089# VSSD 1.91526f $ **FLOATING
C60 x12.D VSSD 6.27447f $ **FLOATING
C61 a_9897_n1883# VSSD 0.167731f $ **FLOATING
C62 a_9694_n2249# VSSD 0.258962f $ **FLOATING
C63 x11.Q VSSD 0.60369f $ **FLOATING
C64 a_10354_n2249# VSSD 0.736061f $ **FLOATING
C65 a_10529_n2275# VSSD 1.13276f $ **FLOATING
C66 a_9789_n2249# VSSD 0.714373f $ **FLOATING
C67 a_10007_n2007# VSSD 0.652907f $ **FLOATING
C68 a_9439_n2249# VSSD 1.56815f $ **FLOATING
C69 a_9273_n2249# VSSD 1.91526f $ **FLOATING
C70 x5.Q VSSD 1.00558f $ **FLOATING
C71 a_7965_n1883# VSSD 0.167731f $ **FLOATING
C72 a_7762_n2249# VSSD 0.258962f $ **FLOATING
C73 a_8422_n2249# VSSD 0.736061f $ **FLOATING
C74 a_8597_n2275# VSSD 1.13276f $ **FLOATING
C75 a_7857_n2249# VSSD 0.714373f $ **FLOATING
C76 a_8075_n2007# VSSD 0.652907f $ **FLOATING
C77 a_7507_n2249# VSSD 1.56815f $ **FLOATING
C78 a_7341_n2249# VSSD 1.91526f $ **FLOATING
C79 x3.Q VSSD 1.00558f $ **FLOATING
C80 a_6033_n1883# VSSD 0.167731f $ **FLOATING
C81 a_5830_n2249# VSSD 0.258962f $ **FLOATING
C82 a_6490_n2249# VSSD 0.736061f $ **FLOATING
C83 a_6665_n2275# VSSD 1.13276f $ **FLOATING
C84 a_5925_n2249# VSSD 0.714373f $ **FLOATING
C85 a_6143_n2007# VSSD 0.652907f $ **FLOATING
C86 a_5575_n2249# VSSD 1.56815f $ **FLOATING
C87 a_5409_n2249# VSSD 1.91526f $ **FLOATING
C88 x2.Q VSSD 1.00558f $ **FLOATING
C89 a_4101_n1883# VSSD 0.167731f $ **FLOATING
C90 a_3898_n2249# VSSD 0.258962f $ **FLOATING
C91 a_4558_n2249# VSSD 0.736061f $ **FLOATING
C92 a_4733_n2275# VSSD 1.13276f $ **FLOATING
C93 a_3993_n2249# VSSD 0.714373f $ **FLOATING
C94 a_4211_n2007# VSSD 0.652907f $ **FLOATING
C95 a_3643_n2249# VSSD 1.56815f $ **FLOATING
C96 a_3477_n2249# VSSD 1.91526f $ **FLOATING
C97 x1.Q VSSD 1.00558f $ **FLOATING
C98 a_2169_n1883# VSSD 0.167731f $ **FLOATING
C99 a_1966_n2249# VSSD 0.258962f $ **FLOATING
C100 a_2626_n2249# VSSD 0.736061f $ **FLOATING
C101 a_2801_n2275# VSSD 1.13276f $ **FLOATING
C102 a_2061_n2249# VSSD 0.714373f $ **FLOATING
C103 a_2279_n2007# VSSD 0.652907f $ **FLOATING
C104 a_1711_n2249# VSSD 1.56815f $ **FLOATING
C105 a_1545_n2249# VSSD 1.91526f $ **FLOATING
C106 x1.D VSSD 1.00558f $ **FLOATING
C107 a_237_n1883# VSSD 0.167731f $ **FLOATING
C108 a_34_n2249# VSSD 0.258962f $ **FLOATING
C109 a_694_n2249# VSSD 0.736061f $ **FLOATING
C110 a_869_n2275# VSSD 1.13276f $ **FLOATING
C111 a_129_n2249# VSSD 0.714373f $ **FLOATING
C112 a_347_n2007# VSSD 0.652907f $ **FLOATING
C113 a_n221_n2249# VSSD 1.56815f $ **FLOATING
C114 x21.Q VSSD 6.16888f $ **FLOATING
C115 a_n387_n2249# VSSD 1.91526f $ **FLOATING
