magic
tech sky130A
magscale 1 2
timestamp 1730624594
<< locali >>
rect 321 -2082 355 -2006
rect 321 -2172 355 -2166
rect 707 -2082 741 -2006
rect 707 -2172 741 -2166
rect 813 -2206 847 -2006
rect 813 -2296 847 -2290
rect 1199 -2206 1233 -2006
rect 1199 -2296 1233 -2290
<< viali >>
rect 321 -2166 355 -2082
rect 707 -2166 741 -2082
rect 813 -2290 847 -2206
rect 1199 -2290 1233 -2206
<< metal1 >>
rect 485 6521 505 6573
rect 557 6521 577 6573
rect 415 6431 421 6483
rect 473 6431 479 6483
rect 415 6359 479 6431
rect 415 6307 421 6359
rect 473 6307 479 6359
rect 415 6235 479 6307
rect 415 6183 421 6235
rect 473 6183 479 6235
rect 583 6431 589 6483
rect 641 6431 647 6483
rect 583 6359 647 6431
rect 583 6307 589 6359
rect 641 6307 647 6359
rect 583 6235 647 6307
rect 583 6183 589 6235
rect 641 6183 647 6235
rect 485 6093 505 6145
rect 557 6093 577 6145
rect 485 5985 505 6037
rect 557 5985 577 6037
rect 415 5895 421 5947
rect 473 5895 479 5947
rect 415 5823 479 5895
rect 415 5771 421 5823
rect 473 5771 479 5823
rect 415 5699 479 5771
rect 415 5647 421 5699
rect 473 5647 479 5699
rect 583 5895 589 5947
rect 641 5895 647 5947
rect 583 5823 647 5895
rect 583 5771 589 5823
rect 641 5771 647 5823
rect 583 5699 647 5771
rect 583 5647 589 5699
rect 641 5647 647 5699
rect 485 5557 505 5609
rect 557 5557 577 5609
rect 485 5449 505 5501
rect 557 5449 577 5501
rect 415 5359 421 5411
rect 473 5359 479 5411
rect 415 5287 479 5359
rect 415 5235 421 5287
rect 473 5235 479 5287
rect 415 5163 479 5235
rect 415 5111 421 5163
rect 473 5111 479 5163
rect 583 5359 589 5411
rect 641 5359 647 5411
rect 583 5287 647 5359
rect 583 5235 589 5287
rect 641 5235 647 5287
rect 583 5163 647 5235
rect 583 5111 589 5163
rect 641 5111 647 5163
rect 485 5021 505 5073
rect 557 5021 577 5073
rect 485 4913 505 4965
rect 557 4913 577 4965
rect 415 4823 421 4875
rect 473 4823 479 4875
rect 415 4751 479 4823
rect 415 4699 421 4751
rect 473 4699 479 4751
rect 415 4627 479 4699
rect 415 4575 421 4627
rect 473 4575 479 4627
rect 583 4823 589 4875
rect 641 4823 647 4875
rect 583 4751 647 4823
rect 583 4699 589 4751
rect 641 4699 647 4751
rect 583 4627 647 4699
rect 583 4575 589 4627
rect 641 4575 647 4627
rect 583 4566 647 4575
rect 485 4485 505 4537
rect 557 4485 577 4537
rect 485 4377 505 4429
rect 557 4377 577 4429
rect 415 4287 421 4339
rect 473 4287 479 4339
rect 415 4215 479 4287
rect 415 4163 421 4215
rect 473 4163 479 4215
rect 415 4091 479 4163
rect 415 4039 421 4091
rect 473 4039 479 4091
rect 583 4287 589 4339
rect 641 4287 647 4339
rect 583 4215 647 4287
rect 583 4163 589 4215
rect 641 4163 647 4215
rect 583 4091 647 4163
rect 583 4039 589 4091
rect 641 4039 647 4091
rect 485 3949 505 4001
rect 557 3949 577 4001
rect 485 3841 505 3893
rect 557 3841 577 3893
rect 415 3751 421 3803
rect 473 3751 479 3803
rect 415 3679 479 3751
rect 415 3627 421 3679
rect 473 3627 479 3679
rect 415 3555 479 3627
rect 415 3503 421 3555
rect 473 3503 479 3555
rect 583 3751 589 3803
rect 641 3751 647 3803
rect 583 3679 647 3751
rect 583 3627 589 3679
rect 641 3627 647 3679
rect 583 3555 647 3627
rect 583 3503 589 3555
rect 641 3503 647 3555
rect 485 3413 505 3465
rect 557 3413 577 3465
rect 485 3305 505 3357
rect 557 3305 577 3357
rect 415 3215 421 3267
rect 473 3215 479 3267
rect 415 3143 479 3215
rect 415 3091 421 3143
rect 473 3091 479 3143
rect 415 3019 479 3091
rect 415 2967 421 3019
rect 473 2967 479 3019
rect 583 3215 589 3267
rect 641 3215 647 3267
rect 583 3143 647 3215
rect 583 3091 589 3143
rect 641 3091 647 3143
rect 583 3019 647 3091
rect 977 3033 997 3085
rect 1049 3033 1069 3085
rect 583 2967 589 3019
rect 641 2967 647 3019
rect 907 2956 971 3004
rect 485 2877 505 2929
rect 557 2877 577 2929
rect 907 2904 913 2956
rect 965 2904 971 2956
rect 1075 2956 1139 3004
rect 1075 2904 1081 2956
rect 1133 2904 1139 2956
rect 977 2823 997 2875
rect 1049 2823 1069 2875
rect 485 2769 505 2821
rect 557 2769 577 2821
rect 415 2679 421 2731
rect 473 2679 479 2731
rect 415 2607 479 2679
rect 415 2555 421 2607
rect 473 2555 479 2607
rect 415 2483 479 2555
rect 415 2431 421 2483
rect 473 2431 479 2483
rect 583 2679 589 2731
rect 641 2686 647 2731
rect 977 2715 997 2767
rect 1049 2715 1069 2767
rect 641 2679 971 2686
rect 583 2638 971 2679
rect 583 2607 913 2638
rect 583 2555 589 2607
rect 641 2586 913 2607
rect 965 2586 971 2638
rect 1075 2638 1139 2686
rect 1075 2586 1081 2638
rect 1133 2586 1139 2638
rect 641 2555 647 2586
rect 583 2483 647 2555
rect 977 2505 997 2557
rect 1049 2505 1069 2557
rect 583 2431 589 2483
rect 641 2431 647 2483
rect 583 2422 647 2431
rect 977 2397 997 2449
rect 1049 2397 1069 2449
rect 485 2341 505 2393
rect 557 2341 577 2393
rect 907 2320 971 2368
rect 485 2233 505 2285
rect 557 2233 577 2285
rect 907 2268 913 2320
rect 965 2268 971 2320
rect 1075 2320 1139 2368
rect 1075 2268 1081 2320
rect 1133 2268 1139 2320
rect 415 2143 421 2195
rect 473 2143 479 2195
rect 415 2071 479 2143
rect 415 2019 421 2071
rect 473 2019 479 2071
rect 415 1947 479 2019
rect 415 1895 421 1947
rect 473 1895 479 1947
rect 583 2143 589 2195
rect 641 2143 647 2195
rect 977 2187 997 2239
rect 1049 2187 1069 2239
rect 583 2071 647 2143
rect 977 2079 997 2131
rect 1049 2079 1069 2131
rect 583 2019 589 2071
rect 641 2050 647 2071
rect 641 2019 971 2050
rect 583 2002 971 2019
rect 583 1950 913 2002
rect 965 1950 971 2002
rect 1075 2002 1139 2050
rect 1075 1950 1081 2002
rect 1133 1950 1139 2002
rect 583 1947 647 1950
rect 583 1895 589 1947
rect 641 1895 647 1947
rect 977 1869 997 1921
rect 1049 1869 1069 1921
rect 485 1805 505 1857
rect 557 1805 577 1857
rect 977 1761 997 1813
rect 1049 1761 1069 1813
rect 485 1697 505 1749
rect 557 1697 577 1749
rect 907 1684 971 1732
rect 415 1607 421 1659
rect 473 1607 479 1659
rect 415 1535 479 1607
rect 415 1483 421 1535
rect 473 1483 479 1535
rect 415 1411 479 1483
rect 415 1359 421 1411
rect 473 1359 479 1411
rect 583 1607 589 1659
rect 641 1607 647 1659
rect 907 1632 913 1684
rect 965 1632 971 1684
rect 1075 1684 1139 1732
rect 1075 1632 1081 1684
rect 1133 1632 1139 1684
rect 583 1535 647 1607
rect 977 1551 997 1603
rect 1049 1551 1069 1603
rect 583 1483 589 1535
rect 641 1483 647 1535
rect 583 1411 647 1483
rect 977 1443 997 1495
rect 1049 1443 1069 1495
rect 583 1359 589 1411
rect 641 1359 647 1411
rect 907 1366 971 1414
rect 485 1269 505 1321
rect 557 1269 577 1321
rect 907 1314 913 1366
rect 965 1314 971 1366
rect 1075 1366 1139 1414
rect 1075 1314 1081 1366
rect 1133 1314 1139 1366
rect 977 1233 997 1285
rect 1049 1233 1069 1285
rect 485 1161 505 1213
rect 557 1161 577 1213
rect 977 1125 997 1177
rect 1049 1125 1069 1177
rect 415 1071 421 1123
rect 473 1071 479 1123
rect 415 999 479 1071
rect 415 947 421 999
rect 473 947 479 999
rect 415 875 479 947
rect 415 823 421 875
rect 473 823 479 875
rect 583 1071 589 1123
rect 641 1096 647 1123
rect 641 1071 971 1096
rect 583 1048 971 1071
rect 583 999 913 1048
rect 583 947 589 999
rect 641 996 913 999
rect 965 996 971 1048
rect 1075 1048 1139 1096
rect 1075 996 1081 1048
rect 1133 996 1139 1048
rect 641 947 647 996
rect 583 875 647 947
rect 977 915 997 967
rect 1049 915 1069 967
rect 583 823 589 875
rect 641 823 647 875
rect 977 807 997 859
rect 1049 807 1069 859
rect 485 733 505 785
rect 557 733 577 785
rect 907 730 971 778
rect 907 678 913 730
rect 965 678 971 730
rect 1075 730 1139 778
rect 1075 678 1081 730
rect 1133 678 1139 730
rect 485 625 505 677
rect 557 625 577 677
rect 977 597 997 649
rect 1049 597 1069 649
rect 415 535 421 587
rect 473 535 479 587
rect 415 463 479 535
rect 415 411 421 463
rect 473 411 479 463
rect 415 339 479 411
rect 415 287 421 339
rect 473 287 479 339
rect 583 535 589 587
rect 641 535 647 587
rect 583 463 647 535
rect 977 489 997 541
rect 1049 489 1069 541
rect 583 411 589 463
rect 641 460 647 463
rect 641 412 971 460
rect 641 411 913 412
rect 583 360 913 411
rect 965 360 971 412
rect 1075 412 1139 460
rect 1075 360 1081 412
rect 1133 360 1139 412
rect 583 339 647 360
rect 583 287 589 339
rect 641 287 647 339
rect 583 278 647 287
rect 977 279 997 331
rect 1049 279 1069 331
rect 485 197 505 249
rect 557 197 577 249
rect 977 171 997 223
rect 1049 171 1069 223
rect 485 89 505 141
rect 557 89 577 141
rect 907 94 971 142
rect 415 -1 421 51
rect 473 -1 479 51
rect 415 -73 479 -1
rect 415 -125 421 -73
rect 473 -125 479 -73
rect 415 -197 479 -125
rect 415 -249 421 -197
rect 473 -249 479 -197
rect 583 -1 589 51
rect 641 -1 647 51
rect 907 42 913 94
rect 965 42 971 94
rect 1075 94 1139 142
rect 1075 42 1081 94
rect 1133 42 1139 94
rect 583 -73 647 -1
rect 977 -39 997 13
rect 1049 -39 1069 13
rect 583 -125 589 -73
rect 641 -125 647 -73
rect 583 -197 647 -125
rect 977 -147 997 -95
rect 1049 -147 1069 -95
rect 583 -249 589 -197
rect 641 -249 647 -197
rect 907 -224 971 -176
rect 907 -276 913 -224
rect 965 -276 971 -224
rect 1075 -224 1139 -176
rect 1075 -276 1081 -224
rect 1133 -276 1139 -224
rect 485 -339 505 -287
rect 557 -339 577 -287
rect 977 -357 997 -305
rect 1049 -357 1069 -305
rect 485 -447 505 -395
rect 557 -447 577 -395
rect 977 -465 997 -413
rect 1049 -465 1069 -413
rect 415 -537 421 -485
rect 473 -537 479 -485
rect 415 -609 479 -537
rect 415 -661 421 -609
rect 473 -661 479 -609
rect 415 -733 479 -661
rect 415 -785 421 -733
rect 473 -785 479 -733
rect 583 -537 589 -485
rect 641 -494 647 -485
rect 641 -537 971 -494
rect 583 -542 971 -537
rect 583 -594 913 -542
rect 965 -594 971 -542
rect 1075 -542 1139 -494
rect 1075 -594 1081 -542
rect 1133 -594 1139 -542
rect 583 -609 647 -594
rect 583 -661 589 -609
rect 641 -661 647 -609
rect 583 -733 647 -661
rect 977 -675 997 -623
rect 1049 -675 1069 -623
rect 583 -785 589 -733
rect 641 -785 647 -733
rect 977 -783 997 -731
rect 1049 -783 1069 -731
rect 485 -875 505 -823
rect 557 -875 577 -823
rect 907 -860 971 -812
rect 907 -912 913 -860
rect 965 -912 971 -860
rect 1075 -860 1139 -812
rect 1075 -912 1081 -860
rect 1133 -912 1139 -860
rect 485 -983 505 -931
rect 557 -983 577 -931
rect 977 -993 997 -941
rect 1049 -993 1069 -941
rect 415 -1073 421 -1021
rect 473 -1073 479 -1021
rect 415 -1145 479 -1073
rect 415 -1197 421 -1145
rect 473 -1197 479 -1145
rect 415 -1269 479 -1197
rect 415 -1321 421 -1269
rect 473 -1321 479 -1269
rect 583 -1073 589 -1021
rect 641 -1073 647 -1021
rect 583 -1130 647 -1073
rect 977 -1101 997 -1049
rect 1049 -1101 1069 -1049
rect 583 -1145 971 -1130
rect 583 -1197 589 -1145
rect 641 -1178 971 -1145
rect 641 -1197 913 -1178
rect 583 -1230 913 -1197
rect 965 -1230 971 -1178
rect 1075 -1178 1139 -1130
rect 1075 -1230 1081 -1178
rect 1133 -1230 1139 -1178
rect 583 -1269 647 -1230
rect 583 -1321 589 -1269
rect 641 -1321 647 -1269
rect 977 -1311 997 -1259
rect 1049 -1311 1069 -1259
rect 485 -1411 505 -1359
rect 557 -1411 577 -1359
rect 977 -1419 997 -1367
rect 1049 -1419 1069 -1367
rect 485 -1519 505 -1467
rect 557 -1519 577 -1467
rect 907 -1496 971 -1448
rect 907 -1548 913 -1496
rect 965 -1548 971 -1496
rect 1075 -1496 1139 -1448
rect 1075 -1548 1081 -1496
rect 1133 -1548 1139 -1496
rect 415 -1609 421 -1557
rect 473 -1609 479 -1557
rect 415 -1681 479 -1609
rect 415 -1733 421 -1681
rect 473 -1733 479 -1681
rect 415 -1805 479 -1733
rect 415 -1857 421 -1805
rect 473 -1857 479 -1805
rect 583 -1609 589 -1557
rect 641 -1609 647 -1557
rect 583 -1681 647 -1609
rect 977 -1629 997 -1577
rect 1049 -1629 1069 -1577
rect 583 -1733 589 -1681
rect 641 -1733 647 -1681
rect 583 -1766 647 -1733
rect 977 -1737 997 -1685
rect 1049 -1737 1069 -1685
rect 583 -1805 971 -1766
rect 583 -1857 589 -1805
rect 641 -1814 971 -1805
rect 641 -1857 913 -1814
rect 583 -1866 913 -1857
rect 965 -1866 971 -1814
rect 1075 -1814 1139 -1766
rect 1075 -1866 1081 -1814
rect 1133 -1866 1139 -1814
rect 485 -1947 505 -1895
rect 557 -1947 577 -1895
rect 977 -1947 997 -1895
rect 1049 -1947 1069 -1895
rect 415 -2033 421 -1981
rect 473 -2033 1081 -1981
rect 1133 -2033 1139 -1981
rect 285 -2082 1269 -2076
rect 285 -2166 321 -2082
rect 355 -2166 707 -2082
rect 741 -2166 1269 -2082
rect 285 -2172 1269 -2166
rect 285 -2206 1269 -2200
rect 285 -2290 813 -2206
rect 847 -2290 1199 -2206
rect 1233 -2290 1269 -2206
rect 285 -2296 1269 -2290
rect 285 -2376 421 -2324
rect 473 -2376 1269 -2324
rect 285 -2382 1269 -2376
<< via1 >>
rect 505 6521 557 6573
rect 421 6431 473 6483
rect 421 6307 473 6359
rect 421 6183 473 6235
rect 589 6431 641 6483
rect 589 6307 641 6359
rect 589 6183 641 6235
rect 505 6093 557 6145
rect 505 5985 557 6037
rect 421 5895 473 5947
rect 421 5771 473 5823
rect 421 5647 473 5699
rect 589 5895 641 5947
rect 589 5771 641 5823
rect 589 5647 641 5699
rect 505 5557 557 5609
rect 505 5449 557 5501
rect 421 5359 473 5411
rect 421 5235 473 5287
rect 421 5111 473 5163
rect 589 5359 641 5411
rect 589 5235 641 5287
rect 589 5111 641 5163
rect 505 5021 557 5073
rect 505 4913 557 4965
rect 421 4823 473 4875
rect 421 4699 473 4751
rect 421 4575 473 4627
rect 589 4823 641 4875
rect 589 4699 641 4751
rect 589 4575 641 4627
rect 505 4485 557 4537
rect 505 4377 557 4429
rect 421 4287 473 4339
rect 421 4163 473 4215
rect 421 4039 473 4091
rect 589 4287 641 4339
rect 589 4163 641 4215
rect 589 4039 641 4091
rect 505 3949 557 4001
rect 505 3841 557 3893
rect 421 3751 473 3803
rect 421 3627 473 3679
rect 421 3503 473 3555
rect 589 3751 641 3803
rect 589 3627 641 3679
rect 589 3503 641 3555
rect 505 3413 557 3465
rect 505 3305 557 3357
rect 421 3215 473 3267
rect 421 3091 473 3143
rect 421 2967 473 3019
rect 589 3215 641 3267
rect 589 3091 641 3143
rect 997 3033 1049 3085
rect 589 2967 641 3019
rect 505 2877 557 2929
rect 913 2904 965 2956
rect 1081 2904 1133 2956
rect 997 2823 1049 2875
rect 505 2769 557 2821
rect 421 2679 473 2731
rect 421 2555 473 2607
rect 421 2431 473 2483
rect 589 2679 641 2731
rect 997 2715 1049 2767
rect 589 2555 641 2607
rect 913 2586 965 2638
rect 1081 2586 1133 2638
rect 997 2505 1049 2557
rect 589 2431 641 2483
rect 997 2397 1049 2449
rect 505 2341 557 2393
rect 505 2233 557 2285
rect 913 2268 965 2320
rect 1081 2268 1133 2320
rect 421 2143 473 2195
rect 421 2019 473 2071
rect 421 1895 473 1947
rect 589 2143 641 2195
rect 997 2187 1049 2239
rect 997 2079 1049 2131
rect 589 2019 641 2071
rect 913 1950 965 2002
rect 1081 1950 1133 2002
rect 589 1895 641 1947
rect 997 1869 1049 1921
rect 505 1805 557 1857
rect 997 1761 1049 1813
rect 505 1697 557 1749
rect 421 1607 473 1659
rect 421 1483 473 1535
rect 421 1359 473 1411
rect 589 1607 641 1659
rect 913 1632 965 1684
rect 1081 1632 1133 1684
rect 997 1551 1049 1603
rect 589 1483 641 1535
rect 997 1443 1049 1495
rect 589 1359 641 1411
rect 505 1269 557 1321
rect 913 1314 965 1366
rect 1081 1314 1133 1366
rect 997 1233 1049 1285
rect 505 1161 557 1213
rect 997 1125 1049 1177
rect 421 1071 473 1123
rect 421 947 473 999
rect 421 823 473 875
rect 589 1071 641 1123
rect 589 947 641 999
rect 913 996 965 1048
rect 1081 996 1133 1048
rect 997 915 1049 967
rect 589 823 641 875
rect 997 807 1049 859
rect 505 733 557 785
rect 913 678 965 730
rect 1081 678 1133 730
rect 505 625 557 677
rect 997 597 1049 649
rect 421 535 473 587
rect 421 411 473 463
rect 421 287 473 339
rect 589 535 641 587
rect 997 489 1049 541
rect 589 411 641 463
rect 913 360 965 412
rect 1081 360 1133 412
rect 589 287 641 339
rect 997 279 1049 331
rect 505 197 557 249
rect 997 171 1049 223
rect 505 89 557 141
rect 421 -1 473 51
rect 421 -125 473 -73
rect 421 -249 473 -197
rect 589 -1 641 51
rect 913 42 965 94
rect 1081 42 1133 94
rect 997 -39 1049 13
rect 589 -125 641 -73
rect 997 -147 1049 -95
rect 589 -249 641 -197
rect 913 -276 965 -224
rect 1081 -276 1133 -224
rect 505 -339 557 -287
rect 997 -357 1049 -305
rect 505 -447 557 -395
rect 997 -465 1049 -413
rect 421 -537 473 -485
rect 421 -661 473 -609
rect 421 -785 473 -733
rect 589 -537 641 -485
rect 913 -594 965 -542
rect 1081 -594 1133 -542
rect 589 -661 641 -609
rect 997 -675 1049 -623
rect 589 -785 641 -733
rect 997 -783 1049 -731
rect 505 -875 557 -823
rect 913 -912 965 -860
rect 1081 -912 1133 -860
rect 505 -983 557 -931
rect 997 -993 1049 -941
rect 421 -1073 473 -1021
rect 421 -1197 473 -1145
rect 421 -1321 473 -1269
rect 589 -1073 641 -1021
rect 997 -1101 1049 -1049
rect 589 -1197 641 -1145
rect 913 -1230 965 -1178
rect 1081 -1230 1133 -1178
rect 589 -1321 641 -1269
rect 997 -1311 1049 -1259
rect 505 -1411 557 -1359
rect 997 -1419 1049 -1367
rect 505 -1519 557 -1467
rect 913 -1548 965 -1496
rect 1081 -1548 1133 -1496
rect 421 -1609 473 -1557
rect 421 -1733 473 -1681
rect 421 -1857 473 -1805
rect 589 -1609 641 -1557
rect 997 -1629 1049 -1577
rect 589 -1733 641 -1681
rect 997 -1737 1049 -1685
rect 589 -1857 641 -1805
rect 913 -1866 965 -1814
rect 1081 -1866 1133 -1814
rect 505 -1947 557 -1895
rect 997 -1947 1049 -1895
rect 421 -2033 473 -1981
rect 1081 -2033 1133 -1981
rect 421 -2376 473 -2324
<< metal2 >>
rect 503 6573 559 6579
rect 503 6521 505 6573
rect 557 6521 559 6573
rect 419 6483 475 6489
rect 419 6431 421 6483
rect 473 6431 475 6483
rect 419 6359 475 6431
rect 419 6307 421 6359
rect 473 6307 475 6359
rect 419 6235 475 6307
rect 419 6183 421 6235
rect 473 6183 475 6235
rect 419 5947 475 6183
rect 419 5895 421 5947
rect 473 5895 475 5947
rect 419 5823 475 5895
rect 419 5771 421 5823
rect 473 5771 475 5823
rect 419 5699 475 5771
rect 419 5647 421 5699
rect 473 5647 475 5699
rect 419 5411 475 5647
rect 419 5359 421 5411
rect 473 5359 475 5411
rect 419 5287 475 5359
rect 419 5235 421 5287
rect 473 5235 475 5287
rect 419 5163 475 5235
rect 419 5111 421 5163
rect 473 5111 475 5163
rect 419 4875 475 5111
rect 419 4823 421 4875
rect 473 4823 475 4875
rect 419 4751 475 4823
rect 419 4699 421 4751
rect 473 4699 475 4751
rect 419 4627 475 4699
rect 419 4575 421 4627
rect 473 4575 475 4627
rect 419 4339 475 4575
rect 419 4287 421 4339
rect 473 4287 475 4339
rect 419 4215 475 4287
rect 419 4163 421 4215
rect 473 4163 475 4215
rect 419 4091 475 4163
rect 419 4039 421 4091
rect 473 4039 475 4091
rect 419 3803 475 4039
rect 419 3751 421 3803
rect 473 3751 475 3803
rect 419 3679 475 3751
rect 419 3627 421 3679
rect 473 3627 475 3679
rect 419 3555 475 3627
rect 419 3503 421 3555
rect 473 3503 475 3555
rect 419 3267 475 3503
rect 419 3215 421 3267
rect 473 3215 475 3267
rect 419 3143 475 3215
rect 419 3091 421 3143
rect 473 3091 475 3143
rect 419 3019 475 3091
rect 419 2967 421 3019
rect 473 2967 475 3019
rect 419 2731 475 2967
rect 419 2679 421 2731
rect 473 2679 475 2731
rect 419 2607 475 2679
rect 419 2555 421 2607
rect 473 2555 475 2607
rect 419 2483 475 2555
rect 419 2431 421 2483
rect 473 2431 475 2483
rect 419 2195 475 2431
rect 419 2143 421 2195
rect 473 2143 475 2195
rect 419 2071 475 2143
rect 419 2019 421 2071
rect 473 2019 475 2071
rect 419 1947 475 2019
rect 419 1895 421 1947
rect 473 1895 475 1947
rect 419 1659 475 1895
rect 419 1607 421 1659
rect 473 1607 475 1659
rect 419 1535 475 1607
rect 419 1483 421 1535
rect 473 1483 475 1535
rect 419 1411 475 1483
rect 419 1359 421 1411
rect 473 1359 475 1411
rect 419 1123 475 1359
rect 419 1071 421 1123
rect 473 1071 475 1123
rect 419 999 475 1071
rect 419 947 421 999
rect 473 947 475 999
rect 419 875 475 947
rect 419 823 421 875
rect 473 823 475 875
rect 419 587 475 823
rect 419 535 421 587
rect 473 535 475 587
rect 419 463 475 535
rect 419 411 421 463
rect 473 411 475 463
rect 419 339 475 411
rect 419 287 421 339
rect 473 287 475 339
rect 419 51 475 287
rect 419 -1 421 51
rect 473 -1 475 51
rect 419 -73 475 -1
rect 419 -125 421 -73
rect 473 -125 475 -73
rect 419 -197 475 -125
rect 419 -249 421 -197
rect 473 -249 475 -197
rect 419 -485 475 -249
rect 419 -537 421 -485
rect 473 -537 475 -485
rect 419 -609 475 -537
rect 419 -661 421 -609
rect 473 -661 475 -609
rect 419 -733 475 -661
rect 419 -785 421 -733
rect 473 -785 475 -733
rect 419 -1021 475 -785
rect 419 -1073 421 -1021
rect 473 -1073 475 -1021
rect 419 -1145 475 -1073
rect 419 -1197 421 -1145
rect 473 -1197 475 -1145
rect 419 -1269 475 -1197
rect 419 -1321 421 -1269
rect 473 -1321 475 -1269
rect 419 -1557 475 -1321
rect 419 -1609 421 -1557
rect 473 -1609 475 -1557
rect 419 -1681 475 -1609
rect 419 -1733 421 -1681
rect 473 -1733 475 -1681
rect 419 -1805 475 -1733
rect 419 -1857 421 -1805
rect 473 -1857 475 -1805
rect 419 -1981 475 -1857
rect 503 6145 559 6521
rect 503 6093 505 6145
rect 557 6093 559 6145
rect 503 6037 559 6093
rect 503 5985 505 6037
rect 557 5985 559 6037
rect 503 5609 559 5985
rect 503 5557 505 5609
rect 557 5557 559 5609
rect 503 5501 559 5557
rect 503 5449 505 5501
rect 557 5449 559 5501
rect 503 5073 559 5449
rect 503 5021 505 5073
rect 557 5021 559 5073
rect 503 4965 559 5021
rect 503 4913 505 4965
rect 557 4913 559 4965
rect 503 4537 559 4913
rect 503 4485 505 4537
rect 557 4485 559 4537
rect 503 4429 559 4485
rect 503 4377 505 4429
rect 557 4377 559 4429
rect 503 4001 559 4377
rect 503 3949 505 4001
rect 557 3949 559 4001
rect 503 3893 559 3949
rect 503 3841 505 3893
rect 557 3841 559 3893
rect 503 3465 559 3841
rect 503 3413 505 3465
rect 557 3413 559 3465
rect 503 3357 559 3413
rect 503 3305 505 3357
rect 557 3305 559 3357
rect 503 2929 559 3305
rect 503 2877 505 2929
rect 557 2877 559 2929
rect 503 2821 559 2877
rect 503 2769 505 2821
rect 557 2769 559 2821
rect 503 2393 559 2769
rect 503 2341 505 2393
rect 557 2341 559 2393
rect 503 2285 559 2341
rect 503 2233 505 2285
rect 557 2233 559 2285
rect 503 1857 559 2233
rect 503 1805 505 1857
rect 557 1805 559 1857
rect 503 1749 559 1805
rect 503 1697 505 1749
rect 557 1697 559 1749
rect 503 1321 559 1697
rect 503 1269 505 1321
rect 557 1269 559 1321
rect 503 1213 559 1269
rect 503 1161 505 1213
rect 557 1161 559 1213
rect 503 785 559 1161
rect 503 733 505 785
rect 557 733 559 785
rect 503 677 559 733
rect 503 625 505 677
rect 557 625 559 677
rect 503 249 559 625
rect 503 197 505 249
rect 557 197 559 249
rect 503 141 559 197
rect 503 89 505 141
rect 557 89 559 141
rect 503 -287 559 89
rect 503 -339 505 -287
rect 557 -339 559 -287
rect 503 -395 559 -339
rect 503 -447 505 -395
rect 557 -447 559 -395
rect 503 -823 559 -447
rect 503 -875 505 -823
rect 557 -875 559 -823
rect 503 -931 559 -875
rect 503 -983 505 -931
rect 557 -983 559 -931
rect 503 -1359 559 -983
rect 503 -1411 505 -1359
rect 557 -1411 559 -1359
rect 503 -1467 559 -1411
rect 503 -1519 505 -1467
rect 557 -1519 559 -1467
rect 503 -1895 559 -1519
rect 587 6483 643 6489
rect 587 6431 589 6483
rect 641 6431 643 6483
rect 587 6359 643 6431
rect 587 6307 589 6359
rect 641 6307 643 6359
rect 587 6235 643 6307
rect 587 6183 589 6235
rect 641 6183 643 6235
rect 587 5947 643 6183
rect 587 5895 589 5947
rect 641 5895 643 5947
rect 587 5823 643 5895
rect 587 5771 589 5823
rect 641 5771 643 5823
rect 587 5699 643 5771
rect 587 5647 589 5699
rect 641 5647 643 5699
rect 587 5411 643 5647
rect 587 5359 589 5411
rect 641 5359 643 5411
rect 587 5287 643 5359
rect 587 5235 589 5287
rect 641 5235 643 5287
rect 587 5163 643 5235
rect 587 5111 589 5163
rect 641 5111 643 5163
rect 587 4875 643 5111
rect 587 4823 589 4875
rect 641 4823 643 4875
rect 587 4751 643 4823
rect 587 4699 589 4751
rect 641 4699 643 4751
rect 587 4627 643 4699
rect 587 4575 589 4627
rect 641 4575 643 4627
rect 587 4339 643 4575
rect 587 4287 589 4339
rect 641 4287 643 4339
rect 587 4215 643 4287
rect 587 4163 589 4215
rect 641 4163 643 4215
rect 587 4091 643 4163
rect 587 4039 589 4091
rect 641 4039 643 4091
rect 587 3803 643 4039
rect 587 3751 589 3803
rect 641 3751 643 3803
rect 587 3679 643 3751
rect 587 3627 589 3679
rect 641 3627 643 3679
rect 587 3555 643 3627
rect 587 3503 589 3555
rect 641 3503 643 3555
rect 587 3267 643 3503
rect 587 3215 589 3267
rect 641 3215 643 3267
rect 587 3143 643 3215
rect 587 3091 589 3143
rect 641 3091 643 3143
rect 587 3019 643 3091
rect 587 2967 589 3019
rect 641 2967 643 3019
rect 995 3085 1051 3091
rect 995 3033 997 3085
rect 1049 3033 1051 3085
rect 587 2731 643 2967
rect 587 2679 589 2731
rect 641 2679 643 2731
rect 587 2607 643 2679
rect 587 2555 589 2607
rect 641 2555 643 2607
rect 587 2483 643 2555
rect 587 2431 589 2483
rect 641 2431 643 2483
rect 587 2195 643 2431
rect 587 2143 589 2195
rect 641 2143 643 2195
rect 587 2071 643 2143
rect 587 2019 589 2071
rect 641 2019 643 2071
rect 587 1947 643 2019
rect 587 1895 589 1947
rect 641 1895 643 1947
rect 587 1659 643 1895
rect 587 1607 589 1659
rect 641 1607 643 1659
rect 587 1535 643 1607
rect 587 1483 589 1535
rect 641 1483 643 1535
rect 587 1411 643 1483
rect 587 1359 589 1411
rect 641 1359 643 1411
rect 587 1123 643 1359
rect 587 1071 589 1123
rect 641 1071 643 1123
rect 587 999 643 1071
rect 587 947 589 999
rect 641 947 643 999
rect 587 875 643 947
rect 587 823 589 875
rect 641 823 643 875
rect 587 587 643 823
rect 587 535 589 587
rect 641 535 643 587
rect 587 463 643 535
rect 587 411 589 463
rect 641 411 643 463
rect 587 339 643 411
rect 587 287 589 339
rect 641 287 643 339
rect 587 51 643 287
rect 587 -1 589 51
rect 641 -1 643 51
rect 587 -73 643 -1
rect 587 -125 589 -73
rect 641 -125 643 -73
rect 587 -197 643 -125
rect 587 -249 589 -197
rect 641 -249 643 -197
rect 587 -485 643 -249
rect 587 -537 589 -485
rect 641 -537 643 -485
rect 587 -609 643 -537
rect 587 -661 589 -609
rect 641 -661 643 -609
rect 587 -733 643 -661
rect 587 -785 589 -733
rect 641 -785 643 -733
rect 587 -1021 643 -785
rect 587 -1073 589 -1021
rect 641 -1073 643 -1021
rect 587 -1145 643 -1073
rect 587 -1197 589 -1145
rect 641 -1197 643 -1145
rect 587 -1269 643 -1197
rect 587 -1321 589 -1269
rect 641 -1321 643 -1269
rect 587 -1557 643 -1321
rect 587 -1609 589 -1557
rect 641 -1609 643 -1557
rect 587 -1681 643 -1609
rect 587 -1733 589 -1681
rect 641 -1733 643 -1681
rect 587 -1805 643 -1733
rect 587 -1857 589 -1805
rect 641 -1857 643 -1805
rect 587 -1863 643 -1857
rect 911 2956 967 3010
rect 911 2904 913 2956
rect 965 2904 967 2956
rect 911 2638 967 2904
rect 911 2586 913 2638
rect 965 2586 967 2638
rect 911 2320 967 2586
rect 911 2268 913 2320
rect 965 2268 967 2320
rect 911 2002 967 2268
rect 911 1950 913 2002
rect 965 1950 967 2002
rect 911 1684 967 1950
rect 911 1632 913 1684
rect 965 1632 967 1684
rect 911 1366 967 1632
rect 911 1314 913 1366
rect 965 1314 967 1366
rect 911 1048 967 1314
rect 911 996 913 1048
rect 965 996 967 1048
rect 911 730 967 996
rect 911 678 913 730
rect 965 678 967 730
rect 911 412 967 678
rect 911 360 913 412
rect 965 360 967 412
rect 911 94 967 360
rect 911 42 913 94
rect 965 42 967 94
rect 911 -224 967 42
rect 911 -276 913 -224
rect 965 -276 967 -224
rect 911 -542 967 -276
rect 911 -594 913 -542
rect 965 -594 967 -542
rect 911 -860 967 -594
rect 911 -912 913 -860
rect 965 -912 967 -860
rect 911 -1178 967 -912
rect 911 -1230 913 -1178
rect 965 -1230 967 -1178
rect 911 -1496 967 -1230
rect 911 -1548 913 -1496
rect 965 -1548 967 -1496
rect 911 -1814 967 -1548
rect 911 -1866 913 -1814
rect 965 -1866 967 -1814
rect 911 -1872 967 -1866
rect 995 2875 1051 3033
rect 995 2823 997 2875
rect 1049 2823 1051 2875
rect 995 2767 1051 2823
rect 995 2715 997 2767
rect 1049 2715 1051 2767
rect 995 2557 1051 2715
rect 995 2505 997 2557
rect 1049 2505 1051 2557
rect 995 2449 1051 2505
rect 995 2397 997 2449
rect 1049 2397 1051 2449
rect 995 2239 1051 2397
rect 995 2187 997 2239
rect 1049 2187 1051 2239
rect 995 2131 1051 2187
rect 995 2079 997 2131
rect 1049 2079 1051 2131
rect 995 1921 1051 2079
rect 995 1869 997 1921
rect 1049 1869 1051 1921
rect 995 1813 1051 1869
rect 995 1761 997 1813
rect 1049 1761 1051 1813
rect 995 1603 1051 1761
rect 995 1551 997 1603
rect 1049 1551 1051 1603
rect 995 1495 1051 1551
rect 995 1443 997 1495
rect 1049 1443 1051 1495
rect 995 1285 1051 1443
rect 995 1233 997 1285
rect 1049 1233 1051 1285
rect 995 1177 1051 1233
rect 995 1125 997 1177
rect 1049 1125 1051 1177
rect 995 967 1051 1125
rect 995 915 997 967
rect 1049 915 1051 967
rect 995 859 1051 915
rect 995 807 997 859
rect 1049 807 1051 859
rect 995 649 1051 807
rect 995 597 997 649
rect 1049 597 1051 649
rect 995 541 1051 597
rect 995 489 997 541
rect 1049 489 1051 541
rect 995 331 1051 489
rect 995 279 997 331
rect 1049 279 1051 331
rect 995 223 1051 279
rect 995 171 997 223
rect 1049 171 1051 223
rect 995 13 1051 171
rect 995 -39 997 13
rect 1049 -39 1051 13
rect 995 -95 1051 -39
rect 995 -147 997 -95
rect 1049 -147 1051 -95
rect 995 -305 1051 -147
rect 995 -357 997 -305
rect 1049 -357 1051 -305
rect 995 -413 1051 -357
rect 995 -465 997 -413
rect 1049 -465 1051 -413
rect 995 -623 1051 -465
rect 995 -675 997 -623
rect 1049 -675 1051 -623
rect 995 -731 1051 -675
rect 995 -783 997 -731
rect 1049 -783 1051 -731
rect 995 -941 1051 -783
rect 995 -993 997 -941
rect 1049 -993 1051 -941
rect 995 -1049 1051 -993
rect 995 -1101 997 -1049
rect 1049 -1101 1051 -1049
rect 995 -1259 1051 -1101
rect 995 -1311 997 -1259
rect 1049 -1311 1051 -1259
rect 995 -1367 1051 -1311
rect 995 -1419 997 -1367
rect 1049 -1419 1051 -1367
rect 995 -1577 1051 -1419
rect 995 -1629 997 -1577
rect 1049 -1629 1051 -1577
rect 995 -1685 1051 -1629
rect 995 -1737 997 -1685
rect 1049 -1737 1051 -1685
rect 503 -1947 505 -1895
rect 557 -1947 559 -1895
rect 503 -1953 559 -1947
rect 995 -1895 1051 -1737
rect 995 -1947 997 -1895
rect 1049 -1947 1051 -1895
rect 995 -1953 1051 -1947
rect 1079 2956 1135 3010
rect 1079 2904 1081 2956
rect 1133 2904 1135 2956
rect 1079 2638 1135 2904
rect 1079 2586 1081 2638
rect 1133 2586 1135 2638
rect 1079 2320 1135 2586
rect 1079 2268 1081 2320
rect 1133 2268 1135 2320
rect 1079 2002 1135 2268
rect 1079 1950 1081 2002
rect 1133 1950 1135 2002
rect 1079 1684 1135 1950
rect 1079 1632 1081 1684
rect 1133 1632 1135 1684
rect 1079 1366 1135 1632
rect 1079 1314 1081 1366
rect 1133 1314 1135 1366
rect 1079 1048 1135 1314
rect 1079 996 1081 1048
rect 1133 996 1135 1048
rect 1079 730 1135 996
rect 1079 678 1081 730
rect 1133 678 1135 730
rect 1079 412 1135 678
rect 1079 360 1081 412
rect 1133 360 1135 412
rect 1079 94 1135 360
rect 1079 42 1081 94
rect 1133 42 1135 94
rect 1079 -224 1135 42
rect 1079 -276 1081 -224
rect 1133 -276 1135 -224
rect 1079 -542 1135 -276
rect 1079 -594 1081 -542
rect 1133 -594 1135 -542
rect 1079 -860 1135 -594
rect 1079 -912 1081 -860
rect 1133 -912 1135 -860
rect 1079 -1178 1135 -912
rect 1079 -1230 1081 -1178
rect 1133 -1230 1135 -1178
rect 1079 -1496 1135 -1230
rect 1079 -1548 1081 -1496
rect 1133 -1548 1135 -1496
rect 1079 -1814 1135 -1548
rect 1079 -1866 1081 -1814
rect 1133 -1866 1135 -1814
rect 419 -2033 421 -1981
rect 473 -2033 475 -1981
rect 419 -2324 475 -2033
rect 1079 -1981 1135 -1866
rect 1079 -2033 1081 -1981
rect 1133 -2033 1135 -1981
rect 1079 -2039 1135 -2033
rect 419 -2376 421 -2324
rect 473 -2376 475 -2324
rect 419 -2382 475 -2376
use sky130_fd_pr__pfet_01v8_GN49S6  XM1
timestamp 1730624594
transform 1 0 531 0 1 2313
box -246 -4389 246 4389
use sky130_fd_pr__nfet_01v8_GPU48F  XM2
timestamp 1730624594
transform 1 0 1023 0 1 569
box -246 -2645 246 2645
<< labels >>
flabel metal1 285 -2172 381 -2076 0 FreeSans 320 0 0 0 vdda
port 1 nsew
flabel metal1 285 -2296 381 -2200 0 FreeSans 320 0 0 0 vssa
port 4 nsew
flabel metal1 285 -2382 343 -2324 0 FreeSans 320 0 0 0 in
port 5 nsew
flabel via1 997 -1947 1049 -1895 0 FreeSans 320 0 0 0 swn
port 3 nsew
flabel via1 505 -1947 557 -1895 0 FreeSans 320 0 0 0 swp
port 2 nsew
flabel via1 589 6431 641 6483 0 FreeSans 320 0 0 0 out
port 6 nsew
<< end >>
