magic
tech sky130A
magscale 1 2
timestamp 1730296483
<< checkpaint >>
rect 2780 -6070 5792 -1530
<< error_s >>
rect 298 -1085 333 -1051
rect 299 -1104 333 -1085
rect 318 -2017 333 -1104
rect 352 -1138 387 -1104
rect 667 -1138 702 -1104
rect 352 -2017 386 -1138
rect 668 -1157 702 -1138
rect 498 -1206 556 -1200
rect 498 -1240 510 -1206
rect 498 -1246 556 -1240
rect 498 -1934 556 -1928
rect 498 -1968 510 -1934
rect 498 -1974 556 -1968
rect 352 -2051 367 -2017
rect 687 -2070 702 -1157
rect 721 -1191 756 -1157
rect 721 -2070 755 -1191
rect 867 -1259 925 -1253
rect 867 -1293 879 -1259
rect 867 -1299 925 -1293
rect 1037 -1592 1071 -1574
rect 1037 -1628 1107 -1592
rect 1054 -1662 1125 -1628
rect 1405 -1662 1440 -1628
rect 867 -1987 925 -1981
rect 867 -2021 879 -1987
rect 867 -2027 925 -2021
rect 721 -2104 736 -2070
rect 1054 -2123 1124 -1662
rect 1406 -1681 1440 -1662
rect 1236 -1730 1294 -1724
rect 1236 -1764 1248 -1730
rect 1236 -1770 1294 -1764
rect 1236 -2040 1294 -2034
rect 1236 -2074 1248 -2040
rect 1236 -2080 1294 -2074
rect 1054 -2159 1107 -2123
rect 1425 -2176 1440 -1681
rect 1459 -1715 1494 -1681
rect 1774 -1715 1809 -1681
rect 1459 -2176 1493 -1715
rect 1775 -1734 1809 -1715
rect 1605 -1783 1663 -1777
rect 1605 -1817 1617 -1783
rect 1605 -1823 1663 -1817
rect 1605 -2093 1663 -2087
rect 1605 -2127 1617 -2093
rect 1605 -2133 1663 -2127
rect 1459 -2210 1474 -2176
rect 1794 -2229 1809 -1734
rect 1828 -1768 1863 -1734
rect 2143 -1768 2178 -1734
rect 1828 -2229 1862 -1768
rect 2144 -1787 2178 -1768
rect 1974 -1836 2032 -1830
rect 1974 -1870 1986 -1836
rect 1974 -1876 2032 -1870
rect 1974 -2146 2032 -2140
rect 1974 -2180 1986 -2146
rect 1974 -2186 2032 -2180
rect 1828 -2263 1843 -2229
rect 2163 -2282 2178 -1787
rect 2197 -1821 2232 -1787
rect 2512 -1821 2547 -1787
rect 2197 -2282 2231 -1821
rect 2513 -1840 2547 -1821
rect 2343 -1889 2401 -1883
rect 2343 -1923 2355 -1889
rect 2343 -1929 2401 -1923
rect 2343 -2199 2401 -2193
rect 2343 -2233 2355 -2199
rect 2343 -2239 2401 -2233
rect 2197 -2316 2212 -2282
rect 2532 -2335 2547 -1840
rect 2566 -1874 2601 -1840
rect 2881 -1874 2916 -1840
rect 2566 -2335 2600 -1874
rect 2882 -1893 2916 -1874
rect 2712 -1942 2770 -1936
rect 2712 -1976 2724 -1942
rect 2712 -1982 2770 -1976
rect 2712 -2252 2770 -2246
rect 2712 -2286 2724 -2252
rect 2712 -2292 2770 -2286
rect 2566 -2369 2581 -2335
rect 2901 -2388 2916 -1893
rect 2935 -1927 2970 -1893
rect 2935 -2388 2969 -1927
rect 3081 -1995 3139 -1989
rect 3081 -2029 3093 -1995
rect 3081 -2035 3139 -2029
rect 3081 -2305 3139 -2299
rect 3081 -2339 3093 -2305
rect 3081 -2345 3139 -2339
rect 2935 -2422 2950 -2388
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__cap_mim_m3_1_V2UT89  XC1
timestamp 0
transform 1 0 3707 0 1 -3317
box -386 -1440 386 1440
use sky130_fd_pr__pfet_01v8_XGSNAL  XM1
timestamp 0
transform 1 0 158 0 1 -1534
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM2
timestamp 0
transform 1 0 527 0 1 -1587
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM3
timestamp 0
transform 1 0 896 0 1 -1640
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 0
transform 1 0 1265 0 1 -1902
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM5
timestamp 0
transform 1 0 1634 0 1 -1955
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM6
timestamp 0
transform 1 0 2003 0 1 -2008
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM7
timestamp 0
transform 1 0 2372 0 1 -2061
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM8
timestamp 0
transform 1 0 2741 0 1 -2114
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM9
timestamp 0
transform 1 0 3110 0 1 -2167
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_RYGWKL  XM10
timestamp 0
transform 1 0 4286 0 1 -3800
box -246 -1010 246 1010
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 clk
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 clkb
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 vi
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vo
port 5 nsew
<< end >>
