magic
tech sky130A
magscale 1 2
timestamp 1730625751
<< metal1 >>
rect 2177 844 2361 850
rect 2177 672 2183 844
rect 2355 672 2361 844
rect 2177 666 2361 672
rect 674 -10318 1617 -10312
rect 674 -10410 680 -10318
rect 772 -10410 1519 -10318
rect 1611 -10410 1617 -10318
rect 674 -10416 1617 -10410
rect 1513 -11038 1961 -11032
rect 1513 -11130 1519 -11038
rect 1611 -11130 1863 -11038
rect 1955 -11130 1961 -11038
rect 1513 -11136 1961 -11130
rect 2697 -12472 2864 -12471
rect 2530 -12478 2968 -12472
rect 2530 -12570 2536 -12478
rect 2628 -12570 2870 -12478
rect 2962 -12570 2968 -12478
rect 2530 -12575 2968 -12570
rect 2530 -12576 2697 -12575
rect 2801 -12576 2968 -12575
rect 2697 -13124 2801 -13020
rect -14221 -21350 17979 -21344
rect -14221 -21442 680 -21350
rect 772 -21442 17979 -21350
rect -14221 -21448 17979 -21442
rect -14221 -21514 17979 -21508
rect -14221 -21606 2703 -21514
rect 2795 -21606 17979 -21514
rect -14221 -21612 17979 -21606
rect -14221 -21678 17979 -21672
rect -14221 -21770 1863 -21678
rect 1955 -21770 17979 -21678
rect -14221 -21776 17979 -21770
rect -14221 -21842 17979 -21836
rect -14221 -21934 1691 -21842
rect 1783 -21934 17979 -21842
rect -14221 -21940 17979 -21934
rect -14221 -22006 17979 -22000
rect -14221 -22098 2870 -22006
rect 2962 -22098 17979 -22006
rect -14221 -22104 17979 -22098
rect -14221 -22170 17979 -22164
rect -14221 -22262 886 -22170
rect 978 -22262 17979 -22170
rect -14221 -22268 17979 -22262
rect -14221 -22334 17979 -22328
rect -14221 -22426 1691 -22334
rect 1783 -22426 2703 -22334
rect 2795 -22426 17979 -22334
rect -14221 -22432 17979 -22426
rect -14221 -22498 17979 -22492
rect -14221 -22590 680 -22498
rect 772 -22590 3713 -22498
rect 3805 -22590 17979 -22498
rect -14221 -22596 17979 -22590
rect -14221 -22662 17979 -22656
rect -14221 -22754 -734 -22662
rect -642 -22754 5231 -22662
rect 5323 -22754 17979 -22662
rect -14221 -22760 17979 -22754
rect -14221 -22826 17979 -22820
rect -14221 -22918 -3874 -22826
rect -3782 -22918 8266 -22826
rect 8358 -22918 17979 -22826
rect -14221 -22924 17979 -22918
rect -14221 -22990 17979 -22984
rect -14221 -23082 -9946 -22990
rect -9854 -23082 14339 -22990
rect 14431 -23082 17979 -22990
rect -14221 -23088 17979 -23082
<< via1 >>
rect 2183 672 2355 844
rect 680 -10410 772 -10318
rect 1519 -10410 1611 -10318
rect 1519 -11130 1611 -11038
rect 1863 -11130 1955 -11038
rect 2536 -12570 2628 -12478
rect 2870 -12570 2962 -12478
rect 680 -21442 772 -21350
rect 2703 -21606 2795 -21514
rect 1863 -21770 1955 -21678
rect 1691 -21934 1783 -21842
rect 2870 -22098 2962 -22006
rect 886 -22262 978 -22170
rect 1691 -22426 1783 -22334
rect 2703 -22426 2795 -22334
rect 680 -22590 772 -22498
rect 3713 -22590 3805 -22498
rect -734 -22754 -642 -22662
rect 5231 -22754 5323 -22662
rect -3874 -22918 -3782 -22826
rect 8266 -22918 8358 -22826
rect -9946 -23082 -9854 -22990
rect 14339 -23082 14431 -22990
<< metal2 >>
rect 1993 844 2545 850
rect 1993 841 2183 844
rect 2355 841 2545 844
rect 1993 755 1998 841
rect 2540 755 2545 841
rect 1993 746 2183 755
rect 2177 672 2183 746
rect 2355 746 2545 755
rect 2355 672 2361 746
rect 2177 666 2361 672
rect 880 -7817 984 -7808
rect 880 -7903 889 -7817
rect 975 -7903 984 -7817
rect 674 -10318 778 -10312
rect 674 -10410 680 -10318
rect 772 -10410 778 -10318
rect 674 -21350 778 -10410
rect 674 -21442 680 -21350
rect 772 -21442 778 -21350
rect 674 -21448 778 -21442
rect 880 -13921 984 -7903
rect 1685 -9977 1789 -9968
rect 1685 -10063 1694 -9977
rect 1780 -10063 1789 -9977
rect 1513 -10318 1617 -10312
rect 1513 -10410 1519 -10318
rect 1611 -10410 1617 -10318
rect 1513 -10416 1617 -10410
rect 1513 -11038 1617 -11032
rect 1513 -11130 1519 -11038
rect 1611 -11130 1617 -11038
rect 1513 -11136 1617 -11130
rect 880 -14007 889 -13921
rect 975 -14007 984 -13921
rect 880 -22170 984 -14007
rect 1685 -11761 1789 -10063
rect 1685 -11847 1694 -11761
rect 1780 -11847 1789 -11761
rect 1685 -21842 1789 -11847
rect 1857 -10697 2801 -10688
rect 1857 -10783 2697 -10697
rect 2796 -10783 2801 -10697
rect 1857 -10792 2801 -10783
rect 1857 -11038 1961 -10792
rect 1857 -11130 1863 -11038
rect 1955 -11130 1961 -11038
rect 1857 -21678 1961 -11130
rect 2697 -11417 2801 -11408
rect 2697 -11503 2706 -11417
rect 2792 -11503 2801 -11417
rect 2530 -12478 2634 -12472
rect 2530 -12570 2536 -12478
rect 2628 -12570 2634 -12478
rect 2530 -12576 2634 -12570
rect 2697 -21514 2801 -11503
rect 2697 -21606 2703 -21514
rect 2795 -21606 2801 -21514
rect 2697 -21612 2801 -21606
rect 2864 -12478 2968 -12472
rect 2864 -12570 2870 -12478
rect 2962 -12570 2968 -12478
rect 1857 -21770 1863 -21678
rect 1955 -21770 1961 -21678
rect 1857 -21776 1961 -21770
rect 1685 -21934 1691 -21842
rect 1783 -21934 1789 -21842
rect 1685 -21940 1789 -21934
rect 2864 -22006 2968 -12570
rect 2864 -22098 2870 -22006
rect 2962 -22098 2968 -22006
rect 2864 -22104 2968 -22098
rect 880 -22262 886 -22170
rect 978 -22262 984 -22170
rect 880 -22268 984 -22262
rect 1685 -22334 1789 -22328
rect 1685 -22426 1691 -22334
rect 1783 -22426 1789 -22334
rect 1685 -22432 1789 -22426
rect 2697 -22334 2801 -22328
rect 2697 -22426 2703 -22334
rect 2795 -22426 2801 -22334
rect 2697 -22432 2801 -22426
rect 674 -22498 778 -22492
rect 674 -22590 680 -22498
rect 772 -22590 778 -22498
rect 674 -22596 778 -22590
rect 3707 -22498 3811 -22492
rect 3707 -22590 3713 -22498
rect 3805 -22590 3811 -22498
rect 3707 -22596 3811 -22590
rect -740 -22662 -636 -22656
rect -740 -22754 -734 -22662
rect -642 -22754 -636 -22662
rect -740 -22760 -636 -22754
rect 5225 -22662 5329 -22656
rect 5225 -22754 5231 -22662
rect 5323 -22754 5329 -22662
rect 5225 -22760 5329 -22754
rect -3880 -22826 -3776 -22820
rect -3880 -22918 -3874 -22826
rect -3782 -22918 -3776 -22826
rect -3880 -22924 -3776 -22918
rect 8260 -22826 8364 -22820
rect 8260 -22918 8266 -22826
rect 8358 -22918 8364 -22826
rect 8260 -22924 8364 -22918
rect -9952 -22990 -9848 -22984
rect -9952 -23082 -9946 -22990
rect -9854 -23082 -9848 -22990
rect -9952 -23088 -9848 -23082
rect 14333 -22990 14437 -22984
rect 14333 -23082 14339 -22990
rect 14431 -23082 14437 -22990
rect 14333 -23088 14437 -23082
<< via2 >>
rect 1998 755 2183 841
rect 2183 755 2355 841
rect 2355 755 2540 841
rect 2186 752 2352 755
rect 889 -7903 975 -7817
rect 1694 -10063 1780 -9977
rect 1522 -10407 1608 -10321
rect 1522 -11127 1608 -11041
rect 889 -14007 975 -13921
rect 1694 -11847 1780 -11761
rect 2697 -10783 2796 -10697
rect 2706 -11503 2792 -11417
rect 2539 -12567 2625 -12481
rect 1694 -22423 1780 -22337
rect 2706 -22423 2792 -22337
rect 683 -22587 769 -22501
rect 3716 -22587 3802 -22501
rect -731 -22751 -645 -22665
rect 5234 -22751 5320 -22665
rect -3871 -22915 -3785 -22829
rect 8269 -22915 8355 -22829
rect -9943 -23079 -9857 -22993
rect 14342 -23079 14428 -22993
<< metal3 >>
rect 1993 841 2545 850
rect 1993 752 2186 755
rect 2352 752 2545 755
rect 1993 746 2545 752
rect 1394 196 2194 300
rect 880 -4929 1071 -4928
rect 875 -5031 881 -4929
rect 983 -5031 1071 -4929
rect 880 -5032 1071 -5031
rect 1685 -5460 1789 -5272
rect 1457 -5564 2257 -5460
rect 880 -7817 1017 -7808
rect 880 -7903 889 -7817
rect 975 -7903 1017 -7817
rect 880 -7912 1017 -7903
rect 1685 -7912 1789 -5564
rect 2697 -7912 2801 -5272
rect 1457 -8444 2257 -8340
rect 1457 -9884 2257 -9780
rect 1685 -9977 1789 -9968
rect 1685 -10063 1694 -9977
rect 1780 -10063 1789 -9977
rect 1685 -10072 1789 -10063
rect 1513 -10321 1617 -10312
rect 1513 -10407 1522 -10321
rect 1608 -10407 1617 -10321
rect 1513 -10416 1617 -10407
rect 1513 -10674 1651 -10478
rect 1513 -11041 1617 -11032
rect 1513 -11127 1522 -11041
rect 1608 -11127 1617 -11041
rect 1513 -11136 1617 -11127
rect 2139 -11324 2257 -11220
rect 2527 -11369 2617 -11232
rect 2697 -11417 2801 -11408
rect 2697 -11503 2706 -11417
rect 2792 -11503 2801 -11417
rect 2697 -11512 2801 -11503
rect 1685 -11761 1789 -11752
rect 1685 -11847 1694 -11761
rect 1780 -11847 1789 -11761
rect 1685 -11856 1789 -11847
rect 1457 -12045 2257 -11941
rect 2530 -12478 2634 -12472
rect 2530 -12570 2536 -12478
rect 2628 -12570 2634 -12478
rect 2530 -12576 2634 -12570
rect 1457 -12764 2257 -12660
rect 2697 -13672 2801 -12472
rect 880 -13921 1017 -13912
rect 880 -14007 889 -13921
rect 975 -14007 1017 -13921
rect 880 -14016 1017 -14007
rect 1457 -14204 2257 -14100
rect 874 -16896 880 -16792
rect 984 -16896 1017 -16792
rect 1457 -17084 2257 -16980
rect 1685 -22337 1789 -22312
rect 1685 -22423 1694 -22337
rect 1780 -22423 1789 -22337
rect 1685 -22432 1789 -22423
rect 2697 -22337 2801 -22312
rect 2697 -22423 2706 -22337
rect 2792 -22423 2801 -22337
rect 2697 -22432 2801 -22423
rect 674 -22498 778 -22492
rect 674 -22590 680 -22498
rect 772 -22590 778 -22498
rect 674 -22596 778 -22590
rect 3707 -22498 3811 -22492
rect 3707 -22590 3713 -22498
rect 3805 -22590 3811 -22498
rect 3707 -22596 3811 -22590
rect -740 -22662 -636 -22656
rect -740 -22754 -734 -22662
rect -642 -22754 -636 -22662
rect -740 -22760 -636 -22754
rect 5225 -22662 5329 -22656
rect 5225 -22754 5231 -22662
rect 5323 -22754 5329 -22662
rect 5225 -22760 5329 -22754
rect -3880 -22826 -3776 -22820
rect -3880 -22918 -3874 -22826
rect -3782 -22918 -3776 -22826
rect -3880 -22924 -3776 -22918
rect 8260 -22826 8364 -22820
rect 8260 -22918 8266 -22826
rect 8358 -22918 8364 -22826
rect 8260 -22924 8364 -22918
rect -9952 -22990 -9848 -22984
rect -9952 -23082 -9946 -22990
rect -9854 -23082 -9848 -22990
rect -9952 -23088 -9848 -23082
rect 14333 -22990 14437 -22984
rect 14333 -23082 14339 -22990
rect 14431 -23082 14437 -22990
rect 14333 -23088 14437 -23082
<< via3 >>
rect 1993 755 1998 841
rect 1998 755 2540 841
rect 2540 755 2545 841
rect 881 -5031 983 -4929
rect 2536 -12481 2628 -12478
rect 2536 -12567 2539 -12481
rect 2539 -12567 2625 -12481
rect 2625 -12567 2628 -12481
rect 2536 -12570 2628 -12567
rect 880 -16896 984 -16792
rect 680 -22501 772 -22498
rect 680 -22587 683 -22501
rect 683 -22587 769 -22501
rect 769 -22587 772 -22501
rect 680 -22590 772 -22587
rect 3713 -22501 3805 -22498
rect 3713 -22587 3716 -22501
rect 3716 -22587 3802 -22501
rect 3802 -22587 3805 -22501
rect 3713 -22590 3805 -22587
rect -734 -22665 -642 -22662
rect -734 -22751 -731 -22665
rect -731 -22751 -645 -22665
rect -645 -22751 -642 -22665
rect -734 -22754 -642 -22751
rect 5231 -22665 5323 -22662
rect 5231 -22751 5234 -22665
rect 5234 -22751 5320 -22665
rect 5320 -22751 5323 -22665
rect 5231 -22754 5323 -22751
rect -3874 -22829 -3782 -22826
rect -3874 -22915 -3871 -22829
rect -3871 -22915 -3785 -22829
rect -3785 -22915 -3782 -22829
rect -3874 -22918 -3782 -22915
rect 8266 -22829 8358 -22826
rect 8266 -22915 8269 -22829
rect 8269 -22915 8355 -22829
rect 8355 -22915 8358 -22829
rect 8266 -22918 8358 -22915
rect -9946 -22993 -9854 -22990
rect -9946 -23079 -9943 -22993
rect -9943 -23079 -9857 -22993
rect -9857 -23079 -9854 -22993
rect -9946 -23082 -9854 -23079
rect 14339 -22993 14431 -22990
rect 14339 -23079 14342 -22993
rect 14342 -23079 14428 -22993
rect 14428 -23079 14431 -22993
rect 14339 -23082 14431 -23079
<< metal4 >>
rect -13974 841 17499 850
rect -13974 755 1993 841
rect 2545 755 17499 841
rect -13974 746 17499 755
rect -13974 500 -13870 746
rect -12962 504 -12858 746
rect -11950 504 -11846 746
rect -10938 504 -10834 746
rect -9926 504 -9822 746
rect -8914 504 -8810 746
rect -7902 504 -7798 746
rect -6890 504 -6786 746
rect -5878 504 -5774 746
rect -4866 500 -4762 746
rect -3854 504 -3750 746
rect -2842 504 -2738 746
rect -1830 504 -1726 746
rect -818 504 -714 746
rect 194 494 298 746
rect 1205 504 1309 746
rect 2217 504 2321 746
rect 3227 504 3331 746
rect 4239 504 4343 746
rect 5251 504 5355 746
rect 6263 504 6367 746
rect 7275 504 7379 746
rect 8287 504 8391 746
rect 9299 504 9403 746
rect 10311 504 10415 746
rect 11323 504 11427 746
rect 12335 504 12439 746
rect 13347 504 13451 746
rect 14359 504 14463 746
rect 15371 504 15475 746
rect 16383 504 16487 746
rect 17395 504 17499 746
rect 880 -4929 984 -4928
rect 880 -5031 881 -4929
rect 983 -5031 984 -4929
rect 880 -16791 984 -5031
rect 1685 -5032 1789 488
rect 2697 -5032 2801 488
rect 1685 -7912 1789 -5272
rect 2697 -7912 2801 -5272
rect 1685 -9352 1789 -8152
rect 2697 -8700 2801 -8152
rect 2697 -8804 2968 -8700
rect 2697 -9352 2801 -8804
rect 2864 -12472 2968 -8804
rect 1685 -13672 1789 -12472
rect 2530 -12478 2968 -12472
rect 2530 -12570 2536 -12478
rect 2628 -12570 2968 -12478
rect 2530 -12576 2968 -12570
rect 2697 -13672 2801 -12576
rect 1685 -16552 1789 -13912
rect 2697 -16552 2801 -13912
rect 879 -16792 985 -16791
rect 879 -16896 880 -16792
rect 984 -16896 985 -16792
rect 879 -16897 985 -16896
rect 1685 -22312 1789 -16792
rect 2697 -22312 2801 -16792
rect -13494 -22492 -13390 -22328
rect -12482 -22492 -12378 -22328
rect -11470 -22492 -11366 -22328
rect -10458 -22492 -10354 -22328
rect -9446 -22492 -9342 -22328
rect -8434 -22492 -8330 -22328
rect -7422 -22492 -7318 -22328
rect -6410 -22492 -6306 -22328
rect -13494 -22596 -6306 -22492
rect -5398 -22492 -5294 -22328
rect -4386 -22492 -4282 -22328
rect -3374 -22492 -3270 -22328
rect -2362 -22492 -2258 -22328
rect -5398 -22596 -2258 -22492
rect -1350 -22492 -1246 -22328
rect -338 -22492 -234 -22328
rect -1350 -22596 -234 -22492
rect 674 -22492 778 -22328
rect 3707 -22492 3811 -22316
rect 674 -22498 3811 -22492
rect 674 -22590 680 -22498
rect 772 -22590 3713 -22498
rect 3805 -22590 3811 -22498
rect 674 -22596 3811 -22590
rect 4719 -22492 4823 -22328
rect 5731 -22492 5835 -22328
rect 4719 -22596 5835 -22492
rect 6743 -22492 6847 -22328
rect 7755 -22492 7859 -22328
rect 8767 -22492 8871 -22318
rect 9779 -22492 9883 -22328
rect 6743 -22596 9883 -22492
rect 10791 -22492 10895 -22328
rect 11803 -22492 11907 -22328
rect 12815 -22492 12919 -22328
rect 13827 -22492 13931 -22328
rect 14839 -22492 14943 -22328
rect 15851 -22492 15955 -22328
rect 16863 -22492 16967 -22328
rect 17875 -22492 17979 -22310
rect 10791 -22596 17979 -22492
rect -9952 -22984 -9848 -22596
rect -3880 -22820 -3776 -22596
rect -844 -22656 -740 -22596
rect 5225 -22656 5329 -22596
rect -844 -22662 5329 -22656
rect -844 -22754 -734 -22662
rect -642 -22754 5231 -22662
rect 5323 -22754 5329 -22662
rect -844 -22760 5329 -22754
rect 8261 -22820 8365 -22596
rect -3880 -22826 8365 -22820
rect -3880 -22918 -3874 -22826
rect -3782 -22918 8266 -22826
rect 8358 -22918 8365 -22826
rect -3880 -22924 8365 -22918
rect 14333 -22984 14437 -22596
rect -9952 -22990 14437 -22984
rect -9952 -23082 -9946 -22990
rect -9854 -23082 14339 -22990
rect 14431 -23082 14437 -22990
rect -9952 -23088 14437 -23082
use sky130_fd_pr__cap_mim_m3_1_DURRY3  sky130_fd_pr__cap_mim_m3_1_DURRY3_0
timestamp 1730624594
transform 1 0 1909 0 1 -10912
box -892 -11520 892 11520
use sky130_fd_pr__cap_mim_m3_1_RV4AQU  sky130_fd_pr__cap_mim_m3_1_RV4AQU_1
timestamp 1730624594
transform 1 0 -6692 0 1 -10912
box -7470 -11520 7470 11520
use sky130_fd_pr__cap_mim_m3_1_RV4AQU  sky130_fd_pr__cap_mim_m3_1_RV4AQU_2
timestamp 1730624594
transform 1 0 10509 0 1 -10912
box -7470 -11520 7470 11520
<< labels >>
flabel metal4 2267 646 2267 648 0 FreeSans 1600 0 0 0 VC
port 0 nsew
flabel metal3 2566 -11300 2566 -11300 0 FreeSans 1600 0 0 0 SW[0]
port 2 nsew
flabel metal4 904 -6972 904 -6972 0 FreeSans 1600 0 0 0 SW[5]
port 7 nsew
flabel metal4 818 -22570 818 -22570 0 FreeSans 1600 0 0 0 SW[6]
port 8 nsew
flabel metal4 1558 -22728 1558 -22728 0 FreeSans 1600 0 0 0 SW[7]
port 9 nsew
flabel metal4 2694 -22882 2694 -22882 0 FreeSans 1600 0 0 0 SW[8]
port 10 nsew
flabel metal4 4062 -23044 4062 -23044 0 FreeSans 1600 0 0 0 SW[9]
port 11 nsew
flabel metal3 1586 -10576 1586 -10576 0 FreeSans 1600 0 0 0 VCM
port 1 nsew
flabel metal2 1898 -10944 1898 -10944 0 FreeSans 1600 0 0 0 SW[1]
port 3 nsew
flabel metal3 1905 -9830 1905 -9830 0 FreeSans 1600 0 0 0 SW[2]
port 4 nsew
flabel metal2 885 -13038 885 -13038 0 FreeSans 1600 0 0 0 SW[4]
port 6 nsew
flabel metal4 2922 -12200 2922 -12200 0 FreeSans 1600 0 0 0 SW[3]
port 5 nsew
<< end >>
