magic
tech sky130A
magscale 1 2
timestamp 1731494802
<< metal2 >>
rect 436952 695977 439452 695982
rect 436948 695960 439456 695977
rect 436948 693504 436959 695960
rect 437495 693504 439456 695960
rect 436948 693487 439456 693504
rect 436952 641422 439452 693487
rect 441476 641430 444961 641442
rect 436952 641400 441050 641422
rect 436956 641022 441050 641400
rect 436956 640634 439452 641022
rect 440650 639028 441050 641022
rect 441476 641054 444564 641430
rect 444940 641054 444961 641430
rect 441476 641042 444961 641054
rect 441476 641036 443784 641042
rect 441476 639060 441876 641036
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 436959 693504 437495 695960
rect 444564 641054 444940 641430
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 414690 688724 417190 702300
rect 466498 695982 468998 702300
rect 435002 695960 468998 695982
rect 435002 693504 436959 695960
rect 437495 693504 468998 695960
rect 435002 693482 468998 693504
rect 510594 702268 515394 704800
rect 520594 702268 525394 704800
rect 414690 686224 445982 688724
rect -800 680242 1700 685242
rect -800 643842 1660 648642
rect 443482 641430 445982 686224
rect 456473 683230 470876 683236
rect 510594 683230 525394 702268
rect 456473 683220 525394 683230
rect 456473 668836 456482 683220
rect 470866 669002 525394 683220
rect 566594 683202 571594 704800
rect 566594 681494 571590 683202
rect 533622 679494 571614 681494
rect 576886 681290 584800 682984
rect 470866 668836 524997 669002
rect 456473 668827 524997 668836
rect 456473 668821 470876 668827
rect 475053 663900 477051 663905
rect 533636 663900 535636 679494
rect 576886 679306 578102 681290
rect 580086 679306 584800 681290
rect 576886 677984 584800 679306
rect 475052 663892 535636 663900
rect 475052 661908 475060 663892
rect 477044 661908 535636 663892
rect 475052 661900 535636 661908
rect 475053 661895 477051 661900
rect 443482 641054 444564 641430
rect 444940 641054 445982 641430
rect 443482 640550 445982 641054
rect 530342 639784 584800 644584
rect 530342 639780 582350 639784
rect -800 633842 1660 638642
rect 530342 634584 582320 639780
rect 530342 629784 584800 634584
rect 530342 629230 545142 629784
rect 493910 629084 545142 629230
rect 493900 629069 545142 629084
rect 456472 625572 470778 625588
rect 456472 623668 456513 625572
rect 470737 623668 470778 625572
rect 456472 623652 470778 623668
rect 412884 619175 415366 619180
rect 412884 619165 412933 619175
rect 412700 618565 412933 619165
rect 412884 618551 412933 618565
rect 415317 618551 415366 619175
rect 412884 618546 415366 618551
rect 450516 617774 452516 617782
rect 450516 615790 450524 617774
rect 452508 615790 452516 617774
rect 450516 615782 452516 615790
rect 493900 614445 493930 629069
rect 495754 614445 545142 629069
rect 493900 614430 545142 614445
rect 583520 589472 584800 589584
rect 512412 588402 583520 588550
rect 512412 588290 584800 588402
rect 512412 588154 583520 588290
rect -800 559442 1660 564242
rect 486008 555294 487844 555322
rect -800 549442 1660 554242
rect 486008 540590 486054 555294
rect 487798 540590 487844 555294
rect 486008 540562 487844 540590
rect 489940 520210 491874 520234
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 489940 505506 489955 520210
rect 491859 505506 491874 520210
rect 489940 505482 491874 505506
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 471554 450324 471948 450329
rect 512412 450324 512808 588154
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 534510 555354 584800 555362
rect 534510 540570 534524 555354
rect 549308 550562 584800 555354
rect 549308 545366 582348 550562
rect 549308 545362 583270 545366
rect 549308 540570 584800 545362
rect 534510 540562 584800 540570
rect 583520 500050 584800 500162
rect 515414 499132 583534 499134
rect 471553 450318 512808 450324
rect 471553 449934 471559 450318
rect 471943 449934 512808 450318
rect 471553 449928 512808 449934
rect 515408 498980 583534 499132
rect 515408 498868 584800 498980
rect 515408 498734 583534 498868
rect 471554 449923 471948 449928
rect 467022 448376 467450 448386
rect 515408 448376 515808 498734
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 583520 455628 584800 455740
rect 467022 448368 515808 448376
rect 467022 447984 467046 448368
rect 467430 447984 515808 448368
rect 467022 447976 515808 447984
rect 518376 454558 583528 454698
rect 518376 454446 584800 454558
rect 518376 454298 583528 454446
rect 467022 447966 467450 447976
rect 462579 445142 462977 445147
rect 518376 445142 518776 454298
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 462578 445134 518776 445142
rect 462578 444750 462586 445134
rect 462970 444750 518776 445134
rect 462578 444742 518776 444750
rect 462579 444737 462977 444742
rect 458254 434996 458654 435010
rect 441574 434927 441975 434928
rect 441569 434919 441980 434927
rect 437667 434875 438068 434876
rect 437662 434867 438073 434875
rect 417206 434826 417605 434848
rect 417205 434817 417606 434826
rect 412630 434796 413031 434797
rect 412625 434788 413036 434796
rect 412625 434404 412638 434788
rect 413022 434404 413036 434788
rect 412625 434397 413036 434404
rect 417205 434433 417213 434817
rect 417597 434433 417606 434817
rect 433586 434796 433987 434797
rect 433581 434788 433992 434796
rect 429600 434740 430001 434741
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect -800 16910 480 17022
rect -800 15728 480 15840
rect -800 14546 480 14658
rect -800 13364 480 13476
rect 412630 12436 413031 434397
rect 417205 18350 417606 434433
rect 429595 434732 430006 434740
rect 429595 434348 429608 434732
rect 429992 434348 430006 434732
rect 433581 434404 433594 434788
rect 433978 434404 433992 434788
rect 437662 434483 437675 434867
rect 438059 434483 438073 434867
rect 441569 434535 441582 434919
rect 441966 434535 441980 434919
rect 441569 434528 441980 434535
rect 445496 434912 445906 434926
rect 445496 434528 445509 434912
rect 445893 434528 445906 434912
rect 437662 434476 438073 434483
rect 433581 434397 433992 434404
rect 429595 434341 430006 434348
rect 417205 17966 417213 18350
rect 417597 17966 417606 18350
rect 417205 17952 417606 17966
rect 429600 19264 430001 434341
rect 433586 228104 433987 434397
rect 433586 227286 433988 228104
rect 433588 23090 433988 227286
rect 437667 49554 438068 434476
rect 441574 94212 441975 434528
rect 445496 434514 445906 434528
rect 450016 434820 450432 434836
rect 445501 282190 445901 434514
rect 450016 434436 450033 434820
rect 450417 434436 450432 434820
rect 450016 434422 450432 434436
rect 453984 434754 454384 434768
rect 450025 318648 450425 434422
rect 453984 434370 453992 434754
rect 454376 434370 454384 434754
rect 453984 432758 454384 434370
rect 458254 434612 458262 434996
rect 458646 434612 458654 434996
rect 453978 363868 454378 432758
rect 458254 410274 458654 434612
rect 583520 411206 584800 411318
rect 458254 410136 583526 410274
rect 458254 410024 584800 410136
rect 458254 409874 583526 410024
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 453978 363714 583524 363868
rect 453978 363602 584800 363714
rect 453978 363468 583524 363602
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 583520 319562 584800 319674
rect 450020 318492 583524 318648
rect 450020 318380 584800 318492
rect 450020 318248 583524 318380
rect 450030 318246 450425 318248
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 445500 282006 445901 282190
rect 445500 274212 445900 282006
rect 583520 275140 584800 275252
rect 445500 274070 583526 274212
rect 445500 273958 584800 274070
rect 445500 273812 583526 273958
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 545546 196230 560302 196236
rect 545546 196204 584800 196230
rect 545546 181500 545572 196204
rect 560276 191430 584800 196204
rect 560276 186230 581188 191430
rect 560276 181500 584800 186230
rect 545546 181474 584800 181500
rect 545546 181468 560302 181474
rect 582340 181430 584800 181474
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect 583520 95118 584800 95230
rect 441574 94048 583524 94212
rect 441574 93936 584800 94048
rect 441574 93812 583524 93936
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 437667 49390 583530 49554
rect 437667 49278 584800 49390
rect 437667 49154 583530 49278
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 583520 24002 584800 24114
rect 433588 22932 583526 23090
rect 433588 22820 584800 22932
rect 433588 22690 583526 22820
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 429600 18348 430000 19264
rect 429600 18204 583522 18348
rect 429600 18092 584800 18204
rect 429600 17948 583522 18092
rect 583520 16910 584800 17022
rect 583520 15728 584800 15840
rect 583520 14546 584800 14658
rect 583520 13364 584800 13476
rect 412630 12294 583538 12436
rect -800 12182 480 12294
rect 412630 12182 584800 12294
rect 412630 12036 583538 12182
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect 417200 7722 417611 7730
rect 417200 7720 417213 7722
rect -800 7454 480 7566
rect 417164 7338 417213 7720
rect 417597 7720 417611 7722
rect 417597 7566 583544 7720
rect 417597 7454 584800 7566
rect 417597 7338 583544 7454
rect 417164 7320 583544 7338
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 456482 668836 470866 683220
rect 578102 679306 580086 681290
rect 475060 661908 477044 663892
rect 456513 623668 470737 625572
rect 412933 618551 415317 619175
rect 450524 615790 452508 617774
rect 493930 614445 495754 629069
rect 486054 540590 487798 555294
rect 489955 505506 491859 520210
rect 534524 540570 549308 555354
rect 471559 449934 471943 450318
rect 467046 447984 467430 448368
rect 462586 444750 462970 445134
rect 412638 434404 413022 434788
rect 417213 434433 417597 434817
rect 429608 434348 429992 434732
rect 433594 434404 433978 434788
rect 437675 434483 438059 434867
rect 441582 434535 441966 434919
rect 445509 434528 445893 434912
rect 417213 17966 417597 18350
rect 450033 434436 450417 434820
rect 453992 434370 454376 434754
rect 458262 434612 458646 434996
rect 545572 181500 560276 196204
rect 417213 7338 417597 7722
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 330544 673274 333044 702300
rect 450516 688276 580094 688358
rect 450516 686440 450598 688276
rect 452434 686440 580094 688276
rect 450516 686358 580094 686440
rect 456472 683220 470877 683231
rect 330544 673262 415394 673274
rect 330544 670786 412906 673262
rect 415382 670786 415394 673262
rect 330544 670774 415394 670786
rect 456472 668836 456482 683220
rect 470866 668836 470877 683220
rect 578094 681290 580094 686358
rect 578094 679306 578102 681290
rect 580086 679306 580094 681290
rect 578094 679298 580094 679306
rect 456472 668826 470877 668836
rect 475052 663892 477052 663900
rect 475052 661908 475060 663892
rect 477044 661908 477052 663892
rect 475052 661900 477052 661908
rect 493909 629069 495775 629085
rect 456481 625572 470769 625589
rect 456481 623668 456513 625572
rect 470737 623668 470769 625572
rect 456481 623651 470769 623668
rect 475052 621713 477052 621795
rect 475052 619877 475134 621713
rect 476970 619877 477052 621713
rect 475052 619795 477052 619877
rect 412893 619175 415357 619181
rect 412893 618551 412933 619175
rect 415317 618551 415357 619175
rect 412893 618545 415357 618551
rect 450515 617774 452517 617783
rect 450515 615790 450524 617774
rect 452508 615790 452517 617774
rect 450515 615781 452517 615790
rect 493909 614445 493930 629069
rect 495754 614445 495775 629069
rect 493909 614429 495775 614445
rect 534515 555354 549317 555363
rect 486017 555294 487835 555323
rect 486017 540590 486054 555294
rect 487798 540590 487835 555294
rect 486017 540561 487835 540590
rect 534515 540570 534524 555354
rect 549308 540570 549317 555354
rect 534515 540561 549317 540570
rect 489949 520210 491865 520235
rect 489949 505506 489955 520210
rect 491859 505506 491865 520210
rect 489949 505481 491865 505506
rect 545546 520178 560302 520238
rect 545546 505542 545606 520178
rect 560242 505542 560302 520178
rect 471553 450318 471949 450324
rect 471553 449934 471559 450318
rect 471943 449934 471949 450318
rect 471553 449928 471949 449934
rect 467038 448368 467438 448376
rect 467038 447984 467046 448368
rect 467430 447984 467438 448368
rect 467038 447976 467438 447984
rect 462578 445134 462978 445142
rect 462578 444750 462586 445134
rect 462970 444750 462978 445134
rect 462578 444742 462978 444750
rect 458253 434996 458655 435005
rect 441574 434919 441975 434928
rect 437667 434867 438068 434876
rect 417205 434817 417606 434843
rect 412630 434788 413031 434797
rect 412630 434404 412638 434788
rect 413022 434404 413031 434788
rect 417205 434433 417213 434817
rect 417597 434433 417606 434817
rect 433586 434788 433987 434797
rect 417205 434408 417606 434433
rect 429600 434732 430001 434741
rect 412630 434396 413031 434404
rect 429600 434348 429608 434732
rect 429992 434348 430001 434732
rect 433586 434404 433594 434788
rect 433978 434404 433987 434788
rect 437667 434483 437675 434867
rect 438059 434483 438068 434867
rect 441574 434535 441582 434919
rect 441966 434535 441975 434919
rect 441574 434527 441975 434535
rect 445501 434912 445901 434920
rect 445501 434528 445509 434912
rect 445893 434528 445901 434912
rect 445501 434520 445901 434528
rect 450025 434820 450425 434828
rect 437667 434475 438068 434483
rect 450025 434436 450033 434820
rect 450417 434436 450425 434820
rect 450025 434428 450425 434436
rect 453983 434754 454385 434763
rect 433586 434396 433987 434404
rect 453983 434370 453992 434754
rect 454376 434370 454385 434754
rect 458253 434612 458262 434996
rect 458646 434612 458655 434996
rect 458253 434603 458655 434612
rect 453983 434361 454385 434370
rect 429600 434340 430001 434348
rect 545546 196231 560302 505542
rect 545545 196204 560303 196231
rect 545545 181500 545572 196204
rect 560276 181500 560303 196204
rect 545545 181473 560303 181500
rect 417204 18350 417607 18360
rect 417204 17966 417213 18350
rect 417597 17966 417607 18350
rect 417204 17957 417607 17966
rect 417205 7722 417606 17957
rect 417205 7338 417213 7722
rect 417597 7338 417606 7722
rect 417205 7330 417606 7338
<< via4 >>
rect 450598 686440 452434 688276
rect 412906 670786 415382 673262
rect 456516 668869 470832 683185
rect 475134 661982 476970 663818
rect 456627 623702 470623 625538
rect 475134 619877 476970 621713
rect 413047 618585 415203 619141
rect 450598 615865 452434 617701
rect 486168 540624 487684 555260
rect 534597 540644 549233 555280
rect 489989 505540 491825 520176
rect 545606 505542 560242 520178
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 450516 688276 452516 688358
rect 450516 686440 450598 688276
rect 452434 686440 452516 688276
rect 412870 673262 415418 673298
rect 412870 670786 412906 673262
rect 415382 670786 415418 673262
rect 412870 670750 415418 670786
rect 412894 619204 415394 670750
rect 412870 619141 415394 619204
rect 412870 618585 413047 619141
rect 415203 618585 415394 619141
rect 412870 618546 415394 618585
rect 412870 618522 415380 618546
rect 450516 617807 452516 686440
rect 456448 683185 470901 683253
rect 456448 668869 456516 683185
rect 470832 668869 470901 683185
rect 456448 668802 470901 668869
rect 456473 625612 470876 668802
rect 456458 625538 470876 625612
rect 456458 623702 456627 625538
rect 470623 623702 470876 625538
rect 456458 623628 470876 623702
rect 456473 623609 470876 623628
rect 475052 663818 477052 663900
rect 475052 661982 475134 663818
rect 476970 661982 477052 663818
rect 475052 621819 477052 661982
rect 475028 621713 477076 621819
rect 475028 619877 475134 621713
rect 476970 619877 477076 621713
rect 475028 619771 477076 619877
rect 450491 617701 452541 617807
rect 450491 615865 450598 617701
rect 452434 615865 452541 617701
rect 450491 615759 452541 615865
rect 534491 555362 549339 555387
rect 486018 555346 549339 555362
rect 485994 555280 549339 555346
rect 485994 555260 534597 555280
rect 485994 540624 486168 555260
rect 487684 540644 534597 555260
rect 549233 540644 549339 555280
rect 487684 540624 549339 540644
rect 485994 540562 549339 540624
rect 485994 540538 487858 540562
rect 534491 540537 549339 540562
rect 489926 520238 491888 520258
rect 545522 520238 560326 520262
rect 489926 520178 560326 520238
rect 489926 520176 545606 520178
rect 489926 505540 489989 520176
rect 491825 505542 545606 520176
rect 560242 505542 560326 520178
rect 491825 505540 560326 505542
rect 489926 505482 560326 505540
rect 489926 505458 491888 505482
rect 545522 505458 560326 505482
use tsar_adc  tsar_adc_0
timestamp 1731494658
transform -1 0 -3592898 0 1 2576019
box -4088868 -2142525 -3979350 -1936460
<< labels >>
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 2188 0 0 0 gpio_analog[2]
port 1 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 2188 0 0 0 gpio_analog[3]
port 2 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 2188 0 0 0 gpio_analog[4]
port 3 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 2188 0 0 0 gpio_analog[5]
port 4 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 2188 0 0 0 gpio_analog[6]
port 5 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 2188 0 0 0 gpio_noesd[2]
port 6 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 2188 0 0 0 gpio_noesd[3]
port 7 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 2188 0 0 0 gpio_noesd[4]
port 8 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 2188 0 0 0 gpio_noesd[5]
port 9 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 2188 0 0 0 gpio_noesd[6]
port 10 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 2188 0 0 0 io_analog[0]
port 11 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 3750 180 0 0 io_analog[1]
port 12 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 3750 180 0 0 io_analog[2]
port 13 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 3750 180 0 0 io_analog[3]
port 14 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 3750 180 0 0 io_analog[4]
port 15 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 3750 180 0 0 io_analog[4]
port 15 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 3750 180 0 0 io_analog[4]
port 15 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 3750 180 0 0 io_analog[4]
port 15 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 3750 180 0 0 io_analog[4]
port 15 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 3750 180 0 0 io_analog[4]
port 15 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 3750 180 0 0 io_clamp_high[0]
port 16 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 3750 180 0 0 io_clamp_low[0]
port 17 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 2188 0 0 0 io_in[10]
port 18 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 2188 0 0 0 io_in[11]
port 19 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 2188 0 0 0 io_in[12]
port 20 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 2188 0 0 0 io_in[13]
port 21 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 2188 0 0 0 io_in[9]
port 22 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 2188 0 0 0 io_in_3v3[10]
port 23 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 2188 0 0 0 io_in_3v3[11]
port 24 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 2188 0 0 0 io_in_3v3[12]
port 25 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 2188 0 0 0 io_in_3v3[13]
port 26 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 2188 0 0 0 io_in_3v3[9]
port 27 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 2188 0 0 0 io_oeb[10]
port 28 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 2188 0 0 0 io_oeb[11]
port 29 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 2188 0 0 0 io_oeb[12]
port 30 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 2188 0 0 0 io_oeb[13]
port 31 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 2188 0 0 0 io_oeb[9]
port 32 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 2188 0 0 0 io_out[10]
port 33 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 2188 0 0 0 io_out[11]
port 34 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 2188 0 0 0 io_out[12]
port 35 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 2188 0 0 0 io_out[13]
port 36 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 2188 0 0 0 io_out[9]
port 37 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 2188 0 0 0 vccd1
port 38 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 2188 0 0 0 vccd1
port 38 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 2188 0 0 0 vdda1
port 39 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 2188 0 0 0 vdda1
port 39 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 2188 0 0 0 vdda1
port 39 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 2188 0 0 0 vdda1
port 39 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 3750 180 0 0 vssa1
port 40 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 3750 180 0 0 vssa1
port 40 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 2188 0 0 0 vssa1
port 40 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 2188 0 0 0 vssa1
port 40 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 2188 0 0 0 io_in[16]
port 41 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 2188 0 0 0 io_in[17]
port 42 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 2188 0 0 0 gpio_analog[9]
port 43 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 2188 0 0 0 gpio_noesd[10]
port 44 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 3750 180 0 0 io_analog[5]
port 45 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 3750 180 0 0 io_analog[5]
port 45 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 3750 180 0 0 io_analog[5]
port 45 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 3750 180 0 0 io_analog[5]
port 45 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 3750 180 0 0 io_analog[5]
port 45 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 3750 180 0 0 io_analog[5]
port 45 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 3750 180 0 0 io_analog[6]
port 46 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 3750 180 0 0 io_analog[6]
port 46 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 3750 180 0 0 io_analog[6]
port 46 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 3750 180 0 0 io_analog[6]
port 46 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 3750 180 0 0 io_analog[6]
port 46 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 3750 180 0 0 io_analog[6]
port 46 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 3750 180 0 0 io_analog[7]
port 47 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 2188 0 0 0 io_in_3v3[14]
port 48 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 2188 0 0 0 io_in_3v3[15]
port 49 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 2188 0 0 0 io_in_3v3[16]
port 50 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 2188 0 0 0 io_in_3v3[17]
port 51 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 3750 180 0 0 io_analog[8]
port 52 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 3750 180 0 0 io_analog[9]
port 53 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 2188 0 0 0 gpio_noesd[7]
port 54 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 2188 0 0 0 io_oeb[14]
port 55 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 2188 0 0 0 io_oeb[15]
port 56 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 2188 0 0 0 io_oeb[16]
port 57 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 2188 0 0 0 io_oeb[17]
port 58 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 2188 0 0 0 gpio_noesd[8]
port 59 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 3750 180 0 0 io_clamp_high[1]
port 60 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 3750 180 0 0 io_clamp_high[2]
port 61 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 2188 0 0 0 gpio_noesd[9]
port 62 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 3750 180 0 0 io_clamp_low[1]
port 63 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 2188 0 0 0 io_out[14]
port 64 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 2188 0 0 0 io_out[15]
port 65 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 2188 0 0 0 io_out[16]
port 66 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 2188 0 0 0 io_out[17]
port 67 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 3750 180 0 0 io_clamp_low[2]
port 68 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 2188 0 0 0 gpio_analog[10]
port 69 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 2188 0 0 0 io_analog[10]
port 70 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 2188 0 0 0 vccd2
port 71 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 2188 0 0 0 vccd2
port 71 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 2188 0 0 0 gpio_analog[7]
port 72 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 2188 0 0 0 gpio_analog[8]
port 73 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 2188 0 0 0 io_in[14]
port 74 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 2188 0 0 0 io_in[15]
port 75 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 2188 0 0 0 vssa2
port 76 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 2188 0 0 0 vssa2
port 76 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 2188 0 0 0 io_in_3v3[24]
port 77 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 2188 0 0 0 io_in_3v3[25]
port 78 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 2188 0 0 0 io_in_3v3[26]
port 79 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 2188 0 0 0 gpio_analog[16]
port 80 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 2188 0 0 0 gpio_analog[17]
port 81 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 2188 0 0 0 gpio_analog[11]
port 82 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 2188 0 0 0 gpio_analog[12]
port 83 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 2188 0 0 0 gpio_noesd[11]
port 84 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 2188 0 0 0 io_in[18]
port 85 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 2188 0 0 0 io_in[19]
port 86 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 2188 0 0 0 io_in[20]
port 87 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 2188 0 0 0 io_in[21]
port 88 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 2188 0 0 0 io_oeb[18]
port 89 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 2188 0 0 0 io_oeb[19]
port 90 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 2188 0 0 0 io_oeb[20]
port 91 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 2188 0 0 0 io_oeb[21]
port 92 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 2188 0 0 0 io_oeb[22]
port 93 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 2188 0 0 0 io_oeb[23]
port 94 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 2188 0 0 0 io_oeb[24]
port 95 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 2188 0 0 0 io_oeb[25]
port 96 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 2188 0 0 0 io_oeb[26]
port 97 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 2188 0 0 0 io_in[22]
port 98 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 2188 0 0 0 io_in[23]
port 99 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 2188 0 0 0 io_in[24]
port 100 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 2188 0 0 0 io_in[25]
port 101 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 2188 0 0 0 io_in[26]
port 102 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 2188 0 0 0 gpio_noesd[12]
port 103 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 2188 0 0 0 gpio_noesd[13]
port 104 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 2188 0 0 0 gpio_noesd[14]
port 105 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 2188 0 0 0 gpio_noesd[15]
port 106 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 2188 0 0 0 io_out[18]
port 107 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 2188 0 0 0 io_out[19]
port 108 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 2188 0 0 0 io_out[20]
port 109 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 2188 0 0 0 io_out[21]
port 110 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 2188 0 0 0 io_out[22]
port 111 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 2188 0 0 0 io_out[23]
port 112 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 2188 0 0 0 io_out[24]
port 113 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 2188 0 0 0 io_out[25]
port 114 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 2188 0 0 0 io_out[26]
port 115 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 2188 0 0 0 gpio_noesd[16]
port 116 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 2188 0 0 0 gpio_noesd[17]
port 117 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 2188 0 0 0 gpio_analog[13]
port 118 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 2188 0 0 0 gpio_analog[14]
port 119 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 2188 0 0 0 gpio_analog[15]
port 120 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 2188 0 0 0 io_in_3v3[18]
port 121 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 2188 0 0 0 io_in_3v3[19]
port 122 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 2188 0 0 0 vdda2
port 123 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 2188 0 0 0 vdda2
port 123 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 2188 0 0 0 io_in_3v3[20]
port 124 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 2188 0 0 0 io_in_3v3[21]
port 125 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 2188 0 0 0 io_in_3v3[22]
port 126 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 2188 0 0 0 io_in_3v3[23]
port 127 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 2188 0 0 0 vssd2
port 128 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 2188 0 0 0 vssd2
port 128 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 2188 0 0 0 io_in_3v3[6]
port 129 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 2188 0 0 0 io_in_3v3[7]
port 130 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 2188 0 0 0 io_in_3v3[8]
port 131 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 2188 0 0 0 io_in[1]
port 132 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 2188 0 0 0 io_oeb[0]
port 133 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 2188 0 0 0 gpio_noesd[0]
port 134 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 2188 0 0 0 io_in[2]
port 135 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 2188 0 0 0 io_in[3]
port 136 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 2188 0 0 0 io_in[4]
port 137 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 2188 0 0 0 io_in[5]
port 138 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 2188 0 0 0 io_out[1]
port 139 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 2188 0 0 0 io_in[6]
port 140 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 2188 0 0 0 io_in_3v3[1]
port 141 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 2188 0 0 0 io_in[7]
port 142 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 2188 0 0 0 io_in[8]
port 143 nsew
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 2188 0 0 0 gpio_analog[0]
port 144 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 2188 0 0 0 io_oeb[1]
port 145 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 2188 0 0 0 io_in_3v3[0]
port 146 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 2188 0 0 0 io_out[2]
port 147 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 2188 0 0 0 io_out[3]
port 148 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 2188 0 0 0 io_out[4]
port 149 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 2188 0 0 0 io_out[5]
port 150 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 2188 0 0 0 io_out[6]
port 151 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 2188 0 0 0 io_out[7]
port 152 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 2188 0 0 0 io_out[8]
port 153 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 2188 0 0 0 gpio_analog[1]
port 154 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 2188 0 0 0 gpio_noesd[1]
port 155 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 2188 0 0 0 io_in[0]
port 156 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 2188 0 0 0 io_in_3v3[2]
port 157 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 2188 0 0 0 io_in_3v3[3]
port 158 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 2188 0 0 0 io_in_3v3[4]
port 159 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 2188 0 0 0 io_oeb[2]
port 160 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 2188 0 0 0 io_oeb[3]
port 161 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 2188 0 0 0 io_oeb[4]
port 162 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 2188 0 0 0 io_oeb[5]
port 163 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 2188 0 0 0 io_oeb[6]
port 164 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 2188 0 0 0 io_oeb[7]
port 165 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 2188 0 0 0 io_oeb[8]
port 166 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 2188 0 0 0 vssd1
port 167 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 2188 0 0 0 vssd1
port 167 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 2188 0 0 0 io_in_3v3[5]
port 168 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 2188 0 0 0 io_out[0]
port 169 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 2188 90 0 0 wb_clk_i
port 170 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 2188 90 0 0 wb_rst_i
port 171 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 2188 90 0 0 wbs_ack_o
port 172 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 2188 90 0 0 wbs_adr_i[0]
port 173 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 2188 90 0 0 wbs_adr_i[10]
port 174 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 2188 90 0 0 wbs_adr_i[11]
port 175 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 2188 90 0 0 wbs_adr_i[12]
port 176 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 2188 90 0 0 wbs_adr_i[13]
port 177 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 2188 90 0 0 wbs_adr_i[14]
port 178 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 2188 90 0 0 wbs_adr_i[15]
port 179 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 2188 90 0 0 wbs_adr_i[16]
port 180 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 2188 90 0 0 wbs_adr_i[17]
port 181 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 2188 90 0 0 wbs_adr_i[1]
port 182 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 2188 90 0 0 wbs_adr_i[2]
port 183 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 2188 90 0 0 wbs_adr_i[3]
port 184 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 2188 90 0 0 wbs_adr_i[4]
port 185 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 2188 90 0 0 wbs_adr_i[5]
port 186 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 2188 90 0 0 wbs_adr_i[6]
port 187 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 2188 90 0 0 wbs_adr_i[7]
port 188 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 2188 90 0 0 wbs_adr_i[8]
port 189 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 2188 90 0 0 wbs_adr_i[9]
port 190 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 2188 90 0 0 wbs_cyc_i
port 191 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 2188 90 0 0 wbs_dat_i[0]
port 192 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 2188 90 0 0 wbs_dat_i[10]
port 193 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 2188 90 0 0 wbs_dat_i[11]
port 194 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 2188 90 0 0 wbs_dat_i[12]
port 195 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 2188 90 0 0 wbs_dat_i[13]
port 196 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 2188 90 0 0 wbs_dat_i[14]
port 197 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 2188 90 0 0 wbs_dat_i[15]
port 198 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 2188 90 0 0 wbs_dat_i[16]
port 199 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 2188 90 0 0 wbs_dat_i[1]
port 200 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 2188 90 0 0 wbs_dat_i[2]
port 201 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 2188 90 0 0 wbs_dat_i[3]
port 202 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 2188 90 0 0 wbs_dat_i[4]
port 203 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 2188 90 0 0 wbs_dat_i[5]
port 204 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 2188 90 0 0 wbs_dat_i[6]
port 205 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 2188 90 0 0 wbs_dat_i[7]
port 206 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 2188 90 0 0 wbs_dat_i[8]
port 207 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 2188 90 0 0 wbs_dat_i[9]
port 208 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 2188 90 0 0 wbs_dat_o[0]
port 209 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 2188 90 0 0 wbs_dat_o[10]
port 210 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 2188 90 0 0 wbs_dat_o[11]
port 211 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 2188 90 0 0 wbs_dat_o[12]
port 212 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 2188 90 0 0 wbs_dat_o[13]
port 213 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 2188 90 0 0 wbs_dat_o[14]
port 214 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 2188 90 0 0 wbs_dat_o[15]
port 215 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 2188 90 0 0 wbs_dat_o[16]
port 216 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 2188 90 0 0 wbs_dat_o[1]
port 217 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 2188 90 0 0 wbs_dat_o[2]
port 218 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 2188 90 0 0 wbs_dat_o[3]
port 219 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 2188 90 0 0 wbs_dat_o[4]
port 220 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 2188 90 0 0 wbs_dat_o[5]
port 221 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 2188 90 0 0 wbs_dat_o[6]
port 222 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 2188 90 0 0 wbs_dat_o[7]
port 223 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 2188 90 0 0 wbs_dat_o[8]
port 224 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 2188 90 0 0 wbs_dat_o[9]
port 225 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 2188 90 0 0 wbs_sel_i[0]
port 226 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 2188 90 0 0 wbs_sel_i[1]
port 227 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 2188 90 0 0 wbs_sel_i[2]
port 228 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 2188 90 0 0 wbs_sel_i[3]
port 229 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 2188 90 0 0 wbs_stb_i
port 230 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 2188 90 0 0 wbs_we_i
port 231 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 2188 90 0 0 wbs_dat_i[17]
port 232 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 2188 90 0 0 wbs_dat_i[18]
port 233 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 2188 90 0 0 wbs_dat_i[19]
port 234 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 2188 90 0 0 wbs_adr_i[18]
port 235 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 2188 90 0 0 wbs_dat_i[20]
port 236 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 2188 90 0 0 wbs_dat_i[21]
port 237 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 2188 90 0 0 wbs_dat_i[22]
port 238 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 2188 90 0 0 wbs_dat_i[23]
port 239 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 2188 90 0 0 wbs_dat_i[24]
port 240 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 2188 90 0 0 wbs_dat_i[25]
port 241 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 2188 90 0 0 wbs_dat_i[26]
port 242 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 2188 90 0 0 wbs_dat_i[27]
port 243 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 2188 90 0 0 wbs_dat_i[28]
port 244 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 2188 90 0 0 wbs_dat_i[29]
port 245 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 2188 90 0 0 wbs_adr_i[19]
port 246 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 2188 90 0 0 wbs_dat_i[30]
port 247 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 2188 90 0 0 wbs_dat_i[31]
port 248 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 2188 90 0 0 la_oenb[0]
port 249 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 2188 90 0 0 wbs_adr_i[20]
port 250 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 2188 90 0 0 wbs_adr_i[21]
port 251 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 2188 90 0 0 wbs_adr_i[22]
port 252 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 2188 90 0 0 wbs_adr_i[23]
port 253 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 2188 90 0 0 wbs_adr_i[24]
port 254 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 2188 90 0 0 wbs_adr_i[25]
port 255 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 2188 90 0 0 wbs_adr_i[26]
port 256 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 2188 90 0 0 wbs_adr_i[27]
port 257 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 2188 90 0 0 wbs_adr_i[28]
port 258 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 2188 90 0 0 wbs_adr_i[29]
port 259 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 2188 90 0 0 la_oenb[1]
port 260 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 2188 90 0 0 wbs_adr_i[30]
port 261 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 2188 90 0 0 wbs_adr_i[31]
port 262 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 2188 90 0 0 la_oenb[2]
port 263 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 2188 90 0 0 wbs_dat_o[17]
port 264 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 2188 90 0 0 wbs_dat_o[18]
port 265 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 2188 90 0 0 wbs_dat_o[19]
port 266 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 2188 90 0 0 la_oenb[3]
port 267 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 2188 90 0 0 wbs_dat_o[20]
port 268 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 2188 90 0 0 wbs_dat_o[21]
port 269 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 2188 90 0 0 wbs_dat_o[22]
port 270 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 2188 90 0 0 wbs_dat_o[23]
port 271 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 2188 90 0 0 wbs_dat_o[24]
port 272 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 2188 90 0 0 wbs_dat_o[25]
port 273 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 2188 90 0 0 wbs_dat_o[26]
port 274 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 2188 90 0 0 wbs_dat_o[27]
port 275 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 2188 90 0 0 wbs_dat_o[28]
port 276 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 2188 90 0 0 wbs_dat_o[29]
port 277 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 2188 90 0 0 la_oenb[4]
port 278 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 2188 90 0 0 wbs_dat_o[30]
port 279 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 2188 90 0 0 wbs_dat_o[31]
port 280 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 2188 90 0 0 la_oenb[5]
port 281 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 2188 90 0 0 la_data_in[0]
port 282 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 2188 90 0 0 la_data_in[1]
port 283 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 2188 90 0 0 la_data_in[2]
port 284 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 2188 90 0 0 la_data_in[3]
port 285 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 2188 90 0 0 la_data_in[4]
port 286 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 2188 90 0 0 la_data_in[5]
port 287 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 2188 90 0 0 la_data_out[0]
port 288 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 2188 90 0 0 la_data_out[1]
port 289 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 2188 90 0 0 la_data_out[2]
port 290 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 2188 90 0 0 la_data_out[3]
port 291 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 2188 90 0 0 la_data_out[4]
port 292 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 2188 90 0 0 la_data_out[5]
port 293 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 2188 90 0 0 la_data_in[23]
port 294 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 2188 90 0 0 la_data_in[24]
port 295 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 2188 90 0 0 la_data_in[25]
port 296 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 2188 90 0 0 la_oenb[6]
port 297 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 2188 90 0 0 la_oenb[7]
port 298 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 2188 90 0 0 la_oenb[8]
port 299 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 2188 90 0 0 la_oenb[9]
port 300 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 2188 90 0 0 la_data_in[26]
port 301 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 2188 90 0 0 la_data_in[11]
port 302 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 2188 90 0 0 la_data_in[12]
port 303 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 2188 90 0 0 la_data_in[13]
port 304 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 2188 90 0 0 la_data_in[14]
port 305 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 2188 90 0 0 la_data_in[6]
port 306 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 2188 90 0 0 la_data_in[7]
port 307 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 2188 90 0 0 la_data_in[8]
port 308 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 2188 90 0 0 la_data_in[9]
port 309 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 2188 90 0 0 la_data_in[15]
port 310 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 2188 90 0 0 la_data_out[10]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 2188 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 2188 90 0 0 la_data_out[12]
port 313 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 2188 90 0 0 la_data_out[13]
port 314 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 2188 90 0 0 la_data_out[14]
port 315 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 2188 90 0 0 la_data_out[15]
port 316 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 2188 90 0 0 la_data_out[16]
port 317 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 2188 90 0 0 la_data_out[17]
port 318 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 2188 90 0 0 la_data_out[18]
port 319 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 2188 90 0 0 la_data_out[19]
port 320 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 2188 90 0 0 la_data_in[16]
port 321 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 2188 90 0 0 la_data_out[20]
port 322 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 2188 90 0 0 la_data_out[21]
port 323 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 2188 90 0 0 la_data_out[22]
port 324 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 2188 90 0 0 la_data_out[23]
port 325 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 2188 90 0 0 la_data_out[24]
port 326 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 2188 90 0 0 la_data_out[25]
port 327 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 2188 90 0 0 la_data_in[17]
port 328 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 2188 90 0 0 la_data_in[18]
port 329 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 2188 90 0 0 la_data_in[19]
port 330 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 2188 90 0 0 la_data_in[10]
port 331 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 2188 90 0 0 la_data_out[6]
port 332 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 2188 90 0 0 la_data_out[7]
port 333 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 2188 90 0 0 la_data_out[8]
port 334 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 2188 90 0 0 la_data_out[9]
port 335 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 2188 90 0 0 la_data_in[20]
port 336 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 2188 90 0 0 la_oenb[10]
port 337 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 2188 90 0 0 la_oenb[11]
port 338 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 2188 90 0 0 la_oenb[12]
port 339 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 2188 90 0 0 la_oenb[13]
port 340 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 2188 90 0 0 la_oenb[14]
port 341 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 2188 90 0 0 la_oenb[15]
port 342 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 2188 90 0 0 la_oenb[16]
port 343 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 2188 90 0 0 la_oenb[17]
port 344 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 2188 90 0 0 la_oenb[18]
port 345 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 2188 90 0 0 la_oenb[19]
port 346 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 2188 90 0 0 la_data_in[21]
port 347 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 2188 90 0 0 la_oenb[20]
port 348 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 2188 90 0 0 la_oenb[21]
port 349 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 2188 90 0 0 la_oenb[22]
port 350 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 2188 90 0 0 la_oenb[23]
port 351 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 2188 90 0 0 la_oenb[24]
port 352 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 2188 90 0 0 la_oenb[25]
port 353 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 2188 90 0 0 la_data_in[22]
port 354 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 2188 90 0 0 la_data_in[39]
port 355 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 2188 90 0 0 la_oenb[45]
port 356 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 2188 90 0 0 la_data_in[40]
port 357 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 2188 90 0 0 la_data_out[26]
port 358 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 2188 90 0 0 la_data_out[27]
port 359 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 2188 90 0 0 la_data_out[28]
port 360 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 2188 90 0 0 la_data_out[29]
port 361 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 2188 90 0 0 la_data_in[41]
port 362 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 2188 90 0 0 la_data_out[30]
port 363 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 2188 90 0 0 la_data_out[31]
port 364 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 2188 90 0 0 la_data_out[32]
port 365 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 2188 90 0 0 la_data_out[33]
port 366 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 2188 90 0 0 la_data_out[34]
port 367 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 2188 90 0 0 la_data_out[35]
port 368 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 2188 90 0 0 la_data_out[36]
port 369 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 2188 90 0 0 la_data_out[37]
port 370 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 2188 90 0 0 la_data_out[38]
port 371 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 2188 90 0 0 la_data_out[39]
port 372 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 2188 90 0 0 la_data_in[42]
port 373 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 2188 90 0 0 la_data_out[40]
port 374 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 2188 90 0 0 la_data_out[41]
port 375 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 2188 90 0 0 la_data_out[42]
port 376 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 2188 90 0 0 la_data_out[43]
port 377 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 2188 90 0 0 la_data_out[44]
port 378 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 2188 90 0 0 la_data_out[45]
port 379 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 2188 90 0 0 la_data_out[46]
port 380 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 2188 90 0 0 la_data_in[43]
port 381 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 2188 90 0 0 la_data_in[44]
port 382 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 2188 90 0 0 la_data_in[45]
port 383 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 2188 90 0 0 la_data_in[46]
port 384 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 2188 90 0 0 la_oenb[46]
port 385 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 2188 90 0 0 la_oenb[38]
port 386 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 2188 90 0 0 la_oenb[39]
port 387 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 2188 90 0 0 la_oenb[37]
port 388 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 2188 90 0 0 la_oenb[40]
port 389 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 2188 90 0 0 la_oenb[41]
port 390 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 2188 90 0 0 la_oenb[42]
port 391 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 2188 90 0 0 la_oenb[43]
port 392 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 2188 90 0 0 la_data_in[27]
port 393 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 2188 90 0 0 la_data_in[28]
port 394 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 2188 90 0 0 la_data_in[29]
port 395 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 2188 90 0 0 la_oenb[44]
port 396 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 2188 90 0 0 la_data_in[30]
port 397 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 2188 90 0 0 la_data_in[31]
port 398 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 2188 90 0 0 la_data_in[32]
port 399 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 2188 90 0 0 la_data_in[33]
port 400 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 2188 90 0 0 la_data_in[34]
port 401 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 2188 90 0 0 la_data_in[35]
port 402 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 2188 90 0 0 la_data_in[36]
port 403 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 2188 90 0 0 la_data_in[37]
port 404 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 2188 90 0 0 la_oenb[26]
port 405 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 2188 90 0 0 la_oenb[27]
port 406 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 2188 90 0 0 la_oenb[28]
port 407 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 2188 90 0 0 la_oenb[29]
port 408 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 2188 90 0 0 la_data_in[38]
port 409 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 2188 90 0 0 la_oenb[30]
port 410 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 2188 90 0 0 la_oenb[31]
port 411 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 2188 90 0 0 la_oenb[32]
port 412 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 2188 90 0 0 la_oenb[33]
port 413 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 2188 90 0 0 la_oenb[34]
port 414 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 2188 90 0 0 la_oenb[35]
port 415 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 2188 90 0 0 la_oenb[36]
port 416 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 2188 90 0 0 la_oenb[47]
port 417 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 2188 90 0 0 la_oenb[48]
port 418 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 2188 90 0 0 la_oenb[49]
port 419 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 2188 90 0 0 la_oenb[50]
port 420 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 2188 90 0 0 la_oenb[51]
port 421 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 2188 90 0 0 la_oenb[52]
port 422 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 2188 90 0 0 la_oenb[53]
port 423 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 2188 90 0 0 la_oenb[54]
port 424 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 2188 90 0 0 la_oenb[55]
port 425 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 2188 90 0 0 la_oenb[56]
port 426 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 2188 90 0 0 la_oenb[57]
port 427 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 2188 90 0 0 la_oenb[58]
port 428 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 2188 90 0 0 la_oenb[59]
port 429 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 2188 90 0 0 la_oenb[60]
port 430 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 2188 90 0 0 la_oenb[61]
port 431 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 2188 90 0 0 la_oenb[62]
port 432 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 2188 90 0 0 la_oenb[63]
port 433 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 2188 90 0 0 la_oenb[64]
port 434 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 2188 90 0 0 la_oenb[65]
port 435 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 2188 90 0 0 la_oenb[66]
port 436 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 2188 90 0 0 la_data_in[47]
port 437 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 2188 90 0 0 la_data_in[48]
port 438 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 2188 90 0 0 la_data_in[49]
port 439 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 2188 90 0 0 la_data_in[50]
port 440 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 2188 90 0 0 la_data_in[51]
port 441 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 2188 90 0 0 la_data_in[52]
port 442 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 2188 90 0 0 la_data_in[53]
port 443 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 2188 90 0 0 la_data_in[54]
port 444 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 2188 90 0 0 la_data_in[55]
port 445 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 2188 90 0 0 la_data_in[56]
port 446 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 2188 90 0 0 la_data_in[57]
port 447 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 2188 90 0 0 la_data_in[58]
port 448 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 2188 90 0 0 la_data_in[59]
port 449 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 2188 90 0 0 la_data_in[60]
port 450 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 2188 90 0 0 la_data_in[61]
port 451 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 2188 90 0 0 la_data_in[62]
port 452 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 2188 90 0 0 la_data_in[63]
port 453 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 2188 90 0 0 la_data_out[47]
port 454 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 2188 90 0 0 la_data_out[48]
port 455 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 2188 90 0 0 la_data_out[49]
port 456 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 2188 90 0 0 la_data_in[64]
port 457 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 2188 90 0 0 la_data_out[50]
port 458 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 2188 90 0 0 la_data_out[51]
port 459 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 2188 90 0 0 la_data_out[52]
port 460 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 2188 90 0 0 la_data_out[53]
port 461 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 2188 90 0 0 la_data_out[54]
port 462 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 2188 90 0 0 la_data_out[55]
port 463 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 2188 90 0 0 la_data_out[56]
port 464 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 2188 90 0 0 la_data_out[57]
port 465 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 2188 90 0 0 la_data_out[58]
port 466 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 2188 90 0 0 la_data_out[59]
port 467 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 2188 90 0 0 la_data_in[65]
port 468 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 2188 90 0 0 la_data_out[60]
port 469 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 2188 90 0 0 la_data_out[61]
port 470 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 2188 90 0 0 la_data_out[62]
port 471 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 2188 90 0 0 la_data_out[63]
port 472 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 2188 90 0 0 la_data_out[64]
port 473 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 2188 90 0 0 la_data_out[65]
port 474 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 2188 90 0 0 la_data_out[66]
port 475 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 2188 90 0 0 la_data_out[67]
port 476 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 2188 90 0 0 la_data_in[66]
port 477 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 2188 90 0 0 la_data_in[67]
port 478 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 2188 90 0 0 la_data_in[72]
port 479 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 2188 90 0 0 la_data_in[73]
port 480 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 2188 90 0 0 la_data_in[74]
port 481 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 2188 90 0 0 la_data_in[75]
port 482 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 2188 90 0 0 la_data_in[76]
port 483 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 2188 90 0 0 la_data_in[77]
port 484 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 2188 90 0 0 la_data_in[78]
port 485 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 2188 90 0 0 la_data_in[79]
port 486 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 2188 90 0 0 la_data_in[80]
port 487 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 2188 90 0 0 la_data_in[81]
port 488 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 2188 90 0 0 la_data_in[82]
port 489 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 2188 90 0 0 la_data_in[83]
port 490 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 2188 90 0 0 la_data_in[84]
port 491 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 2188 90 0 0 la_data_in[85]
port 492 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 2188 90 0 0 la_data_in[86]
port 493 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 2188 90 0 0 la_data_in[87]
port 494 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 2188 90 0 0 la_data_in[69]
port 495 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 2188 90 0 0 la_oenb[67]
port 496 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 2188 90 0 0 la_oenb[68]
port 497 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 2188 90 0 0 la_oenb[69]
port 498 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 2188 90 0 0 la_oenb[70]
port 499 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 2188 90 0 0 la_oenb[71]
port 500 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 2188 90 0 0 la_oenb[72]
port 501 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 2188 90 0 0 la_oenb[73]
port 502 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 2188 90 0 0 la_oenb[74]
port 503 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 2188 90 0 0 la_oenb[75]
port 504 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 2188 90 0 0 la_oenb[76]
port 505 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 2188 90 0 0 la_oenb[77]
port 506 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 2188 90 0 0 la_oenb[78]
port 507 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 2188 90 0 0 la_oenb[79]
port 508 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 2188 90 0 0 la_oenb[80]
port 509 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 2188 90 0 0 la_oenb[81]
port 510 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 2188 90 0 0 la_oenb[82]
port 511 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 2188 90 0 0 la_oenb[83]
port 512 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 2188 90 0 0 la_oenb[84]
port 513 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 2188 90 0 0 la_oenb[85]
port 514 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 2188 90 0 0 la_oenb[86]
port 515 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 2188 90 0 0 la_oenb[87]
port 516 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 2188 90 0 0 la_data_out[68]
port 517 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 2188 90 0 0 la_data_out[69]
port 518 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 2188 90 0 0 la_data_in[70]
port 519 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 2188 90 0 0 la_data_out[70]
port 520 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 2188 90 0 0 la_data_out[71]
port 521 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 2188 90 0 0 la_data_out[72]
port 522 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 2188 90 0 0 la_data_out[73]
port 523 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 2188 90 0 0 la_data_out[74]
port 524 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 2188 90 0 0 la_data_out[75]
port 525 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 2188 90 0 0 la_data_out[76]
port 526 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 2188 90 0 0 la_data_out[77]
port 527 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 2188 90 0 0 la_data_out[78]
port 528 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 2188 90 0 0 la_data_out[79]
port 529 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 2188 90 0 0 la_data_in[71]
port 530 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 2188 90 0 0 la_data_out[80]
port 531 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 2188 90 0 0 la_data_out[81]
port 532 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 2188 90 0 0 la_data_out[82]
port 533 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 2188 90 0 0 la_data_out[83]
port 534 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 2188 90 0 0 la_data_out[84]
port 535 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 2188 90 0 0 la_data_out[85]
port 536 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 2188 90 0 0 la_data_out[86]
port 537 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 2188 90 0 0 la_data_out[87]
port 538 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 2188 90 0 0 la_data_in[68]
port 539 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 2188 90 0 0 la_oenb[88]
port 540 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 2188 90 0 0 la_oenb[89]
port 541 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 2188 90 0 0 la_oenb[90]
port 542 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 2188 90 0 0 la_oenb[91]
port 543 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 2188 90 0 0 la_oenb[92]
port 544 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 2188 90 0 0 la_oenb[93]
port 545 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 2188 90 0 0 la_oenb[94]
port 546 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 2188 90 0 0 la_oenb[95]
port 547 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 2188 90 0 0 la_oenb[96]
port 548 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 2188 90 0 0 la_oenb[97]
port 549 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 2188 90 0 0 la_oenb[98]
port 550 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 2188 90 0 0 la_oenb[99]
port 551 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 2188 90 0 0 la_data_in[101]
port 552 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 2188 90 0 0 la_data_in[102]
port 553 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 2188 90 0 0 la_data_in[103]
port 554 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 2188 90 0 0 la_data_in[104]
port 555 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 2188 90 0 0 la_data_in[105]
port 556 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 2188 90 0 0 la_data_in[106]
port 557 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 2188 90 0 0 la_data_in[107]
port 558 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 2188 90 0 0 la_data_in[108]
port 559 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 2188 90 0 0 la_data_in[100]
port 560 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 2188 90 0 0 la_data_in[90]
port 561 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 2188 90 0 0 la_data_in[91]
port 562 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 2188 90 0 0 la_data_in[92]
port 563 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 2188 90 0 0 la_data_in[93]
port 564 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 2188 90 0 0 la_data_in[94]
port 565 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 2188 90 0 0 la_data_in[95]
port 566 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 2188 90 0 0 la_data_in[96]
port 567 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 2188 90 0 0 la_data_in[97]
port 568 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 2188 90 0 0 la_data_in[98]
port 569 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 2188 90 0 0 la_data_in[99]
port 570 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 2188 90 0 0 la_data_out[100]
port 571 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 2188 90 0 0 la_data_out[101]
port 572 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 2188 90 0 0 la_data_out[102]
port 573 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 2188 90 0 0 la_data_out[103]
port 574 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 2188 90 0 0 la_data_out[104]
port 575 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 2188 90 0 0 la_data_out[105]
port 576 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 2188 90 0 0 la_data_out[93]
port 577 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 2188 90 0 0 la_data_out[106]
port 578 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 2188 90 0 0 la_data_out[94]
port 579 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 2188 90 0 0 la_data_out[107]
port 580 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 2188 90 0 0 la_data_out[95]
port 581 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 2188 90 0 0 la_data_out[96]
port 582 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 2188 90 0 0 la_data_out[108]
port 583 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 2188 90 0 0 la_data_out[97]
port 584 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 2188 90 0 0 la_data_out[98]
port 585 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 2188 90 0 0 la_data_out[99]
port 586 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 2188 90 0 0 la_data_out[92]
port 587 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 2188 90 0 0 la_oenb[100]
port 588 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 2188 90 0 0 la_oenb[101]
port 589 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 2188 90 0 0 la_oenb[102]
port 590 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 2188 90 0 0 la_oenb[103]
port 591 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 2188 90 0 0 la_oenb[104]
port 592 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 2188 90 0 0 la_oenb[105]
port 593 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 2188 90 0 0 la_oenb[106]
port 594 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 2188 90 0 0 la_oenb[107]
port 595 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 2188 90 0 0 la_data_in[88]
port 596 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 2188 90 0 0 la_data_in[89]
port 597 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 2188 90 0 0 la_data_out[88]
port 598 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 2188 90 0 0 la_data_out[89]
port 599 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 2188 90 0 0 la_data_out[90]
port 600 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 2188 90 0 0 la_data_out[91]
port 601 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 2188 90 0 0 la_data_in[119]
port 602 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 2188 90 0 0 la_data_out[120]
port 603 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 2188 90 0 0 la_data_out[121]
port 604 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 2188 90 0 0 la_data_out[122]
port 605 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 2188 90 0 0 la_data_in[116]
port 606 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 2188 90 0 0 la_data_in[117]
port 607 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 2188 90 0 0 la_data_out[123]
port 608 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 2188 90 0 0 la_data_in[112]
port 609 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 2188 90 0 0 la_data_out[124]
port 610 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 2188 90 0 0 la_data_out[125]
port 611 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 2188 90 0 0 la_data_out[126]
port 612 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 2188 90 0 0 la_data_out[127]
port 613 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 2188 90 0 0 la_data_in[118]
port 614 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 2188 90 0 0 la_oenb[109]
port 615 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 2188 90 0 0 la_data_in[120]
port 616 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 2188 90 0 0 la_oenb[110]
port 617 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 2188 90 0 0 la_data_in[121]
port 618 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 2188 90 0 0 la_oenb[111]
port 619 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 2188 90 0 0 la_oenb[112]
port 620 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 2188 90 0 0 la_oenb[113]
port 621 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 2188 90 0 0 la_oenb[114]
port 622 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 2188 90 0 0 la_oenb[115]
port 623 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 2188 90 0 0 la_oenb[116]
port 624 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 2188 90 0 0 la_oenb[117]
port 625 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 2188 90 0 0 la_oenb[118]
port 626 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 2188 90 0 0 la_oenb[119]
port 627 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 2188 90 0 0 la_data_in[122]
port 628 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 2188 90 0 0 la_data_in[123]
port 629 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 2188 90 0 0 la_oenb[120]
port 630 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 2188 90 0 0 la_oenb[121]
port 631 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 2188 90 0 0 la_oenb[122]
port 632 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 2188 90 0 0 la_oenb[123]
port 633 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 2188 90 0 0 la_oenb[124]
port 634 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 2188 90 0 0 la_oenb[125]
port 635 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 2188 90 0 0 la_oenb[126]
port 636 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 2188 90 0 0 la_oenb[127]
port 637 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 2188 90 0 0 la_data_in[124]
port 638 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 2188 90 0 0 la_data_in[125]
port 639 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 2188 90 0 0 la_data_in[126]
port 640 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 2188 90 0 0 la_data_in[127]
port 641 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 2188 90 0 0 la_data_out[110]
port 642 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 2188 90 0 0 user_clock2
port 643 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 2188 90 0 0 user_irq[0]
port 644 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 2188 90 0 0 la_data_in[113]
port 645 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 2188 90 0 0 user_irq[1]
port 646 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 2188 90 0 0 la_data_in[114]
port 647 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 2188 90 0 0 user_irq[2]
port 648 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 2188 90 0 0 la_data_out[111]
port 649 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 2188 90 0 0 la_data_out[112]
port 650 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 2188 90 0 0 la_data_out[109]
port 651 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 2188 90 0 0 la_data_in[109]
port 652 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 2188 90 0 0 la_data_out[113]
port 653 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 2188 90 0 0 la_data_in[110]
port 654 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 2188 90 0 0 la_data_out[114]
port 655 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 2188 90 0 0 la_oenb[108]
port 656 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 2188 90 0 0 la_data_out[115]
port 657 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 2188 90 0 0 la_data_out[116]
port 658 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 2188 90 0 0 la_data_in[111]
port 659 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 2188 90 0 0 la_data_out[117]
port 660 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 2188 90 0 0 la_data_in[115]
port 661 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 2188 90 0 0 la_data_out[118]
port 662 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 2188 90 0 0 la_data_out[119]
port 663 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
